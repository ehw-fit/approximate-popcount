// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.09375
// WCE=4.0
// EP=0.726562%
// Printed PDK parameters:
//  Area=28946192.0
//  Delay=54040800.0
//  Power=1322300.0

module popcount18_yobk(input [17:0] input_a, output [4:0] popcount18_yobk_out);
  wire popcount18_yobk_core_020;
  wire popcount18_yobk_core_021;
  wire popcount18_yobk_core_022;
  wire popcount18_yobk_core_023;
  wire popcount18_yobk_core_024_not;
  wire popcount18_yobk_core_026;
  wire popcount18_yobk_core_027;
  wire popcount18_yobk_core_028;
  wire popcount18_yobk_core_030;
  wire popcount18_yobk_core_031;
  wire popcount18_yobk_core_033;
  wire popcount18_yobk_core_035;
  wire popcount18_yobk_core_036;
  wire popcount18_yobk_core_037;
  wire popcount18_yobk_core_038;
  wire popcount18_yobk_core_040;
  wire popcount18_yobk_core_041_not;
  wire popcount18_yobk_core_042;
  wire popcount18_yobk_core_045;
  wire popcount18_yobk_core_048;
  wire popcount18_yobk_core_049;
  wire popcount18_yobk_core_050;
  wire popcount18_yobk_core_051;
  wire popcount18_yobk_core_052;
  wire popcount18_yobk_core_053;
  wire popcount18_yobk_core_054;
  wire popcount18_yobk_core_057;
  wire popcount18_yobk_core_058;
  wire popcount18_yobk_core_061;
  wire popcount18_yobk_core_062;
  wire popcount18_yobk_core_063;
  wire popcount18_yobk_core_064;
  wire popcount18_yobk_core_065;
  wire popcount18_yobk_core_066;
  wire popcount18_yobk_core_067;
  wire popcount18_yobk_core_068;
  wire popcount18_yobk_core_069;
  wire popcount18_yobk_core_070;
  wire popcount18_yobk_core_071_not;
  wire popcount18_yobk_core_073;
  wire popcount18_yobk_core_074;
  wire popcount18_yobk_core_075;
  wire popcount18_yobk_core_076;
  wire popcount18_yobk_core_078;
  wire popcount18_yobk_core_082;
  wire popcount18_yobk_core_083;
  wire popcount18_yobk_core_084;
  wire popcount18_yobk_core_085;
  wire popcount18_yobk_core_086;
  wire popcount18_yobk_core_087;
  wire popcount18_yobk_core_090;
  wire popcount18_yobk_core_091;
  wire popcount18_yobk_core_092;
  wire popcount18_yobk_core_093;
  wire popcount18_yobk_core_094;
  wire popcount18_yobk_core_095;
  wire popcount18_yobk_core_096;
  wire popcount18_yobk_core_097;
  wire popcount18_yobk_core_098;
  wire popcount18_yobk_core_099;
  wire popcount18_yobk_core_100;
  wire popcount18_yobk_core_101;
  wire popcount18_yobk_core_103;
  wire popcount18_yobk_core_106;
  wire popcount18_yobk_core_107;
  wire popcount18_yobk_core_108;
  wire popcount18_yobk_core_111;
  wire popcount18_yobk_core_112;
  wire popcount18_yobk_core_113;
  wire popcount18_yobk_core_114;
  wire popcount18_yobk_core_115;
  wire popcount18_yobk_core_116;
  wire popcount18_yobk_core_117;
  wire popcount18_yobk_core_118;
  wire popcount18_yobk_core_119;
  wire popcount18_yobk_core_120;
  wire popcount18_yobk_core_122;
  wire popcount18_yobk_core_124;

  assign popcount18_yobk_core_020 = ~input_a[4];
  assign popcount18_yobk_core_021 = ~(input_a[1] & input_a[5]);
  assign popcount18_yobk_core_022 = input_a[4] & input_a[16];
  assign popcount18_yobk_core_023 = input_a[7] | input_a[0];
  assign popcount18_yobk_core_024_not = ~input_a[0];
  assign popcount18_yobk_core_026 = input_a[7] | input_a[2];
  assign popcount18_yobk_core_027 = input_a[2] ^ input_a[7];
  assign popcount18_yobk_core_028 = ~popcount18_yobk_core_026;
  assign popcount18_yobk_core_030 = input_a[7] | input_a[2];
  assign popcount18_yobk_core_031 = input_a[16] ^ input_a[10];
  assign popcount18_yobk_core_033 = input_a[11] | input_a[0];
  assign popcount18_yobk_core_035 = input_a[15] | input_a[12];
  assign popcount18_yobk_core_036 = ~input_a[9];
  assign popcount18_yobk_core_037 = input_a[6] | input_a[9];
  assign popcount18_yobk_core_038 = input_a[12] | input_a[16];
  assign popcount18_yobk_core_040 = ~(input_a[2] ^ input_a[2]);
  assign popcount18_yobk_core_041_not = ~input_a[1];
  assign popcount18_yobk_core_042 = ~(input_a[14] | input_a[6]);
  assign popcount18_yobk_core_045 = ~(input_a[14] | input_a[2]);
  assign popcount18_yobk_core_048 = input_a[4] & input_a[1];
  assign popcount18_yobk_core_049 = input_a[17] & input_a[3];
  assign popcount18_yobk_core_050 = popcount18_yobk_core_028 ^ input_a[6];
  assign popcount18_yobk_core_051 = popcount18_yobk_core_028 & input_a[6];
  assign popcount18_yobk_core_052 = popcount18_yobk_core_050 ^ popcount18_yobk_core_049;
  assign popcount18_yobk_core_053 = popcount18_yobk_core_050 & popcount18_yobk_core_049;
  assign popcount18_yobk_core_054 = popcount18_yobk_core_051 | popcount18_yobk_core_053;
  assign popcount18_yobk_core_057 = popcount18_yobk_core_030 ^ popcount18_yobk_core_054;
  assign popcount18_yobk_core_058 = popcount18_yobk_core_030 & popcount18_yobk_core_054;
  assign popcount18_yobk_core_061 = ~(input_a[13] | input_a[8]);
  assign popcount18_yobk_core_062 = input_a[9] ^ input_a[10];
  assign popcount18_yobk_core_063 = input_a[9] & input_a[10];
  assign popcount18_yobk_core_064 = input_a[11] ^ input_a[12];
  assign popcount18_yobk_core_065 = input_a[11] & input_a[12];
  assign popcount18_yobk_core_066 = popcount18_yobk_core_062 ^ popcount18_yobk_core_064;
  assign popcount18_yobk_core_067 = popcount18_yobk_core_062 & popcount18_yobk_core_064;
  assign popcount18_yobk_core_068 = popcount18_yobk_core_063 ^ popcount18_yobk_core_065;
  assign popcount18_yobk_core_069 = popcount18_yobk_core_063 & popcount18_yobk_core_065;
  assign popcount18_yobk_core_070 = popcount18_yobk_core_068 | popcount18_yobk_core_067;
  assign popcount18_yobk_core_071_not = ~input_a[11];
  assign popcount18_yobk_core_073 = input_a[13] ^ input_a[14];
  assign popcount18_yobk_core_074 = input_a[13] & input_a[14];
  assign popcount18_yobk_core_075 = ~(input_a[0] ^ input_a[0]);
  assign popcount18_yobk_core_076 = input_a[0] & input_a[15];
  assign popcount18_yobk_core_078 = ~(input_a[9] ^ input_a[16]);
  assign popcount18_yobk_core_082 = popcount18_yobk_core_073 & input_a[1];
  assign popcount18_yobk_core_083 = popcount18_yobk_core_074 ^ popcount18_yobk_core_076;
  assign popcount18_yobk_core_084 = popcount18_yobk_core_074 & popcount18_yobk_core_076;
  assign popcount18_yobk_core_085 = popcount18_yobk_core_083 ^ popcount18_yobk_core_082;
  assign popcount18_yobk_core_086 = popcount18_yobk_core_083 & popcount18_yobk_core_082;
  assign popcount18_yobk_core_087 = popcount18_yobk_core_084 | popcount18_yobk_core_086;
  assign popcount18_yobk_core_090 = ~(input_a[16] | input_a[1]);
  assign popcount18_yobk_core_091 = popcount18_yobk_core_066 & input_a[8];
  assign popcount18_yobk_core_092 = popcount18_yobk_core_070 ^ popcount18_yobk_core_085;
  assign popcount18_yobk_core_093 = popcount18_yobk_core_070 & popcount18_yobk_core_085;
  assign popcount18_yobk_core_094 = popcount18_yobk_core_092 ^ popcount18_yobk_core_091;
  assign popcount18_yobk_core_095 = popcount18_yobk_core_092 & popcount18_yobk_core_091;
  assign popcount18_yobk_core_096 = popcount18_yobk_core_093 | popcount18_yobk_core_095;
  assign popcount18_yobk_core_097 = popcount18_yobk_core_069 ^ popcount18_yobk_core_087;
  assign popcount18_yobk_core_098 = popcount18_yobk_core_069 & popcount18_yobk_core_087;
  assign popcount18_yobk_core_099 = popcount18_yobk_core_097 ^ popcount18_yobk_core_096;
  assign popcount18_yobk_core_100 = popcount18_yobk_core_097 & popcount18_yobk_core_096;
  assign popcount18_yobk_core_101 = popcount18_yobk_core_098 | popcount18_yobk_core_100;
  assign popcount18_yobk_core_103 = input_a[1] & input_a[16];
  assign popcount18_yobk_core_106 = popcount18_yobk_core_052 ^ popcount18_yobk_core_094;
  assign popcount18_yobk_core_107 = popcount18_yobk_core_052 & popcount18_yobk_core_094;
  assign popcount18_yobk_core_108 = input_a[12] | input_a[0];
  assign popcount18_yobk_core_111 = popcount18_yobk_core_057 ^ popcount18_yobk_core_099;
  assign popcount18_yobk_core_112 = popcount18_yobk_core_057 & popcount18_yobk_core_099;
  assign popcount18_yobk_core_113 = popcount18_yobk_core_111 ^ popcount18_yobk_core_107;
  assign popcount18_yobk_core_114 = popcount18_yobk_core_111 & popcount18_yobk_core_107;
  assign popcount18_yobk_core_115 = popcount18_yobk_core_112 | popcount18_yobk_core_114;
  assign popcount18_yobk_core_116 = popcount18_yobk_core_058 ^ popcount18_yobk_core_101;
  assign popcount18_yobk_core_117 = popcount18_yobk_core_058 & popcount18_yobk_core_101;
  assign popcount18_yobk_core_118 = popcount18_yobk_core_116 | popcount18_yobk_core_115;
  assign popcount18_yobk_core_119 = ~(input_a[16] & input_a[8]);
  assign popcount18_yobk_core_120 = ~input_a[5];
  assign popcount18_yobk_core_122 = input_a[5] ^ input_a[1];
  assign popcount18_yobk_core_124 = ~input_a[7];

  assign popcount18_yobk_out[0] = input_a[5];
  assign popcount18_yobk_out[1] = popcount18_yobk_core_106;
  assign popcount18_yobk_out[2] = popcount18_yobk_core_113;
  assign popcount18_yobk_out[3] = popcount18_yobk_core_118;
  assign popcount18_yobk_out[4] = popcount18_yobk_core_117;
endmodule