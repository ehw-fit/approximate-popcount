// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.18645
// WCE=12.0
// EP=0.859843%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_c58h(input [22:0] input_a, output [4:0] popcount23_c58h_out);
  wire popcount23_c58h_core_025;
  wire popcount23_c58h_core_028;
  wire popcount23_c58h_core_029;
  wire popcount23_c58h_core_031;
  wire popcount23_c58h_core_032;
  wire popcount23_c58h_core_033;
  wire popcount23_c58h_core_038;
  wire popcount23_c58h_core_042;
  wire popcount23_c58h_core_043;
  wire popcount23_c58h_core_044;
  wire popcount23_c58h_core_045;
  wire popcount23_c58h_core_047;
  wire popcount23_c58h_core_048;
  wire popcount23_c58h_core_051;
  wire popcount23_c58h_core_053;
  wire popcount23_c58h_core_054;
  wire popcount23_c58h_core_056_not;
  wire popcount23_c58h_core_058;
  wire popcount23_c58h_core_059;
  wire popcount23_c58h_core_060;
  wire popcount23_c58h_core_061;
  wire popcount23_c58h_core_063;
  wire popcount23_c58h_core_064;
  wire popcount23_c58h_core_065;
  wire popcount23_c58h_core_067;
  wire popcount23_c58h_core_068;
  wire popcount23_c58h_core_069_not;
  wire popcount23_c58h_core_070;
  wire popcount23_c58h_core_071;
  wire popcount23_c58h_core_072;
  wire popcount23_c58h_core_073;
  wire popcount23_c58h_core_074;
  wire popcount23_c58h_core_076;
  wire popcount23_c58h_core_077;
  wire popcount23_c58h_core_078;
  wire popcount23_c58h_core_080;
  wire popcount23_c58h_core_082_not;
  wire popcount23_c58h_core_083;
  wire popcount23_c58h_core_084;
  wire popcount23_c58h_core_087;
  wire popcount23_c58h_core_088;
  wire popcount23_c58h_core_089;
  wire popcount23_c58h_core_090;
  wire popcount23_c58h_core_093;
  wire popcount23_c58h_core_094;
  wire popcount23_c58h_core_098;
  wire popcount23_c58h_core_099;
  wire popcount23_c58h_core_100;
  wire popcount23_c58h_core_102;
  wire popcount23_c58h_core_103;
  wire popcount23_c58h_core_104;
  wire popcount23_c58h_core_105;
  wire popcount23_c58h_core_106;
  wire popcount23_c58h_core_107;
  wire popcount23_c58h_core_108;
  wire popcount23_c58h_core_109;
  wire popcount23_c58h_core_112;
  wire popcount23_c58h_core_114;
  wire popcount23_c58h_core_116;
  wire popcount23_c58h_core_118;
  wire popcount23_c58h_core_119;
  wire popcount23_c58h_core_121;
  wire popcount23_c58h_core_122;
  wire popcount23_c58h_core_124;
  wire popcount23_c58h_core_126;
  wire popcount23_c58h_core_127;
  wire popcount23_c58h_core_128;
  wire popcount23_c58h_core_129;
  wire popcount23_c58h_core_130_not;
  wire popcount23_c58h_core_132;
  wire popcount23_c58h_core_133;
  wire popcount23_c58h_core_138;
  wire popcount23_c58h_core_139;
  wire popcount23_c58h_core_140;
  wire popcount23_c58h_core_141;
  wire popcount23_c58h_core_143;
  wire popcount23_c58h_core_144;
  wire popcount23_c58h_core_145;
  wire popcount23_c58h_core_147;
  wire popcount23_c58h_core_148;
  wire popcount23_c58h_core_149;
  wire popcount23_c58h_core_151_not;
  wire popcount23_c58h_core_152;
  wire popcount23_c58h_core_155;
  wire popcount23_c58h_core_156;
  wire popcount23_c58h_core_157;
  wire popcount23_c58h_core_158;
  wire popcount23_c58h_core_160;
  wire popcount23_c58h_core_161;
  wire popcount23_c58h_core_162;
  wire popcount23_c58h_core_163_not;
  wire popcount23_c58h_core_164;
  wire popcount23_c58h_core_166;

  assign popcount23_c58h_core_025 = input_a[17] & input_a[2];
  assign popcount23_c58h_core_028 = input_a[21] | input_a[14];
  assign popcount23_c58h_core_029 = ~(input_a[4] ^ input_a[18]);
  assign popcount23_c58h_core_031 = input_a[11] | input_a[5];
  assign popcount23_c58h_core_032 = ~(input_a[13] | input_a[1]);
  assign popcount23_c58h_core_033 = ~input_a[10];
  assign popcount23_c58h_core_038 = ~(input_a[6] & input_a[21]);
  assign popcount23_c58h_core_042 = input_a[7] | input_a[1];
  assign popcount23_c58h_core_043 = input_a[5] | input_a[22];
  assign popcount23_c58h_core_044 = ~input_a[11];
  assign popcount23_c58h_core_045 = input_a[18] | input_a[2];
  assign popcount23_c58h_core_047 = ~input_a[18];
  assign popcount23_c58h_core_048 = ~input_a[6];
  assign popcount23_c58h_core_051 = input_a[22] & input_a[14];
  assign popcount23_c58h_core_053 = input_a[4] | input_a[13];
  assign popcount23_c58h_core_054 = ~input_a[22];
  assign popcount23_c58h_core_056_not = ~input_a[19];
  assign popcount23_c58h_core_058 = input_a[5] ^ input_a[3];
  assign popcount23_c58h_core_059 = input_a[6] ^ input_a[7];
  assign popcount23_c58h_core_060 = ~(input_a[6] | input_a[10]);
  assign popcount23_c58h_core_061 = input_a[14] ^ input_a[0];
  assign popcount23_c58h_core_063 = input_a[11] & input_a[11];
  assign popcount23_c58h_core_064 = ~(input_a[21] & input_a[14]);
  assign popcount23_c58h_core_065 = input_a[22] | input_a[20];
  assign popcount23_c58h_core_067 = ~input_a[16];
  assign popcount23_c58h_core_068 = input_a[4] & input_a[1];
  assign popcount23_c58h_core_069_not = ~input_a[12];
  assign popcount23_c58h_core_070 = ~(input_a[4] ^ input_a[2]);
  assign popcount23_c58h_core_071 = ~input_a[0];
  assign popcount23_c58h_core_072 = input_a[11] ^ input_a[7];
  assign popcount23_c58h_core_073 = input_a[2] | input_a[6];
  assign popcount23_c58h_core_074 = ~(input_a[18] & input_a[17]);
  assign popcount23_c58h_core_076 = ~(input_a[7] ^ input_a[14]);
  assign popcount23_c58h_core_077 = ~(input_a[5] ^ input_a[10]);
  assign popcount23_c58h_core_078 = ~(input_a[6] ^ input_a[11]);
  assign popcount23_c58h_core_080 = ~(input_a[1] | input_a[12]);
  assign popcount23_c58h_core_082_not = ~input_a[2];
  assign popcount23_c58h_core_083 = ~(input_a[10] ^ input_a[11]);
  assign popcount23_c58h_core_084 = ~(input_a[19] | input_a[20]);
  assign popcount23_c58h_core_087 = input_a[17] ^ input_a[18];
  assign popcount23_c58h_core_088 = ~(input_a[14] | input_a[7]);
  assign popcount23_c58h_core_089 = ~(input_a[7] ^ input_a[11]);
  assign popcount23_c58h_core_090 = input_a[16] ^ input_a[10];
  assign popcount23_c58h_core_093 = ~(input_a[6] & input_a[12]);
  assign popcount23_c58h_core_094 = input_a[13] ^ input_a[9];
  assign popcount23_c58h_core_098 = ~(input_a[12] | input_a[13]);
  assign popcount23_c58h_core_099 = input_a[14] | input_a[7];
  assign popcount23_c58h_core_100 = ~(input_a[3] & input_a[4]);
  assign popcount23_c58h_core_102 = ~(input_a[9] ^ input_a[3]);
  assign popcount23_c58h_core_103 = ~(input_a[11] ^ input_a[5]);
  assign popcount23_c58h_core_104 = input_a[15] ^ input_a[5];
  assign popcount23_c58h_core_105 = input_a[4] & input_a[10];
  assign popcount23_c58h_core_106 = input_a[1] ^ input_a[4];
  assign popcount23_c58h_core_107 = ~(input_a[0] ^ input_a[17]);
  assign popcount23_c58h_core_108 = ~(input_a[3] ^ input_a[1]);
  assign popcount23_c58h_core_109 = input_a[11] ^ input_a[7];
  assign popcount23_c58h_core_112 = input_a[13] & input_a[16];
  assign popcount23_c58h_core_114 = input_a[14] & input_a[6];
  assign popcount23_c58h_core_116 = ~input_a[19];
  assign popcount23_c58h_core_118 = ~(input_a[8] | input_a[19]);
  assign popcount23_c58h_core_119 = ~(input_a[18] & input_a[3]);
  assign popcount23_c58h_core_121 = ~(input_a[16] | input_a[13]);
  assign popcount23_c58h_core_122 = ~(input_a[11] ^ input_a[11]);
  assign popcount23_c58h_core_124 = ~(input_a[18] ^ input_a[8]);
  assign popcount23_c58h_core_126 = input_a[1] ^ input_a[16];
  assign popcount23_c58h_core_127 = ~(input_a[6] & input_a[18]);
  assign popcount23_c58h_core_128 = input_a[5] ^ input_a[8];
  assign popcount23_c58h_core_129 = ~input_a[1];
  assign popcount23_c58h_core_130_not = ~input_a[20];
  assign popcount23_c58h_core_132 = input_a[22] | input_a[22];
  assign popcount23_c58h_core_133 = ~(input_a[0] | input_a[9]);
  assign popcount23_c58h_core_138 = ~input_a[8];
  assign popcount23_c58h_core_139 = ~(input_a[15] & input_a[14]);
  assign popcount23_c58h_core_140 = input_a[3] & input_a[8];
  assign popcount23_c58h_core_141 = ~(input_a[4] | input_a[3]);
  assign popcount23_c58h_core_143 = ~(input_a[13] ^ input_a[17]);
  assign popcount23_c58h_core_144 = ~(input_a[4] | input_a[6]);
  assign popcount23_c58h_core_145 = input_a[5] & input_a[1];
  assign popcount23_c58h_core_147 = ~(input_a[0] | input_a[11]);
  assign popcount23_c58h_core_148 = input_a[21] & input_a[1];
  assign popcount23_c58h_core_149 = input_a[5] & input_a[21];
  assign popcount23_c58h_core_151_not = ~input_a[0];
  assign popcount23_c58h_core_152 = input_a[15] | input_a[2];
  assign popcount23_c58h_core_155 = ~(input_a[18] & input_a[15]);
  assign popcount23_c58h_core_156 = ~(input_a[3] & input_a[7]);
  assign popcount23_c58h_core_157 = ~(input_a[11] | input_a[12]);
  assign popcount23_c58h_core_158 = input_a[18] ^ input_a[16];
  assign popcount23_c58h_core_160 = ~input_a[10];
  assign popcount23_c58h_core_161 = ~(input_a[1] ^ input_a[13]);
  assign popcount23_c58h_core_162 = ~(input_a[15] | input_a[22]);
  assign popcount23_c58h_core_163_not = ~input_a[11];
  assign popcount23_c58h_core_164 = ~(input_a[18] & input_a[14]);
  assign popcount23_c58h_core_166 = input_a[1] ^ input_a[9];

  assign popcount23_c58h_out[0] = input_a[17];
  assign popcount23_c58h_out[1] = input_a[21];
  assign popcount23_c58h_out[2] = input_a[5];
  assign popcount23_c58h_out[3] = 1'b1;
  assign popcount23_c58h_out[4] = 1'b0;
endmodule