// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5
// WCE=35.0
// EP=0.999994%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_cvsc(input [31:0] input_a, output [5:0] popcount32_cvsc_out);
  wire popcount32_cvsc_core_034;
  wire popcount32_cvsc_core_035;
  wire popcount32_cvsc_core_037;
  wire popcount32_cvsc_core_038_not;
  wire popcount32_cvsc_core_039;
  wire popcount32_cvsc_core_046_not;
  wire popcount32_cvsc_core_048;
  wire popcount32_cvsc_core_049;
  wire popcount32_cvsc_core_052;
  wire popcount32_cvsc_core_053;
  wire popcount32_cvsc_core_056;
  wire popcount32_cvsc_core_057_not;
  wire popcount32_cvsc_core_058;
  wire popcount32_cvsc_core_059;
  wire popcount32_cvsc_core_060;
  wire popcount32_cvsc_core_061;
  wire popcount32_cvsc_core_062;
  wire popcount32_cvsc_core_063;
  wire popcount32_cvsc_core_068;
  wire popcount32_cvsc_core_069;
  wire popcount32_cvsc_core_070;
  wire popcount32_cvsc_core_071;
  wire popcount32_cvsc_core_073;
  wire popcount32_cvsc_core_075;
  wire popcount32_cvsc_core_076;
  wire popcount32_cvsc_core_077;
  wire popcount32_cvsc_core_079;
  wire popcount32_cvsc_core_081;
  wire popcount32_cvsc_core_082;
  wire popcount32_cvsc_core_083;
  wire popcount32_cvsc_core_084;
  wire popcount32_cvsc_core_085;
  wire popcount32_cvsc_core_086;
  wire popcount32_cvsc_core_087;
  wire popcount32_cvsc_core_090;
  wire popcount32_cvsc_core_091;
  wire popcount32_cvsc_core_092;
  wire popcount32_cvsc_core_093;
  wire popcount32_cvsc_core_095;
  wire popcount32_cvsc_core_096;
  wire popcount32_cvsc_core_098;
  wire popcount32_cvsc_core_099_not;
  wire popcount32_cvsc_core_100;
  wire popcount32_cvsc_core_101;
  wire popcount32_cvsc_core_103;
  wire popcount32_cvsc_core_104;
  wire popcount32_cvsc_core_105;
  wire popcount32_cvsc_core_107;
  wire popcount32_cvsc_core_108;
  wire popcount32_cvsc_core_109;
  wire popcount32_cvsc_core_110;
  wire popcount32_cvsc_core_112;
  wire popcount32_cvsc_core_113;
  wire popcount32_cvsc_core_114;
  wire popcount32_cvsc_core_115;
  wire popcount32_cvsc_core_120;
  wire popcount32_cvsc_core_121;
  wire popcount32_cvsc_core_122;
  wire popcount32_cvsc_core_124;
  wire popcount32_cvsc_core_125;
  wire popcount32_cvsc_core_126;
  wire popcount32_cvsc_core_127;
  wire popcount32_cvsc_core_130;
  wire popcount32_cvsc_core_132;
  wire popcount32_cvsc_core_133;
  wire popcount32_cvsc_core_134;
  wire popcount32_cvsc_core_136_not;
  wire popcount32_cvsc_core_138;
  wire popcount32_cvsc_core_139;
  wire popcount32_cvsc_core_141;
  wire popcount32_cvsc_core_142;
  wire popcount32_cvsc_core_144;
  wire popcount32_cvsc_core_145;
  wire popcount32_cvsc_core_147;
  wire popcount32_cvsc_core_148;
  wire popcount32_cvsc_core_151;
  wire popcount32_cvsc_core_152;
  wire popcount32_cvsc_core_155;
  wire popcount32_cvsc_core_156;
  wire popcount32_cvsc_core_159;
  wire popcount32_cvsc_core_166;
  wire popcount32_cvsc_core_167;
  wire popcount32_cvsc_core_168;
  wire popcount32_cvsc_core_169;
  wire popcount32_cvsc_core_171;
  wire popcount32_cvsc_core_172;
  wire popcount32_cvsc_core_173;
  wire popcount32_cvsc_core_174;
  wire popcount32_cvsc_core_175;
  wire popcount32_cvsc_core_179;
  wire popcount32_cvsc_core_180;
  wire popcount32_cvsc_core_181;
  wire popcount32_cvsc_core_182;
  wire popcount32_cvsc_core_183;
  wire popcount32_cvsc_core_186;
  wire popcount32_cvsc_core_187;
  wire popcount32_cvsc_core_188;
  wire popcount32_cvsc_core_192;
  wire popcount32_cvsc_core_193;
  wire popcount32_cvsc_core_197;
  wire popcount32_cvsc_core_199;
  wire popcount32_cvsc_core_200;
  wire popcount32_cvsc_core_202;
  wire popcount32_cvsc_core_203;
  wire popcount32_cvsc_core_204;
  wire popcount32_cvsc_core_205;
  wire popcount32_cvsc_core_206;
  wire popcount32_cvsc_core_207;
  wire popcount32_cvsc_core_208;
  wire popcount32_cvsc_core_209;
  wire popcount32_cvsc_core_210;
  wire popcount32_cvsc_core_211;
  wire popcount32_cvsc_core_212;
  wire popcount32_cvsc_core_213;
  wire popcount32_cvsc_core_214;
  wire popcount32_cvsc_core_215;
  wire popcount32_cvsc_core_216;
  wire popcount32_cvsc_core_217;
  wire popcount32_cvsc_core_218;
  wire popcount32_cvsc_core_220;
  wire popcount32_cvsc_core_222;
  wire popcount32_cvsc_core_223;
  wire popcount32_cvsc_core_224;
  wire popcount32_cvsc_core_225;

  assign popcount32_cvsc_core_034 = ~input_a[31];
  assign popcount32_cvsc_core_035 = input_a[21] & input_a[13];
  assign popcount32_cvsc_core_037 = input_a[21] | input_a[30];
  assign popcount32_cvsc_core_038_not = ~input_a[27];
  assign popcount32_cvsc_core_039 = ~(input_a[9] & input_a[23]);
  assign popcount32_cvsc_core_046_not = ~input_a[16];
  assign popcount32_cvsc_core_048 = input_a[2] & input_a[22];
  assign popcount32_cvsc_core_049 = input_a[1] & input_a[16];
  assign popcount32_cvsc_core_052 = input_a[11] & input_a[0];
  assign popcount32_cvsc_core_053 = ~(input_a[26] & input_a[12]);
  assign popcount32_cvsc_core_056 = input_a[25] ^ input_a[19];
  assign popcount32_cvsc_core_057_not = ~input_a[26];
  assign popcount32_cvsc_core_058 = ~(input_a[7] & input_a[0]);
  assign popcount32_cvsc_core_059 = input_a[13] & input_a[13];
  assign popcount32_cvsc_core_060 = ~(input_a[3] ^ input_a[24]);
  assign popcount32_cvsc_core_061 = ~(input_a[16] | input_a[11]);
  assign popcount32_cvsc_core_062 = input_a[23] & input_a[11];
  assign popcount32_cvsc_core_063 = ~(input_a[30] ^ input_a[14]);
  assign popcount32_cvsc_core_068 = ~(input_a[6] ^ input_a[21]);
  assign popcount32_cvsc_core_069 = ~(input_a[14] & input_a[20]);
  assign popcount32_cvsc_core_070 = ~(input_a[22] & input_a[31]);
  assign popcount32_cvsc_core_071 = ~(input_a[29] ^ input_a[9]);
  assign popcount32_cvsc_core_073 = input_a[25] | input_a[6];
  assign popcount32_cvsc_core_075 = ~(input_a[19] & input_a[13]);
  assign popcount32_cvsc_core_076 = ~input_a[0];
  assign popcount32_cvsc_core_077 = input_a[27] | input_a[7];
  assign popcount32_cvsc_core_079 = ~input_a[15];
  assign popcount32_cvsc_core_081 = ~(input_a[10] | input_a[31]);
  assign popcount32_cvsc_core_082 = ~(input_a[15] ^ input_a[16]);
  assign popcount32_cvsc_core_083 = ~(input_a[23] & input_a[17]);
  assign popcount32_cvsc_core_084 = ~(input_a[25] | input_a[27]);
  assign popcount32_cvsc_core_085 = input_a[5] | input_a[4];
  assign popcount32_cvsc_core_086 = input_a[26] & input_a[17];
  assign popcount32_cvsc_core_087 = input_a[25] ^ input_a[26];
  assign popcount32_cvsc_core_090 = ~input_a[21];
  assign popcount32_cvsc_core_091 = input_a[31] | input_a[25];
  assign popcount32_cvsc_core_092 = ~input_a[13];
  assign popcount32_cvsc_core_093 = ~(input_a[30] ^ input_a[6]);
  assign popcount32_cvsc_core_095 = input_a[7] & input_a[2];
  assign popcount32_cvsc_core_096 = input_a[22] | input_a[23];
  assign popcount32_cvsc_core_098 = ~(input_a[0] ^ input_a[27]);
  assign popcount32_cvsc_core_099_not = ~input_a[25];
  assign popcount32_cvsc_core_100 = ~input_a[15];
  assign popcount32_cvsc_core_101 = ~(input_a[15] ^ input_a[18]);
  assign popcount32_cvsc_core_103 = ~(input_a[22] | input_a[5]);
  assign popcount32_cvsc_core_104 = ~input_a[2];
  assign popcount32_cvsc_core_105 = ~(input_a[25] | input_a[26]);
  assign popcount32_cvsc_core_107 = input_a[30] | input_a[4];
  assign popcount32_cvsc_core_108 = ~(input_a[19] & input_a[18]);
  assign popcount32_cvsc_core_109 = ~(input_a[28] | input_a[7]);
  assign popcount32_cvsc_core_110 = input_a[26] | input_a[11];
  assign popcount32_cvsc_core_112 = ~(input_a[6] & input_a[29]);
  assign popcount32_cvsc_core_113 = ~(input_a[12] & input_a[22]);
  assign popcount32_cvsc_core_114 = ~input_a[20];
  assign popcount32_cvsc_core_115 = input_a[29] & input_a[13];
  assign popcount32_cvsc_core_120 = ~(input_a[18] & input_a[9]);
  assign popcount32_cvsc_core_121 = input_a[12] & input_a[27];
  assign popcount32_cvsc_core_122 = input_a[7] | input_a[20];
  assign popcount32_cvsc_core_124 = input_a[15] ^ input_a[13];
  assign popcount32_cvsc_core_125 = input_a[10] ^ input_a[18];
  assign popcount32_cvsc_core_126 = ~(input_a[29] ^ input_a[29]);
  assign popcount32_cvsc_core_127 = ~(input_a[23] | input_a[8]);
  assign popcount32_cvsc_core_130 = ~(input_a[21] | input_a[15]);
  assign popcount32_cvsc_core_132 = ~input_a[23];
  assign popcount32_cvsc_core_133 = input_a[2] & input_a[11];
  assign popcount32_cvsc_core_134 = ~(input_a[26] ^ input_a[30]);
  assign popcount32_cvsc_core_136_not = ~input_a[3];
  assign popcount32_cvsc_core_138 = ~(input_a[20] ^ input_a[18]);
  assign popcount32_cvsc_core_139 = ~(input_a[1] & input_a[9]);
  assign popcount32_cvsc_core_141 = ~(input_a[10] | input_a[11]);
  assign popcount32_cvsc_core_142 = input_a[18] & input_a[20];
  assign popcount32_cvsc_core_144 = input_a[9] & input_a[22];
  assign popcount32_cvsc_core_145 = ~(input_a[12] ^ input_a[27]);
  assign popcount32_cvsc_core_147 = ~input_a[2];
  assign popcount32_cvsc_core_148 = input_a[21] & input_a[6];
  assign popcount32_cvsc_core_151 = ~input_a[7];
  assign popcount32_cvsc_core_152 = input_a[10] ^ input_a[29];
  assign popcount32_cvsc_core_155 = ~(input_a[4] & input_a[27]);
  assign popcount32_cvsc_core_156 = ~(input_a[15] & input_a[27]);
  assign popcount32_cvsc_core_159 = input_a[16] | input_a[3];
  assign popcount32_cvsc_core_166 = input_a[26] & input_a[8];
  assign popcount32_cvsc_core_167 = input_a[12] ^ input_a[0];
  assign popcount32_cvsc_core_168 = ~(input_a[25] | input_a[31]);
  assign popcount32_cvsc_core_169 = input_a[25] | input_a[15];
  assign popcount32_cvsc_core_171 = input_a[18] & input_a[3];
  assign popcount32_cvsc_core_172 = input_a[3] | input_a[19];
  assign popcount32_cvsc_core_173 = input_a[2] | input_a[31];
  assign popcount32_cvsc_core_174 = ~(input_a[27] & input_a[7]);
  assign popcount32_cvsc_core_175 = input_a[12] & input_a[26];
  assign popcount32_cvsc_core_179 = input_a[31] | input_a[6];
  assign popcount32_cvsc_core_180 = input_a[1] & input_a[30];
  assign popcount32_cvsc_core_181 = input_a[31] ^ input_a[15];
  assign popcount32_cvsc_core_182 = ~input_a[18];
  assign popcount32_cvsc_core_183 = input_a[14] | input_a[1];
  assign popcount32_cvsc_core_186 = input_a[29] | input_a[7];
  assign popcount32_cvsc_core_187 = input_a[2] | input_a[19];
  assign popcount32_cvsc_core_188 = ~(input_a[0] & input_a[24]);
  assign popcount32_cvsc_core_192 = input_a[16] & input_a[28];
  assign popcount32_cvsc_core_193 = ~(input_a[20] | input_a[8]);
  assign popcount32_cvsc_core_197 = ~(input_a[0] & input_a[30]);
  assign popcount32_cvsc_core_199 = ~(input_a[9] ^ input_a[18]);
  assign popcount32_cvsc_core_200 = input_a[3] & input_a[3];
  assign popcount32_cvsc_core_202 = input_a[16] ^ input_a[30];
  assign popcount32_cvsc_core_203 = ~input_a[3];
  assign popcount32_cvsc_core_204 = ~(input_a[24] | input_a[0]);
  assign popcount32_cvsc_core_205 = input_a[26] & input_a[7];
  assign popcount32_cvsc_core_206 = ~input_a[2];
  assign popcount32_cvsc_core_207 = input_a[21] & input_a[28];
  assign popcount32_cvsc_core_208 = input_a[14] ^ input_a[22];
  assign popcount32_cvsc_core_209 = input_a[2] | input_a[1];
  assign popcount32_cvsc_core_210 = input_a[26] ^ input_a[28];
  assign popcount32_cvsc_core_211 = ~(input_a[18] & input_a[9]);
  assign popcount32_cvsc_core_212 = ~(input_a[1] ^ input_a[19]);
  assign popcount32_cvsc_core_213 = input_a[21] | input_a[21];
  assign popcount32_cvsc_core_214 = input_a[8] & input_a[13];
  assign popcount32_cvsc_core_215 = ~(input_a[19] ^ input_a[9]);
  assign popcount32_cvsc_core_216 = ~(input_a[31] | input_a[7]);
  assign popcount32_cvsc_core_217 = ~(input_a[23] | input_a[7]);
  assign popcount32_cvsc_core_218 = input_a[16] | input_a[15];
  assign popcount32_cvsc_core_220 = ~(input_a[15] & input_a[26]);
  assign popcount32_cvsc_core_222 = ~input_a[14];
  assign popcount32_cvsc_core_223 = ~(input_a[19] & input_a[9]);
  assign popcount32_cvsc_core_224 = ~input_a[6];
  assign popcount32_cvsc_core_225 = ~(input_a[10] & input_a[20]);

  assign popcount32_cvsc_out[0] = 1'b0;
  assign popcount32_cvsc_out[1] = input_a[11];
  assign popcount32_cvsc_out[2] = input_a[6];
  assign popcount32_cvsc_out[3] = 1'b0;
  assign popcount32_cvsc_out[4] = 1'b0;
  assign popcount32_cvsc_out[5] = input_a[22];
endmodule