// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.09835
// WCE=12.0
// EP=0.851834%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_rb4r(input [20:0] input_a, output [4:0] popcount21_rb4r_out);
  wire popcount21_rb4r_core_025;
  wire popcount21_rb4r_core_026;
  wire popcount21_rb4r_core_027;
  wire popcount21_rb4r_core_028;
  wire popcount21_rb4r_core_029;
  wire popcount21_rb4r_core_032;
  wire popcount21_rb4r_core_033;
  wire popcount21_rb4r_core_034;
  wire popcount21_rb4r_core_035;
  wire popcount21_rb4r_core_036;
  wire popcount21_rb4r_core_037;
  wire popcount21_rb4r_core_039;
  wire popcount21_rb4r_core_043;
  wire popcount21_rb4r_core_044;
  wire popcount21_rb4r_core_045;
  wire popcount21_rb4r_core_046;
  wire popcount21_rb4r_core_047;
  wire popcount21_rb4r_core_048;
  wire popcount21_rb4r_core_049;
  wire popcount21_rb4r_core_050;
  wire popcount21_rb4r_core_051;
  wire popcount21_rb4r_core_053;
  wire popcount21_rb4r_core_054;
  wire popcount21_rb4r_core_055;
  wire popcount21_rb4r_core_056;
  wire popcount21_rb4r_core_057;
  wire popcount21_rb4r_core_058;
  wire popcount21_rb4r_core_059;
  wire popcount21_rb4r_core_061;
  wire popcount21_rb4r_core_063;
  wire popcount21_rb4r_core_064;
  wire popcount21_rb4r_core_065;
  wire popcount21_rb4r_core_066;
  wire popcount21_rb4r_core_067;
  wire popcount21_rb4r_core_070;
  wire popcount21_rb4r_core_072;
  wire popcount21_rb4r_core_073;
  wire popcount21_rb4r_core_076;
  wire popcount21_rb4r_core_077;
  wire popcount21_rb4r_core_078;
  wire popcount21_rb4r_core_080;
  wire popcount21_rb4r_core_081;
  wire popcount21_rb4r_core_082;
  wire popcount21_rb4r_core_084;
  wire popcount21_rb4r_core_086;
  wire popcount21_rb4r_core_087;
  wire popcount21_rb4r_core_088;
  wire popcount21_rb4r_core_089;
  wire popcount21_rb4r_core_091;
  wire popcount21_rb4r_core_092;
  wire popcount21_rb4r_core_094;
  wire popcount21_rb4r_core_095;
  wire popcount21_rb4r_core_097;
  wire popcount21_rb4r_core_098;
  wire popcount21_rb4r_core_099;
  wire popcount21_rb4r_core_100;
  wire popcount21_rb4r_core_105;
  wire popcount21_rb4r_core_106;
  wire popcount21_rb4r_core_107;
  wire popcount21_rb4r_core_108;
  wire popcount21_rb4r_core_109;
  wire popcount21_rb4r_core_111;
  wire popcount21_rb4r_core_113;
  wire popcount21_rb4r_core_114;
  wire popcount21_rb4r_core_115;
  wire popcount21_rb4r_core_117;
  wire popcount21_rb4r_core_118_not;
  wire popcount21_rb4r_core_119;
  wire popcount21_rb4r_core_121_not;
  wire popcount21_rb4r_core_122_not;
  wire popcount21_rb4r_core_124;
  wire popcount21_rb4r_core_125;
  wire popcount21_rb4r_core_127;
  wire popcount21_rb4r_core_129;
  wire popcount21_rb4r_core_130_not;
  wire popcount21_rb4r_core_131;
  wire popcount21_rb4r_core_133;
  wire popcount21_rb4r_core_134;
  wire popcount21_rb4r_core_136;
  wire popcount21_rb4r_core_139;
  wire popcount21_rb4r_core_140;
  wire popcount21_rb4r_core_141;
  wire popcount21_rb4r_core_143;
  wire popcount21_rb4r_core_145;
  wire popcount21_rb4r_core_146;
  wire popcount21_rb4r_core_147;
  wire popcount21_rb4r_core_149;
  wire popcount21_rb4r_core_151;
  wire popcount21_rb4r_core_152;
  wire popcount21_rb4r_core_153;

  assign popcount21_rb4r_core_025 = input_a[7] | input_a[9];
  assign popcount21_rb4r_core_026 = ~input_a[3];
  assign popcount21_rb4r_core_027 = input_a[1] | input_a[14];
  assign popcount21_rb4r_core_028 = input_a[7] & input_a[10];
  assign popcount21_rb4r_core_029 = ~(input_a[18] ^ input_a[9]);
  assign popcount21_rb4r_core_032 = ~(input_a[14] ^ input_a[7]);
  assign popcount21_rb4r_core_033 = ~(input_a[14] ^ input_a[13]);
  assign popcount21_rb4r_core_034 = input_a[5] ^ input_a[6];
  assign popcount21_rb4r_core_035 = ~input_a[7];
  assign popcount21_rb4r_core_036 = input_a[3] & input_a[16];
  assign popcount21_rb4r_core_037 = ~(input_a[3] ^ input_a[6]);
  assign popcount21_rb4r_core_039 = ~input_a[20];
  assign popcount21_rb4r_core_043 = input_a[20] | input_a[20];
  assign popcount21_rb4r_core_044 = input_a[13] | input_a[12];
  assign popcount21_rb4r_core_045 = ~input_a[6];
  assign popcount21_rb4r_core_046 = input_a[13] & input_a[19];
  assign popcount21_rb4r_core_047 = ~input_a[20];
  assign popcount21_rb4r_core_048 = ~input_a[2];
  assign popcount21_rb4r_core_049 = input_a[17] & input_a[7];
  assign popcount21_rb4r_core_050 = ~(input_a[3] & input_a[20]);
  assign popcount21_rb4r_core_051 = input_a[7] | input_a[8];
  assign popcount21_rb4r_core_053 = ~(input_a[14] ^ input_a[5]);
  assign popcount21_rb4r_core_054 = ~(input_a[20] ^ input_a[13]);
  assign popcount21_rb4r_core_055 = input_a[15] | input_a[14];
  assign popcount21_rb4r_core_056 = ~input_a[17];
  assign popcount21_rb4r_core_057 = ~(input_a[15] | input_a[6]);
  assign popcount21_rb4r_core_058 = ~(input_a[18] & input_a[7]);
  assign popcount21_rb4r_core_059 = ~(input_a[11] & input_a[4]);
  assign popcount21_rb4r_core_061 = input_a[20] | input_a[0];
  assign popcount21_rb4r_core_063 = ~(input_a[16] & input_a[11]);
  assign popcount21_rb4r_core_064 = input_a[11] | input_a[7];
  assign popcount21_rb4r_core_065 = ~(input_a[4] | input_a[0]);
  assign popcount21_rb4r_core_066 = ~(input_a[8] ^ input_a[14]);
  assign popcount21_rb4r_core_067 = ~(input_a[19] & input_a[7]);
  assign popcount21_rb4r_core_070 = input_a[20] & input_a[15];
  assign popcount21_rb4r_core_072 = input_a[20] & input_a[19];
  assign popcount21_rb4r_core_073 = ~(input_a[2] ^ input_a[14]);
  assign popcount21_rb4r_core_076 = input_a[12] ^ input_a[9];
  assign popcount21_rb4r_core_077 = input_a[3] | input_a[5];
  assign popcount21_rb4r_core_078 = input_a[15] | input_a[0];
  assign popcount21_rb4r_core_080 = ~(input_a[12] | input_a[11]);
  assign popcount21_rb4r_core_081 = input_a[15] | input_a[20];
  assign popcount21_rb4r_core_082 = input_a[5] ^ input_a[18];
  assign popcount21_rb4r_core_084 = ~(input_a[15] ^ input_a[9]);
  assign popcount21_rb4r_core_086 = ~(input_a[4] ^ input_a[14]);
  assign popcount21_rb4r_core_087 = input_a[14] & input_a[17];
  assign popcount21_rb4r_core_088 = ~(input_a[17] & input_a[17]);
  assign popcount21_rb4r_core_089 = ~input_a[0];
  assign popcount21_rb4r_core_091 = ~input_a[3];
  assign popcount21_rb4r_core_092 = input_a[11] | input_a[4];
  assign popcount21_rb4r_core_094 = input_a[15] ^ input_a[8];
  assign popcount21_rb4r_core_095 = ~(input_a[9] & input_a[3]);
  assign popcount21_rb4r_core_097 = ~input_a[13];
  assign popcount21_rb4r_core_098 = input_a[7] & input_a[16];
  assign popcount21_rb4r_core_099 = input_a[14] & input_a[7];
  assign popcount21_rb4r_core_100 = ~input_a[3];
  assign popcount21_rb4r_core_105 = input_a[16] | input_a[12];
  assign popcount21_rb4r_core_106 = ~(input_a[15] & input_a[6]);
  assign popcount21_rb4r_core_107 = input_a[15] | input_a[15];
  assign popcount21_rb4r_core_108 = ~(input_a[15] & input_a[15]);
  assign popcount21_rb4r_core_109 = input_a[6] ^ input_a[20];
  assign popcount21_rb4r_core_111 = ~input_a[7];
  assign popcount21_rb4r_core_113 = input_a[6] | input_a[5];
  assign popcount21_rb4r_core_114 = ~(input_a[3] ^ input_a[13]);
  assign popcount21_rb4r_core_115 = ~(input_a[1] & input_a[18]);
  assign popcount21_rb4r_core_117 = ~(input_a[2] | input_a[10]);
  assign popcount21_rb4r_core_118_not = ~input_a[5];
  assign popcount21_rb4r_core_119 = input_a[3] | input_a[2];
  assign popcount21_rb4r_core_121_not = ~input_a[11];
  assign popcount21_rb4r_core_122_not = ~input_a[4];
  assign popcount21_rb4r_core_124 = ~(input_a[14] ^ input_a[5]);
  assign popcount21_rb4r_core_125 = input_a[13] & input_a[12];
  assign popcount21_rb4r_core_127 = ~(input_a[3] | input_a[14]);
  assign popcount21_rb4r_core_129 = ~(input_a[11] | input_a[0]);
  assign popcount21_rb4r_core_130_not = ~input_a[16];
  assign popcount21_rb4r_core_131 = ~input_a[7];
  assign popcount21_rb4r_core_133 = ~(input_a[8] ^ input_a[2]);
  assign popcount21_rb4r_core_134 = input_a[11] & input_a[3];
  assign popcount21_rb4r_core_136 = ~(input_a[5] ^ input_a[19]);
  assign popcount21_rb4r_core_139 = ~input_a[13];
  assign popcount21_rb4r_core_140 = input_a[17] | input_a[12];
  assign popcount21_rb4r_core_141 = input_a[3] | input_a[11];
  assign popcount21_rb4r_core_143 = ~input_a[1];
  assign popcount21_rb4r_core_145 = input_a[12] | input_a[10];
  assign popcount21_rb4r_core_146 = ~(input_a[9] ^ input_a[16]);
  assign popcount21_rb4r_core_147 = ~(input_a[4] | input_a[20]);
  assign popcount21_rb4r_core_149 = input_a[16] | input_a[2];
  assign popcount21_rb4r_core_151 = input_a[19] | input_a[4];
  assign popcount21_rb4r_core_152 = input_a[16] ^ input_a[11];
  assign popcount21_rb4r_core_153 = ~input_a[4];

  assign popcount21_rb4r_out[0] = input_a[8];
  assign popcount21_rb4r_out[1] = 1'b1;
  assign popcount21_rb4r_out[2] = 1'b0;
  assign popcount21_rb4r_out[3] = 1'b1;
  assign popcount21_rb4r_out[4] = 1'b0;
endmodule