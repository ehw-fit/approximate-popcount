// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.56096
// WCE=28.0
// EP=0.98188%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_8ly7(input [30:0] input_a, output [4:0] popcount31_8ly7_out);
  wire popcount31_8ly7_core_034;
  wire popcount31_8ly7_core_037_not;
  wire popcount31_8ly7_core_038;
  wire popcount31_8ly7_core_039;
  wire popcount31_8ly7_core_040;
  wire popcount31_8ly7_core_041;
  wire popcount31_8ly7_core_042;
  wire popcount31_8ly7_core_044;
  wire popcount31_8ly7_core_045;
  wire popcount31_8ly7_core_047;
  wire popcount31_8ly7_core_049;
  wire popcount31_8ly7_core_050;
  wire popcount31_8ly7_core_052;
  wire popcount31_8ly7_core_054_not;
  wire popcount31_8ly7_core_055;
  wire popcount31_8ly7_core_056;
  wire popcount31_8ly7_core_057;
  wire popcount31_8ly7_core_058;
  wire popcount31_8ly7_core_059;
  wire popcount31_8ly7_core_060;
  wire popcount31_8ly7_core_061;
  wire popcount31_8ly7_core_062;
  wire popcount31_8ly7_core_063;
  wire popcount31_8ly7_core_068;
  wire popcount31_8ly7_core_069;
  wire popcount31_8ly7_core_071;
  wire popcount31_8ly7_core_072;
  wire popcount31_8ly7_core_075;
  wire popcount31_8ly7_core_077;
  wire popcount31_8ly7_core_079;
  wire popcount31_8ly7_core_081;
  wire popcount31_8ly7_core_082;
  wire popcount31_8ly7_core_083;
  wire popcount31_8ly7_core_086;
  wire popcount31_8ly7_core_087;
  wire popcount31_8ly7_core_088;
  wire popcount31_8ly7_core_089;
  wire popcount31_8ly7_core_090;
  wire popcount31_8ly7_core_092;
  wire popcount31_8ly7_core_094_not;
  wire popcount31_8ly7_core_095;
  wire popcount31_8ly7_core_096;
  wire popcount31_8ly7_core_097;
  wire popcount31_8ly7_core_099;
  wire popcount31_8ly7_core_101;
  wire popcount31_8ly7_core_102;
  wire popcount31_8ly7_core_104;
  wire popcount31_8ly7_core_105;
  wire popcount31_8ly7_core_106;
  wire popcount31_8ly7_core_107;
  wire popcount31_8ly7_core_108;
  wire popcount31_8ly7_core_109;
  wire popcount31_8ly7_core_111;
  wire popcount31_8ly7_core_112;
  wire popcount31_8ly7_core_113;
  wire popcount31_8ly7_core_114;
  wire popcount31_8ly7_core_115;
  wire popcount31_8ly7_core_118;
  wire popcount31_8ly7_core_119;
  wire popcount31_8ly7_core_121;
  wire popcount31_8ly7_core_123;
  wire popcount31_8ly7_core_124;
  wire popcount31_8ly7_core_127;
  wire popcount31_8ly7_core_128;
  wire popcount31_8ly7_core_131;
  wire popcount31_8ly7_core_132;
  wire popcount31_8ly7_core_133;
  wire popcount31_8ly7_core_134;
  wire popcount31_8ly7_core_135;
  wire popcount31_8ly7_core_136_not;
  wire popcount31_8ly7_core_137;
  wire popcount31_8ly7_core_138;
  wire popcount31_8ly7_core_141;
  wire popcount31_8ly7_core_142;
  wire popcount31_8ly7_core_143;
  wire popcount31_8ly7_core_144;
  wire popcount31_8ly7_core_145;
  wire popcount31_8ly7_core_146;
  wire popcount31_8ly7_core_147;
  wire popcount31_8ly7_core_148;
  wire popcount31_8ly7_core_149;
  wire popcount31_8ly7_core_150;
  wire popcount31_8ly7_core_151;
  wire popcount31_8ly7_core_152;
  wire popcount31_8ly7_core_154;
  wire popcount31_8ly7_core_155;
  wire popcount31_8ly7_core_156;
  wire popcount31_8ly7_core_158;
  wire popcount31_8ly7_core_159_not;
  wire popcount31_8ly7_core_160;
  wire popcount31_8ly7_core_162;
  wire popcount31_8ly7_core_165;
  wire popcount31_8ly7_core_166;
  wire popcount31_8ly7_core_167;
  wire popcount31_8ly7_core_168;
  wire popcount31_8ly7_core_169;
  wire popcount31_8ly7_core_170;
  wire popcount31_8ly7_core_174;
  wire popcount31_8ly7_core_175;
  wire popcount31_8ly7_core_177;
  wire popcount31_8ly7_core_179;
  wire popcount31_8ly7_core_182;
  wire popcount31_8ly7_core_184;
  wire popcount31_8ly7_core_185;
  wire popcount31_8ly7_core_186;
  wire popcount31_8ly7_core_187;
  wire popcount31_8ly7_core_189;
  wire popcount31_8ly7_core_191;
  wire popcount31_8ly7_core_192;
  wire popcount31_8ly7_core_193;
  wire popcount31_8ly7_core_195;
  wire popcount31_8ly7_core_196;
  wire popcount31_8ly7_core_197;
  wire popcount31_8ly7_core_198;
  wire popcount31_8ly7_core_199;
  wire popcount31_8ly7_core_200;
  wire popcount31_8ly7_core_201;
  wire popcount31_8ly7_core_202;
  wire popcount31_8ly7_core_203;
  wire popcount31_8ly7_core_204;
  wire popcount31_8ly7_core_205;
  wire popcount31_8ly7_core_207;
  wire popcount31_8ly7_core_208;
  wire popcount31_8ly7_core_209;
  wire popcount31_8ly7_core_210;
  wire popcount31_8ly7_core_211;
  wire popcount31_8ly7_core_215;
  wire popcount31_8ly7_core_217;
  wire popcount31_8ly7_core_218;
  wire popcount31_8ly7_core_219;

  assign popcount31_8ly7_core_034 = input_a[16] | input_a[1];
  assign popcount31_8ly7_core_037_not = ~input_a[3];
  assign popcount31_8ly7_core_038 = ~(input_a[22] | input_a[4]);
  assign popcount31_8ly7_core_039 = ~(input_a[1] | input_a[4]);
  assign popcount31_8ly7_core_040 = ~(input_a[18] ^ input_a[9]);
  assign popcount31_8ly7_core_041 = input_a[17] ^ input_a[7];
  assign popcount31_8ly7_core_042 = ~(input_a[22] | input_a[13]);
  assign popcount31_8ly7_core_044 = ~(input_a[10] & input_a[20]);
  assign popcount31_8ly7_core_045 = ~(input_a[6] ^ input_a[21]);
  assign popcount31_8ly7_core_047 = ~(input_a[3] | input_a[25]);
  assign popcount31_8ly7_core_049 = ~(input_a[27] & input_a[29]);
  assign popcount31_8ly7_core_050 = input_a[13] & input_a[15];
  assign popcount31_8ly7_core_052 = ~input_a[24];
  assign popcount31_8ly7_core_054_not = ~input_a[17];
  assign popcount31_8ly7_core_055 = input_a[0] & input_a[0];
  assign popcount31_8ly7_core_056 = input_a[30] | input_a[7];
  assign popcount31_8ly7_core_057 = ~(input_a[13] ^ input_a[10]);
  assign popcount31_8ly7_core_058 = ~input_a[5];
  assign popcount31_8ly7_core_059 = input_a[4] ^ input_a[14];
  assign popcount31_8ly7_core_060 = input_a[26] | input_a[15];
  assign popcount31_8ly7_core_061 = input_a[17] | input_a[22];
  assign popcount31_8ly7_core_062 = ~(input_a[6] & input_a[2]);
  assign popcount31_8ly7_core_063 = ~input_a[5];
  assign popcount31_8ly7_core_068 = input_a[23] ^ input_a[18];
  assign popcount31_8ly7_core_069 = input_a[8] ^ input_a[19];
  assign popcount31_8ly7_core_071 = ~(input_a[26] | input_a[30]);
  assign popcount31_8ly7_core_072 = ~(input_a[8] | input_a[23]);
  assign popcount31_8ly7_core_075 = input_a[24] & input_a[9];
  assign popcount31_8ly7_core_077 = input_a[7] | input_a[25];
  assign popcount31_8ly7_core_079 = ~(input_a[17] & input_a[10]);
  assign popcount31_8ly7_core_081 = input_a[12] ^ input_a[1];
  assign popcount31_8ly7_core_082 = ~(input_a[16] & input_a[8]);
  assign popcount31_8ly7_core_083 = input_a[22] ^ input_a[6];
  assign popcount31_8ly7_core_086 = input_a[27] ^ input_a[13];
  assign popcount31_8ly7_core_087 = ~(input_a[9] | input_a[17]);
  assign popcount31_8ly7_core_088 = input_a[26] & input_a[26];
  assign popcount31_8ly7_core_089 = ~input_a[1];
  assign popcount31_8ly7_core_090 = ~(input_a[5] ^ input_a[8]);
  assign popcount31_8ly7_core_092 = input_a[4] & input_a[29];
  assign popcount31_8ly7_core_094_not = ~input_a[5];
  assign popcount31_8ly7_core_095 = ~input_a[5];
  assign popcount31_8ly7_core_096 = input_a[0] ^ input_a[1];
  assign popcount31_8ly7_core_097 = ~(input_a[21] & input_a[29]);
  assign popcount31_8ly7_core_099 = input_a[12] ^ input_a[1];
  assign popcount31_8ly7_core_101 = ~input_a[10];
  assign popcount31_8ly7_core_102 = input_a[26] ^ input_a[0];
  assign popcount31_8ly7_core_104 = ~input_a[2];
  assign popcount31_8ly7_core_105 = ~input_a[11];
  assign popcount31_8ly7_core_106 = input_a[1] | input_a[6];
  assign popcount31_8ly7_core_107 = ~(input_a[23] | input_a[6]);
  assign popcount31_8ly7_core_108 = ~(input_a[25] | input_a[10]);
  assign popcount31_8ly7_core_109 = input_a[23] ^ input_a[8];
  assign popcount31_8ly7_core_111 = ~(input_a[30] & input_a[20]);
  assign popcount31_8ly7_core_112 = input_a[26] ^ input_a[8];
  assign popcount31_8ly7_core_113 = input_a[9] & input_a[6];
  assign popcount31_8ly7_core_114 = input_a[14] & input_a[9];
  assign popcount31_8ly7_core_115 = ~(input_a[11] & input_a[27]);
  assign popcount31_8ly7_core_118 = input_a[10] | input_a[8];
  assign popcount31_8ly7_core_119 = ~(input_a[26] & input_a[5]);
  assign popcount31_8ly7_core_121 = ~input_a[13];
  assign popcount31_8ly7_core_123 = ~(input_a[15] | input_a[10]);
  assign popcount31_8ly7_core_124 = ~(input_a[20] ^ input_a[2]);
  assign popcount31_8ly7_core_127 = ~(input_a[14] ^ input_a[2]);
  assign popcount31_8ly7_core_128 = ~(input_a[1] ^ input_a[1]);
  assign popcount31_8ly7_core_131 = input_a[17] ^ input_a[22];
  assign popcount31_8ly7_core_132 = ~(input_a[13] ^ input_a[18]);
  assign popcount31_8ly7_core_133 = ~input_a[19];
  assign popcount31_8ly7_core_134 = ~input_a[29];
  assign popcount31_8ly7_core_135 = input_a[0] | input_a[24];
  assign popcount31_8ly7_core_136_not = ~input_a[20];
  assign popcount31_8ly7_core_137 = input_a[26] ^ input_a[0];
  assign popcount31_8ly7_core_138 = ~(input_a[26] ^ input_a[19]);
  assign popcount31_8ly7_core_141 = ~(input_a[15] | input_a[15]);
  assign popcount31_8ly7_core_142 = ~input_a[19];
  assign popcount31_8ly7_core_143 = input_a[19] & input_a[1];
  assign popcount31_8ly7_core_144 = ~(input_a[28] | input_a[8]);
  assign popcount31_8ly7_core_145 = ~input_a[17];
  assign popcount31_8ly7_core_146 = ~(input_a[30] & input_a[28]);
  assign popcount31_8ly7_core_147 = input_a[4] ^ input_a[18];
  assign popcount31_8ly7_core_148 = ~(input_a[10] ^ input_a[18]);
  assign popcount31_8ly7_core_149 = input_a[17] & input_a[9];
  assign popcount31_8ly7_core_150 = ~input_a[23];
  assign popcount31_8ly7_core_151 = ~(input_a[18] | input_a[20]);
  assign popcount31_8ly7_core_152 = input_a[15] & input_a[11];
  assign popcount31_8ly7_core_154 = ~(input_a[18] | input_a[10]);
  assign popcount31_8ly7_core_155 = ~(input_a[24] ^ input_a[13]);
  assign popcount31_8ly7_core_156 = ~(input_a[26] & input_a[0]);
  assign popcount31_8ly7_core_158 = input_a[13] ^ input_a[1];
  assign popcount31_8ly7_core_159_not = ~input_a[6];
  assign popcount31_8ly7_core_160 = input_a[7] & input_a[25];
  assign popcount31_8ly7_core_162 = ~(input_a[3] & input_a[5]);
  assign popcount31_8ly7_core_165 = input_a[24] | input_a[11];
  assign popcount31_8ly7_core_166 = ~(input_a[19] & input_a[4]);
  assign popcount31_8ly7_core_167 = input_a[20] | input_a[20];
  assign popcount31_8ly7_core_168 = input_a[25] ^ input_a[27];
  assign popcount31_8ly7_core_169 = ~input_a[19];
  assign popcount31_8ly7_core_170 = input_a[21] | input_a[15];
  assign popcount31_8ly7_core_174 = input_a[13] ^ input_a[16];
  assign popcount31_8ly7_core_175 = ~(input_a[28] & input_a[10]);
  assign popcount31_8ly7_core_177 = ~(input_a[2] & input_a[11]);
  assign popcount31_8ly7_core_179 = ~(input_a[21] & input_a[20]);
  assign popcount31_8ly7_core_182 = ~(input_a[2] & input_a[9]);
  assign popcount31_8ly7_core_184 = ~(input_a[9] | input_a[30]);
  assign popcount31_8ly7_core_185 = ~(input_a[12] ^ input_a[20]);
  assign popcount31_8ly7_core_186 = ~(input_a[20] | input_a[20]);
  assign popcount31_8ly7_core_187 = ~(input_a[21] | input_a[29]);
  assign popcount31_8ly7_core_189 = ~(input_a[17] ^ input_a[3]);
  assign popcount31_8ly7_core_191 = ~(input_a[17] | input_a[27]);
  assign popcount31_8ly7_core_192 = ~input_a[21];
  assign popcount31_8ly7_core_193 = ~input_a[28];
  assign popcount31_8ly7_core_195 = ~input_a[9];
  assign popcount31_8ly7_core_196 = ~(input_a[25] | input_a[18]);
  assign popcount31_8ly7_core_197 = ~(input_a[19] ^ input_a[21]);
  assign popcount31_8ly7_core_198 = input_a[4] | input_a[8];
  assign popcount31_8ly7_core_199 = input_a[16] ^ input_a[28];
  assign popcount31_8ly7_core_200 = ~(input_a[20] | input_a[29]);
  assign popcount31_8ly7_core_201 = input_a[20] ^ input_a[25];
  assign popcount31_8ly7_core_202 = ~input_a[6];
  assign popcount31_8ly7_core_203 = input_a[24] | input_a[2];
  assign popcount31_8ly7_core_204 = ~(input_a[27] & input_a[13]);
  assign popcount31_8ly7_core_205 = input_a[22] ^ input_a[4];
  assign popcount31_8ly7_core_207 = input_a[16] | input_a[17];
  assign popcount31_8ly7_core_208 = input_a[14] ^ input_a[4];
  assign popcount31_8ly7_core_209 = ~input_a[10];
  assign popcount31_8ly7_core_210 = ~(input_a[13] ^ input_a[9]);
  assign popcount31_8ly7_core_211 = input_a[29] & input_a[17];
  assign popcount31_8ly7_core_215 = ~(input_a[29] | input_a[10]);
  assign popcount31_8ly7_core_217 = ~(input_a[0] & input_a[22]);
  assign popcount31_8ly7_core_218 = input_a[30] | input_a[4];
  assign popcount31_8ly7_core_219 = ~(input_a[5] & input_a[10]);

  assign popcount31_8ly7_out[0] = 1'b1;
  assign popcount31_8ly7_out[1] = 1'b0;
  assign popcount31_8ly7_out[2] = input_a[10];
  assign popcount31_8ly7_out[3] = input_a[11];
  assign popcount31_8ly7_out[4] = 1'b0;
endmodule