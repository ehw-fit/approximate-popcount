// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.97587
// WCE=23.0
// EP=0.894228%
// Printed PDK parameters:
//  Area=17247315.0
//  Delay=44464396.0
//  Power=799580.0

module popcount45_0xd7(input [44:0] input_a, output [5:0] popcount45_0xd7_out);
  wire popcount45_0xd7_core_047;
  wire popcount45_0xd7_core_048;
  wire popcount45_0xd7_core_049;
  wire popcount45_0xd7_core_050;
  wire popcount45_0xd7_core_051;
  wire popcount45_0xd7_core_052;
  wire popcount45_0xd7_core_054;
  wire popcount45_0xd7_core_056;
  wire popcount45_0xd7_core_057;
  wire popcount45_0xd7_core_058;
  wire popcount45_0xd7_core_059;
  wire popcount45_0xd7_core_060;
  wire popcount45_0xd7_core_061;
  wire popcount45_0xd7_core_062;
  wire popcount45_0xd7_core_063;
  wire popcount45_0xd7_core_068;
  wire popcount45_0xd7_core_069;
  wire popcount45_0xd7_core_070;
  wire popcount45_0xd7_core_072;
  wire popcount45_0xd7_core_073;
  wire popcount45_0xd7_core_074;
  wire popcount45_0xd7_core_075_not;
  wire popcount45_0xd7_core_076;
  wire popcount45_0xd7_core_077;
  wire popcount45_0xd7_core_079;
  wire popcount45_0xd7_core_081;
  wire popcount45_0xd7_core_084;
  wire popcount45_0xd7_core_086;
  wire popcount45_0xd7_core_087;
  wire popcount45_0xd7_core_089;
  wire popcount45_0xd7_core_090;
  wire popcount45_0xd7_core_093;
  wire popcount45_0xd7_core_094_not;
  wire popcount45_0xd7_core_095;
  wire popcount45_0xd7_core_099;
  wire popcount45_0xd7_core_100;
  wire popcount45_0xd7_core_101;
  wire popcount45_0xd7_core_104;
  wire popcount45_0xd7_core_105;
  wire popcount45_0xd7_core_106;
  wire popcount45_0xd7_core_107;
  wire popcount45_0xd7_core_109;
  wire popcount45_0xd7_core_110;
  wire popcount45_0xd7_core_114;
  wire popcount45_0xd7_core_117;
  wire popcount45_0xd7_core_118;
  wire popcount45_0xd7_core_121;
  wire popcount45_0xd7_core_122;
  wire popcount45_0xd7_core_123;
  wire popcount45_0xd7_core_124;
  wire popcount45_0xd7_core_125;
  wire popcount45_0xd7_core_126;
  wire popcount45_0xd7_core_127;
  wire popcount45_0xd7_core_128;
  wire popcount45_0xd7_core_130;
  wire popcount45_0xd7_core_131;
  wire popcount45_0xd7_core_132;
  wire popcount45_0xd7_core_133;
  wire popcount45_0xd7_core_134;
  wire popcount45_0xd7_core_136;
  wire popcount45_0xd7_core_137;
  wire popcount45_0xd7_core_139;
  wire popcount45_0xd7_core_140;
  wire popcount45_0xd7_core_141;
  wire popcount45_0xd7_core_142;
  wire popcount45_0xd7_core_143;
  wire popcount45_0xd7_core_145;
  wire popcount45_0xd7_core_147;
  wire popcount45_0xd7_core_149;
  wire popcount45_0xd7_core_150;
  wire popcount45_0xd7_core_151;
  wire popcount45_0xd7_core_153;
  wire popcount45_0xd7_core_154;
  wire popcount45_0xd7_core_155;
  wire popcount45_0xd7_core_156;
  wire popcount45_0xd7_core_157;
  wire popcount45_0xd7_core_159;
  wire popcount45_0xd7_core_167;
  wire popcount45_0xd7_core_168;
  wire popcount45_0xd7_core_170;
  wire popcount45_0xd7_core_171;
  wire popcount45_0xd7_core_172;
  wire popcount45_0xd7_core_173;
  wire popcount45_0xd7_core_174;
  wire popcount45_0xd7_core_177;
  wire popcount45_0xd7_core_178;
  wire popcount45_0xd7_core_181;
  wire popcount45_0xd7_core_185;
  wire popcount45_0xd7_core_191;
  wire popcount45_0xd7_core_194;
  wire popcount45_0xd7_core_195;
  wire popcount45_0xd7_core_196;
  wire popcount45_0xd7_core_200;
  wire popcount45_0xd7_core_201;
  wire popcount45_0xd7_core_202;
  wire popcount45_0xd7_core_206;
  wire popcount45_0xd7_core_207;
  wire popcount45_0xd7_core_208;
  wire popcount45_0xd7_core_209;
  wire popcount45_0xd7_core_210;
  wire popcount45_0xd7_core_211;
  wire popcount45_0xd7_core_213;
  wire popcount45_0xd7_core_216;
  wire popcount45_0xd7_core_220;
  wire popcount45_0xd7_core_221;
  wire popcount45_0xd7_core_224;
  wire popcount45_0xd7_core_228;
  wire popcount45_0xd7_core_229;
  wire popcount45_0xd7_core_231;
  wire popcount45_0xd7_core_234;
  wire popcount45_0xd7_core_240;
  wire popcount45_0xd7_core_241;
  wire popcount45_0xd7_core_249;
  wire popcount45_0xd7_core_250;
  wire popcount45_0xd7_core_252;
  wire popcount45_0xd7_core_253;
  wire popcount45_0xd7_core_254;
  wire popcount45_0xd7_core_255;
  wire popcount45_0xd7_core_257;
  wire popcount45_0xd7_core_258;
  wire popcount45_0xd7_core_259;
  wire popcount45_0xd7_core_260;
  wire popcount45_0xd7_core_263;
  wire popcount45_0xd7_core_265;
  wire popcount45_0xd7_core_266;
  wire popcount45_0xd7_core_267_not;
  wire popcount45_0xd7_core_268;
  wire popcount45_0xd7_core_269;
  wire popcount45_0xd7_core_271;
  wire popcount45_0xd7_core_275;
  wire popcount45_0xd7_core_277;
  wire popcount45_0xd7_core_278;
  wire popcount45_0xd7_core_281;
  wire popcount45_0xd7_core_282;
  wire popcount45_0xd7_core_283;
  wire popcount45_0xd7_core_284;
  wire popcount45_0xd7_core_286;
  wire popcount45_0xd7_core_287;
  wire popcount45_0xd7_core_288_not;
  wire popcount45_0xd7_core_289;
  wire popcount45_0xd7_core_290;
  wire popcount45_0xd7_core_291;
  wire popcount45_0xd7_core_292;
  wire popcount45_0xd7_core_293;
  wire popcount45_0xd7_core_294;
  wire popcount45_0xd7_core_295;
  wire popcount45_0xd7_core_298;
  wire popcount45_0xd7_core_299;
  wire popcount45_0xd7_core_300;
  wire popcount45_0xd7_core_301;
  wire popcount45_0xd7_core_302;
  wire popcount45_0xd7_core_303;
  wire popcount45_0xd7_core_305;
  wire popcount45_0xd7_core_306;
  wire popcount45_0xd7_core_309;
  wire popcount45_0xd7_core_310;
  wire popcount45_0xd7_core_312;
  wire popcount45_0xd7_core_316;
  wire popcount45_0xd7_core_318;
  wire popcount45_0xd7_core_319;
  wire popcount45_0xd7_core_320;
  wire popcount45_0xd7_core_321;
  wire popcount45_0xd7_core_323;
  wire popcount45_0xd7_core_324;
  wire popcount45_0xd7_core_326;
  wire popcount45_0xd7_core_327;
  wire popcount45_0xd7_core_328;
  wire popcount45_0xd7_core_329;
  wire popcount45_0xd7_core_330;
  wire popcount45_0xd7_core_332;
  wire popcount45_0xd7_core_333;
  wire popcount45_0xd7_core_336;
  wire popcount45_0xd7_core_337;
  wire popcount45_0xd7_core_338;
  wire popcount45_0xd7_core_342;
  wire popcount45_0xd7_core_344;
  wire popcount45_0xd7_core_345;
  wire popcount45_0xd7_core_346;
  wire popcount45_0xd7_core_347;
  wire popcount45_0xd7_core_348;
  wire popcount45_0xd7_core_349;
  wire popcount45_0xd7_core_350;
  wire popcount45_0xd7_core_351;
  wire popcount45_0xd7_core_352;
  wire popcount45_0xd7_core_353;
  wire popcount45_0xd7_core_354;
  wire popcount45_0xd7_core_355;
  wire popcount45_0xd7_core_356;

  assign popcount45_0xd7_core_047 = input_a[13] | input_a[31];
  assign popcount45_0xd7_core_048 = ~(input_a[11] ^ input_a[34]);
  assign popcount45_0xd7_core_049 = input_a[8] ^ input_a[41];
  assign popcount45_0xd7_core_050 = ~input_a[22];
  assign popcount45_0xd7_core_051 = input_a[1] ^ input_a[16];
  assign popcount45_0xd7_core_052 = input_a[25] | input_a[10];
  assign popcount45_0xd7_core_054 = input_a[37] | input_a[18];
  assign popcount45_0xd7_core_056 = input_a[1] | input_a[31];
  assign popcount45_0xd7_core_057 = input_a[12] ^ input_a[18];
  assign popcount45_0xd7_core_058 = input_a[22] ^ input_a[32];
  assign popcount45_0xd7_core_059 = input_a[36] ^ input_a[44];
  assign popcount45_0xd7_core_060 = ~(input_a[42] | input_a[13]);
  assign popcount45_0xd7_core_061 = input_a[11] ^ input_a[37];
  assign popcount45_0xd7_core_062 = ~(input_a[41] ^ input_a[31]);
  assign popcount45_0xd7_core_063 = ~(input_a[35] ^ input_a[14]);
  assign popcount45_0xd7_core_068 = ~(input_a[29] & input_a[22]);
  assign popcount45_0xd7_core_069 = input_a[27] ^ input_a[25];
  assign popcount45_0xd7_core_070 = input_a[35] & input_a[26];
  assign popcount45_0xd7_core_072 = input_a[33] ^ input_a[40];
  assign popcount45_0xd7_core_073 = input_a[36] ^ input_a[44];
  assign popcount45_0xd7_core_074 = ~(input_a[32] ^ input_a[31]);
  assign popcount45_0xd7_core_075_not = ~input_a[25];
  assign popcount45_0xd7_core_076 = input_a[21] & input_a[11];
  assign popcount45_0xd7_core_077 = input_a[20] & input_a[26];
  assign popcount45_0xd7_core_079 = ~(input_a[36] & input_a[6]);
  assign popcount45_0xd7_core_081 = ~(input_a[12] & input_a[20]);
  assign popcount45_0xd7_core_084 = ~(input_a[17] | input_a[3]);
  assign popcount45_0xd7_core_086 = input_a[19] ^ input_a[3];
  assign popcount45_0xd7_core_087 = ~(input_a[11] ^ input_a[12]);
  assign popcount45_0xd7_core_089 = ~(input_a[39] | input_a[24]);
  assign popcount45_0xd7_core_090 = ~(input_a[2] & input_a[4]);
  assign popcount45_0xd7_core_093 = input_a[37] & input_a[40];
  assign popcount45_0xd7_core_094_not = ~input_a[22];
  assign popcount45_0xd7_core_095 = ~(input_a[38] | input_a[20]);
  assign popcount45_0xd7_core_099 = ~(input_a[14] | input_a[33]);
  assign popcount45_0xd7_core_100 = ~(input_a[15] & input_a[39]);
  assign popcount45_0xd7_core_101 = input_a[31] & input_a[19];
  assign popcount45_0xd7_core_104 = ~input_a[28];
  assign popcount45_0xd7_core_105 = ~(input_a[27] ^ input_a[35]);
  assign popcount45_0xd7_core_106 = input_a[5] & input_a[41];
  assign popcount45_0xd7_core_107 = ~(input_a[3] | input_a[4]);
  assign popcount45_0xd7_core_109 = ~(input_a[21] & input_a[43]);
  assign popcount45_0xd7_core_110 = ~(input_a[32] | input_a[24]);
  assign popcount45_0xd7_core_114 = input_a[20] & input_a[8];
  assign popcount45_0xd7_core_117 = ~(input_a[43] | input_a[24]);
  assign popcount45_0xd7_core_118 = popcount45_0xd7_core_106 & popcount45_0xd7_core_114;
  assign popcount45_0xd7_core_121 = input_a[0] | input_a[36];
  assign popcount45_0xd7_core_122 = ~input_a[4];
  assign popcount45_0xd7_core_123 = ~(input_a[14] ^ input_a[13]);
  assign popcount45_0xd7_core_124 = input_a[34] | input_a[19];
  assign popcount45_0xd7_core_125 = ~(input_a[32] & input_a[16]);
  assign popcount45_0xd7_core_126 = ~(input_a[12] & input_a[28]);
  assign popcount45_0xd7_core_127 = input_a[43] & input_a[34];
  assign popcount45_0xd7_core_128 = ~(input_a[42] ^ input_a[20]);
  assign popcount45_0xd7_core_130 = ~(input_a[10] & input_a[35]);
  assign popcount45_0xd7_core_131 = ~(input_a[14] | input_a[19]);
  assign popcount45_0xd7_core_132 = input_a[16] & input_a[42];
  assign popcount45_0xd7_core_133 = input_a[26] ^ input_a[21];
  assign popcount45_0xd7_core_134 = input_a[40] | input_a[13];
  assign popcount45_0xd7_core_136 = ~input_a[44];
  assign popcount45_0xd7_core_137 = ~input_a[11];
  assign popcount45_0xd7_core_139 = ~(input_a[22] & input_a[37]);
  assign popcount45_0xd7_core_140 = input_a[12] ^ input_a[10];
  assign popcount45_0xd7_core_141 = ~(input_a[1] ^ input_a[19]);
  assign popcount45_0xd7_core_142 = ~(input_a[38] | input_a[44]);
  assign popcount45_0xd7_core_143 = input_a[11] | input_a[26];
  assign popcount45_0xd7_core_145 = input_a[36] | input_a[34];
  assign popcount45_0xd7_core_147 = input_a[38] & input_a[41];
  assign popcount45_0xd7_core_149 = input_a[15] & popcount45_0xd7_core_136;
  assign popcount45_0xd7_core_150 = ~(input_a[10] ^ input_a[12]);
  assign popcount45_0xd7_core_151 = input_a[18] ^ input_a[21];
  assign popcount45_0xd7_core_153 = popcount45_0xd7_core_118 ^ popcount45_0xd7_core_143;
  assign popcount45_0xd7_core_154 = popcount45_0xd7_core_118 & popcount45_0xd7_core_143;
  assign popcount45_0xd7_core_155 = popcount45_0xd7_core_153 ^ popcount45_0xd7_core_149;
  assign popcount45_0xd7_core_156 = popcount45_0xd7_core_153 & popcount45_0xd7_core_149;
  assign popcount45_0xd7_core_157 = popcount45_0xd7_core_154 | popcount45_0xd7_core_156;
  assign popcount45_0xd7_core_159 = ~(input_a[35] & input_a[26]);
  assign popcount45_0xd7_core_167 = input_a[0] | input_a[7];
  assign popcount45_0xd7_core_168 = input_a[10] & input_a[1];
  assign popcount45_0xd7_core_170 = input_a[44] ^ popcount45_0xd7_core_155;
  assign popcount45_0xd7_core_171 = input_a[44] & popcount45_0xd7_core_155;
  assign popcount45_0xd7_core_172 = popcount45_0xd7_core_170 ^ popcount45_0xd7_core_168;
  assign popcount45_0xd7_core_173 = popcount45_0xd7_core_170 & popcount45_0xd7_core_168;
  assign popcount45_0xd7_core_174 = popcount45_0xd7_core_171 | popcount45_0xd7_core_173;
  assign popcount45_0xd7_core_177 = popcount45_0xd7_core_157 ^ popcount45_0xd7_core_174;
  assign popcount45_0xd7_core_178 = popcount45_0xd7_core_157 & popcount45_0xd7_core_174;
  assign popcount45_0xd7_core_181 = ~(input_a[44] | input_a[0]);
  assign popcount45_0xd7_core_185 = ~(input_a[12] ^ input_a[42]);
  assign popcount45_0xd7_core_191 = ~input_a[5];
  assign popcount45_0xd7_core_194 = ~(input_a[6] | input_a[0]);
  assign popcount45_0xd7_core_195 = ~(input_a[12] | input_a[35]);
  assign popcount45_0xd7_core_196 = input_a[12] ^ input_a[41];
  assign popcount45_0xd7_core_200 = input_a[39] & input_a[3];
  assign popcount45_0xd7_core_201 = ~(input_a[14] & input_a[1]);
  assign popcount45_0xd7_core_202 = ~(input_a[20] ^ input_a[9]);
  assign popcount45_0xd7_core_206 = ~input_a[37];
  assign popcount45_0xd7_core_207 = ~(input_a[26] | input_a[13]);
  assign popcount45_0xd7_core_208 = ~(input_a[37] | input_a[17]);
  assign popcount45_0xd7_core_209 = input_a[14] | input_a[44];
  assign popcount45_0xd7_core_210 = input_a[12] & input_a[7];
  assign popcount45_0xd7_core_211 = ~(input_a[34] & input_a[24]);
  assign popcount45_0xd7_core_213 = input_a[22] | input_a[41];
  assign popcount45_0xd7_core_216 = ~(input_a[10] & input_a[19]);
  assign popcount45_0xd7_core_220 = ~(input_a[7] & input_a[18]);
  assign popcount45_0xd7_core_221 = ~(input_a[23] & input_a[39]);
  assign popcount45_0xd7_core_224 = ~(input_a[35] & input_a[15]);
  assign popcount45_0xd7_core_228 = input_a[6] & input_a[5];
  assign popcount45_0xd7_core_229 = ~(input_a[8] & input_a[31]);
  assign popcount45_0xd7_core_231 = ~(input_a[30] | input_a[43]);
  assign popcount45_0xd7_core_234 = ~input_a[14];
  assign popcount45_0xd7_core_240 = ~(input_a[20] & input_a[12]);
  assign popcount45_0xd7_core_241 = ~(input_a[13] ^ input_a[25]);
  assign popcount45_0xd7_core_249 = ~input_a[23];
  assign popcount45_0xd7_core_250 = ~(input_a[10] ^ input_a[30]);
  assign popcount45_0xd7_core_252 = ~(input_a[34] | input_a[9]);
  assign popcount45_0xd7_core_253 = ~(input_a[43] | input_a[3]);
  assign popcount45_0xd7_core_254 = ~(input_a[21] & input_a[43]);
  assign popcount45_0xd7_core_255 = ~(input_a[32] & input_a[33]);
  assign popcount45_0xd7_core_257 = ~(input_a[34] | input_a[27]);
  assign popcount45_0xd7_core_258 = ~(input_a[20] & input_a[15]);
  assign popcount45_0xd7_core_259 = ~(input_a[35] | input_a[41]);
  assign popcount45_0xd7_core_260 = input_a[15] | input_a[42];
  assign popcount45_0xd7_core_263 = ~(input_a[27] & input_a[2]);
  assign popcount45_0xd7_core_265 = ~input_a[24];
  assign popcount45_0xd7_core_266 = input_a[2] & input_a[41];
  assign popcount45_0xd7_core_267_not = ~input_a[13];
  assign popcount45_0xd7_core_268 = input_a[24] | input_a[43];
  assign popcount45_0xd7_core_269 = ~input_a[43];
  assign popcount45_0xd7_core_271 = input_a[33] & input_a[6];
  assign popcount45_0xd7_core_275 = input_a[11] ^ input_a[21];
  assign popcount45_0xd7_core_277 = ~(input_a[20] | input_a[17]);
  assign popcount45_0xd7_core_278 = ~(input_a[35] | input_a[17]);
  assign popcount45_0xd7_core_281 = ~input_a[14];
  assign popcount45_0xd7_core_282 = input_a[27] ^ input_a[23];
  assign popcount45_0xd7_core_283 = ~input_a[2];
  assign popcount45_0xd7_core_284 = ~input_a[30];
  assign popcount45_0xd7_core_286 = ~input_a[21];
  assign popcount45_0xd7_core_287 = ~input_a[17];
  assign popcount45_0xd7_core_288_not = ~input_a[8];
  assign popcount45_0xd7_core_289 = ~(input_a[2] ^ input_a[23]);
  assign popcount45_0xd7_core_290 = ~(input_a[15] & input_a[25]);
  assign popcount45_0xd7_core_291 = ~input_a[15];
  assign popcount45_0xd7_core_292 = ~(input_a[2] & input_a[1]);
  assign popcount45_0xd7_core_293 = ~(input_a[35] ^ input_a[1]);
  assign popcount45_0xd7_core_294 = ~(input_a[40] ^ input_a[30]);
  assign popcount45_0xd7_core_295 = input_a[11] | input_a[13];
  assign popcount45_0xd7_core_298 = ~input_a[39];
  assign popcount45_0xd7_core_299 = ~(input_a[1] | input_a[30]);
  assign popcount45_0xd7_core_300 = ~input_a[35];
  assign popcount45_0xd7_core_301 = ~(input_a[0] ^ input_a[24]);
  assign popcount45_0xd7_core_302 = ~(input_a[11] | input_a[10]);
  assign popcount45_0xd7_core_303 = ~(input_a[32] & input_a[37]);
  assign popcount45_0xd7_core_305 = input_a[1] | input_a[20];
  assign popcount45_0xd7_core_306 = ~input_a[26];
  assign popcount45_0xd7_core_309 = input_a[35] ^ input_a[17];
  assign popcount45_0xd7_core_310 = input_a[27] ^ input_a[7];
  assign popcount45_0xd7_core_312 = input_a[33] & input_a[30];
  assign popcount45_0xd7_core_316 = ~input_a[29];
  assign popcount45_0xd7_core_318 = input_a[5] & input_a[2];
  assign popcount45_0xd7_core_319 = ~(input_a[28] & input_a[43]);
  assign popcount45_0xd7_core_320 = ~input_a[35];
  assign popcount45_0xd7_core_321 = input_a[31] & input_a[0];
  assign popcount45_0xd7_core_323 = ~input_a[40];
  assign popcount45_0xd7_core_324 = ~(input_a[23] & input_a[33]);
  assign popcount45_0xd7_core_326 = input_a[1] ^ input_a[6];
  assign popcount45_0xd7_core_327 = ~input_a[4];
  assign popcount45_0xd7_core_328 = input_a[33] & input_a[40];
  assign popcount45_0xd7_core_329 = input_a[41] | input_a[27];
  assign popcount45_0xd7_core_330 = ~(input_a[3] | input_a[37]);
  assign popcount45_0xd7_core_332 = input_a[38] ^ input_a[39];
  assign popcount45_0xd7_core_333 = input_a[13] | input_a[26];
  assign popcount45_0xd7_core_336 = input_a[4] & input_a[12];
  assign popcount45_0xd7_core_337 = popcount45_0xd7_core_172 ^ popcount45_0xd7_core_300;
  assign popcount45_0xd7_core_338 = popcount45_0xd7_core_172 & popcount45_0xd7_core_300;
  assign popcount45_0xd7_core_342 = popcount45_0xd7_core_177 ^ popcount45_0xd7_core_320;
  assign popcount45_0xd7_core_344 = popcount45_0xd7_core_342 ^ popcount45_0xd7_core_338;
  assign popcount45_0xd7_core_345 = popcount45_0xd7_core_342 & popcount45_0xd7_core_338;
  assign popcount45_0xd7_core_346 = popcount45_0xd7_core_177 | popcount45_0xd7_core_345;
  assign popcount45_0xd7_core_347 = popcount45_0xd7_core_178 ^ input_a[35];
  assign popcount45_0xd7_core_348 = popcount45_0xd7_core_178 & input_a[35];
  assign popcount45_0xd7_core_349 = popcount45_0xd7_core_347 | popcount45_0xd7_core_346;
  assign popcount45_0xd7_core_350 = input_a[27] | input_a[14];
  assign popcount45_0xd7_core_351 = ~input_a[26];
  assign popcount45_0xd7_core_352 = ~(input_a[37] & input_a[20]);
  assign popcount45_0xd7_core_353 = ~(input_a[5] & input_a[12]);
  assign popcount45_0xd7_core_354 = ~(input_a[42] | input_a[35]);
  assign popcount45_0xd7_core_355 = ~(input_a[8] ^ input_a[15]);
  assign popcount45_0xd7_core_356 = ~(input_a[13] | input_a[13]);

  assign popcount45_0xd7_out[0] = input_a[23];
  assign popcount45_0xd7_out[1] = popcount45_0xd7_core_300;
  assign popcount45_0xd7_out[2] = popcount45_0xd7_core_337;
  assign popcount45_0xd7_out[3] = popcount45_0xd7_core_344;
  assign popcount45_0xd7_out[4] = popcount45_0xd7_core_349;
  assign popcount45_0xd7_out[5] = popcount45_0xd7_core_348;
endmodule