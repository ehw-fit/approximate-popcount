// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=9.00067
// WCE=25.0
// EP=0.999216%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_d3ei(input [31:0] input_a, output [5:0] popcount32_d3ei_out);
  wire popcount32_d3ei_core_035;
  wire popcount32_d3ei_core_037;
  wire popcount32_d3ei_core_038;
  wire popcount32_d3ei_core_041;
  wire popcount32_d3ei_core_042;
  wire popcount32_d3ei_core_043;
  wire popcount32_d3ei_core_045;
  wire popcount32_d3ei_core_047;
  wire popcount32_d3ei_core_048;
  wire popcount32_d3ei_core_050;
  wire popcount32_d3ei_core_051;
  wire popcount32_d3ei_core_054;
  wire popcount32_d3ei_core_055;
  wire popcount32_d3ei_core_056;
  wire popcount32_d3ei_core_057;
  wire popcount32_d3ei_core_058;
  wire popcount32_d3ei_core_060;
  wire popcount32_d3ei_core_061;
  wire popcount32_d3ei_core_062;
  wire popcount32_d3ei_core_064;
  wire popcount32_d3ei_core_065;
  wire popcount32_d3ei_core_066;
  wire popcount32_d3ei_core_067;
  wire popcount32_d3ei_core_068;
  wire popcount32_d3ei_core_070;
  wire popcount32_d3ei_core_072;
  wire popcount32_d3ei_core_074;
  wire popcount32_d3ei_core_075;
  wire popcount32_d3ei_core_076;
  wire popcount32_d3ei_core_077;
  wire popcount32_d3ei_core_078;
  wire popcount32_d3ei_core_080;
  wire popcount32_d3ei_core_081;
  wire popcount32_d3ei_core_084;
  wire popcount32_d3ei_core_085;
  wire popcount32_d3ei_core_086;
  wire popcount32_d3ei_core_090;
  wire popcount32_d3ei_core_093;
  wire popcount32_d3ei_core_094_not;
  wire popcount32_d3ei_core_096;
  wire popcount32_d3ei_core_097;
  wire popcount32_d3ei_core_098;
  wire popcount32_d3ei_core_102;
  wire popcount32_d3ei_core_105;
  wire popcount32_d3ei_core_107;
  wire popcount32_d3ei_core_110;
  wire popcount32_d3ei_core_111_not;
  wire popcount32_d3ei_core_112;
  wire popcount32_d3ei_core_114;
  wire popcount32_d3ei_core_116;
  wire popcount32_d3ei_core_118;
  wire popcount32_d3ei_core_119;
  wire popcount32_d3ei_core_120;
  wire popcount32_d3ei_core_122;
  wire popcount32_d3ei_core_124;
  wire popcount32_d3ei_core_125;
  wire popcount32_d3ei_core_126;
  wire popcount32_d3ei_core_127;
  wire popcount32_d3ei_core_129_not;
  wire popcount32_d3ei_core_130;
  wire popcount32_d3ei_core_132;
  wire popcount32_d3ei_core_135;
  wire popcount32_d3ei_core_138;
  wire popcount32_d3ei_core_139;
  wire popcount32_d3ei_core_142;
  wire popcount32_d3ei_core_143;
  wire popcount32_d3ei_core_144;
  wire popcount32_d3ei_core_145;
  wire popcount32_d3ei_core_146;
  wire popcount32_d3ei_core_147;
  wire popcount32_d3ei_core_148;
  wire popcount32_d3ei_core_149;
  wire popcount32_d3ei_core_150;
  wire popcount32_d3ei_core_151;
  wire popcount32_d3ei_core_152;
  wire popcount32_d3ei_core_155;
  wire popcount32_d3ei_core_156;
  wire popcount32_d3ei_core_157;
  wire popcount32_d3ei_core_158;
  wire popcount32_d3ei_core_159;
  wire popcount32_d3ei_core_160;
  wire popcount32_d3ei_core_161;
  wire popcount32_d3ei_core_163;
  wire popcount32_d3ei_core_164;
  wire popcount32_d3ei_core_165;
  wire popcount32_d3ei_core_167;
  wire popcount32_d3ei_core_169;
  wire popcount32_d3ei_core_170;
  wire popcount32_d3ei_core_172;
  wire popcount32_d3ei_core_173;
  wire popcount32_d3ei_core_175;
  wire popcount32_d3ei_core_176;
  wire popcount32_d3ei_core_178;
  wire popcount32_d3ei_core_179;
  wire popcount32_d3ei_core_182;
  wire popcount32_d3ei_core_184;
  wire popcount32_d3ei_core_186;
  wire popcount32_d3ei_core_187;
  wire popcount32_d3ei_core_188;
  wire popcount32_d3ei_core_189;
  wire popcount32_d3ei_core_190;
  wire popcount32_d3ei_core_191;
  wire popcount32_d3ei_core_192;
  wire popcount32_d3ei_core_193;
  wire popcount32_d3ei_core_194;
  wire popcount32_d3ei_core_195;
  wire popcount32_d3ei_core_196;
  wire popcount32_d3ei_core_198;
  wire popcount32_d3ei_core_200;
  wire popcount32_d3ei_core_201;
  wire popcount32_d3ei_core_202;
  wire popcount32_d3ei_core_203_not;
  wire popcount32_d3ei_core_205;
  wire popcount32_d3ei_core_207;
  wire popcount32_d3ei_core_208;
  wire popcount32_d3ei_core_211;
  wire popcount32_d3ei_core_212;
  wire popcount32_d3ei_core_213;
  wire popcount32_d3ei_core_216;
  wire popcount32_d3ei_core_217;
  wire popcount32_d3ei_core_218;
  wire popcount32_d3ei_core_219;
  wire popcount32_d3ei_core_220;
  wire popcount32_d3ei_core_221;
  wire popcount32_d3ei_core_224;
  wire popcount32_d3ei_core_225;

  assign popcount32_d3ei_core_035 = input_a[13] | input_a[23];
  assign popcount32_d3ei_core_037 = ~input_a[12];
  assign popcount32_d3ei_core_038 = ~(input_a[14] ^ input_a[17]);
  assign popcount32_d3ei_core_041 = input_a[24] ^ input_a[0];
  assign popcount32_d3ei_core_042 = input_a[18] & input_a[2];
  assign popcount32_d3ei_core_043 = ~input_a[7];
  assign popcount32_d3ei_core_045 = input_a[2] | input_a[8];
  assign popcount32_d3ei_core_047 = input_a[24] & input_a[28];
  assign popcount32_d3ei_core_048 = ~input_a[29];
  assign popcount32_d3ei_core_050 = ~(input_a[23] ^ input_a[24]);
  assign popcount32_d3ei_core_051 = input_a[4] | input_a[13];
  assign popcount32_d3ei_core_054 = ~(input_a[21] ^ input_a[7]);
  assign popcount32_d3ei_core_055 = input_a[18] ^ input_a[27];
  assign popcount32_d3ei_core_056 = input_a[12] | input_a[17];
  assign popcount32_d3ei_core_057 = input_a[15] | input_a[9];
  assign popcount32_d3ei_core_058 = ~(input_a[6] ^ input_a[1]);
  assign popcount32_d3ei_core_060 = input_a[19] | input_a[18];
  assign popcount32_d3ei_core_061 = input_a[11] ^ input_a[0];
  assign popcount32_d3ei_core_062 = ~input_a[19];
  assign popcount32_d3ei_core_064 = input_a[1] ^ input_a[30];
  assign popcount32_d3ei_core_065 = input_a[18] & input_a[17];
  assign popcount32_d3ei_core_066 = input_a[19] & input_a[0];
  assign popcount32_d3ei_core_067 = input_a[15] | input_a[22];
  assign popcount32_d3ei_core_068 = ~(input_a[14] ^ input_a[10]);
  assign popcount32_d3ei_core_070 = ~input_a[10];
  assign popcount32_d3ei_core_072 = input_a[11] & input_a[21];
  assign popcount32_d3ei_core_074 = ~(input_a[24] & input_a[20]);
  assign popcount32_d3ei_core_075 = input_a[29] ^ input_a[1];
  assign popcount32_d3ei_core_076 = input_a[2] & input_a[18];
  assign popcount32_d3ei_core_077 = ~(input_a[29] ^ input_a[27]);
  assign popcount32_d3ei_core_078 = ~input_a[17];
  assign popcount32_d3ei_core_080 = input_a[12] | input_a[22];
  assign popcount32_d3ei_core_081 = ~(input_a[17] | input_a[18]);
  assign popcount32_d3ei_core_084 = ~(input_a[26] | input_a[8]);
  assign popcount32_d3ei_core_085 = ~(input_a[15] | input_a[6]);
  assign popcount32_d3ei_core_086 = input_a[26] | input_a[29];
  assign popcount32_d3ei_core_090 = input_a[8] ^ input_a[23];
  assign popcount32_d3ei_core_093 = input_a[13] & input_a[1];
  assign popcount32_d3ei_core_094_not = ~input_a[29];
  assign popcount32_d3ei_core_096 = input_a[3] ^ input_a[25];
  assign popcount32_d3ei_core_097 = ~(input_a[17] | input_a[20]);
  assign popcount32_d3ei_core_098 = input_a[29] & input_a[4];
  assign popcount32_d3ei_core_102 = ~(input_a[25] ^ input_a[2]);
  assign popcount32_d3ei_core_105 = ~(input_a[0] & input_a[19]);
  assign popcount32_d3ei_core_107 = input_a[19] & input_a[12];
  assign popcount32_d3ei_core_110 = ~(input_a[27] | input_a[15]);
  assign popcount32_d3ei_core_111_not = ~input_a[8];
  assign popcount32_d3ei_core_112 = ~(input_a[0] & input_a[7]);
  assign popcount32_d3ei_core_114 = input_a[23] | input_a[18];
  assign popcount32_d3ei_core_116 = ~(input_a[11] ^ input_a[9]);
  assign popcount32_d3ei_core_118 = input_a[13] ^ input_a[19];
  assign popcount32_d3ei_core_119 = input_a[0] ^ input_a[6];
  assign popcount32_d3ei_core_120 = ~(input_a[22] & input_a[18]);
  assign popcount32_d3ei_core_122 = ~(input_a[28] | input_a[12]);
  assign popcount32_d3ei_core_124 = ~(input_a[2] | input_a[28]);
  assign popcount32_d3ei_core_125 = ~input_a[5];
  assign popcount32_d3ei_core_126 = input_a[8] & input_a[24];
  assign popcount32_d3ei_core_127 = input_a[22] & input_a[14];
  assign popcount32_d3ei_core_129_not = ~input_a[14];
  assign popcount32_d3ei_core_130 = input_a[5] | input_a[16];
  assign popcount32_d3ei_core_132 = ~input_a[2];
  assign popcount32_d3ei_core_135 = ~(input_a[28] | input_a[2]);
  assign popcount32_d3ei_core_138 = input_a[6] | input_a[13];
  assign popcount32_d3ei_core_139 = ~(input_a[13] ^ input_a[6]);
  assign popcount32_d3ei_core_142 = input_a[29] | input_a[26];
  assign popcount32_d3ei_core_143 = input_a[26] ^ input_a[21];
  assign popcount32_d3ei_core_144 = ~(input_a[17] | input_a[31]);
  assign popcount32_d3ei_core_145 = ~(input_a[10] & input_a[19]);
  assign popcount32_d3ei_core_146 = input_a[8] & input_a[11];
  assign popcount32_d3ei_core_147 = input_a[25] & input_a[0];
  assign popcount32_d3ei_core_148 = ~(input_a[22] ^ input_a[1]);
  assign popcount32_d3ei_core_149 = input_a[18] ^ input_a[31];
  assign popcount32_d3ei_core_150 = input_a[18] | input_a[12];
  assign popcount32_d3ei_core_151 = ~(input_a[31] ^ input_a[12]);
  assign popcount32_d3ei_core_152 = input_a[1] | input_a[30];
  assign popcount32_d3ei_core_155 = ~(input_a[7] & input_a[3]);
  assign popcount32_d3ei_core_156 = ~(input_a[1] & input_a[8]);
  assign popcount32_d3ei_core_157 = ~(input_a[26] ^ input_a[29]);
  assign popcount32_d3ei_core_158 = input_a[12] & input_a[17];
  assign popcount32_d3ei_core_159 = ~(input_a[19] & input_a[10]);
  assign popcount32_d3ei_core_160 = input_a[19] ^ input_a[10];
  assign popcount32_d3ei_core_161 = input_a[31] & input_a[22];
  assign popcount32_d3ei_core_163 = input_a[18] ^ input_a[10];
  assign popcount32_d3ei_core_164 = ~(input_a[21] ^ input_a[19]);
  assign popcount32_d3ei_core_165 = input_a[30] & input_a[30];
  assign popcount32_d3ei_core_167 = ~(input_a[16] & input_a[12]);
  assign popcount32_d3ei_core_169 = input_a[2] | input_a[30];
  assign popcount32_d3ei_core_170 = input_a[15] ^ input_a[13];
  assign popcount32_d3ei_core_172 = ~(input_a[0] | input_a[31]);
  assign popcount32_d3ei_core_173 = ~(input_a[15] | input_a[29]);
  assign popcount32_d3ei_core_175 = ~(input_a[1] | input_a[13]);
  assign popcount32_d3ei_core_176 = ~input_a[28];
  assign popcount32_d3ei_core_178 = input_a[8] & input_a[15];
  assign popcount32_d3ei_core_179 = input_a[1] ^ input_a[26];
  assign popcount32_d3ei_core_182 = ~(input_a[15] & input_a[15]);
  assign popcount32_d3ei_core_184 = input_a[30] ^ input_a[24];
  assign popcount32_d3ei_core_186 = ~(input_a[13] ^ input_a[4]);
  assign popcount32_d3ei_core_187 = ~(input_a[17] & input_a[28]);
  assign popcount32_d3ei_core_188 = input_a[12] ^ input_a[13];
  assign popcount32_d3ei_core_189 = input_a[24] ^ input_a[27];
  assign popcount32_d3ei_core_190 = ~(input_a[17] ^ input_a[7]);
  assign popcount32_d3ei_core_191 = input_a[24] & input_a[5];
  assign popcount32_d3ei_core_192 = ~(input_a[16] & input_a[16]);
  assign popcount32_d3ei_core_193 = input_a[31] | input_a[3];
  assign popcount32_d3ei_core_194 = ~input_a[5];
  assign popcount32_d3ei_core_195 = input_a[30] & input_a[13];
  assign popcount32_d3ei_core_196 = input_a[15] & input_a[14];
  assign popcount32_d3ei_core_198 = ~(input_a[9] & input_a[1]);
  assign popcount32_d3ei_core_200 = input_a[16] & input_a[28];
  assign popcount32_d3ei_core_201 = input_a[26] & input_a[3];
  assign popcount32_d3ei_core_202 = ~(input_a[29] | input_a[10]);
  assign popcount32_d3ei_core_203_not = ~input_a[5];
  assign popcount32_d3ei_core_205 = input_a[2] ^ input_a[26];
  assign popcount32_d3ei_core_207 = ~(input_a[19] & input_a[11]);
  assign popcount32_d3ei_core_208 = ~(input_a[20] | input_a[11]);
  assign popcount32_d3ei_core_211 = input_a[24] ^ input_a[14];
  assign popcount32_d3ei_core_212 = ~input_a[0];
  assign popcount32_d3ei_core_213 = input_a[0] ^ input_a[25];
  assign popcount32_d3ei_core_216 = input_a[9] & input_a[25];
  assign popcount32_d3ei_core_217 = input_a[29] & input_a[12];
  assign popcount32_d3ei_core_218 = input_a[20] | input_a[21];
  assign popcount32_d3ei_core_219 = ~input_a[0];
  assign popcount32_d3ei_core_220 = input_a[20] ^ input_a[15];
  assign popcount32_d3ei_core_221 = input_a[1] ^ input_a[7];
  assign popcount32_d3ei_core_224 = ~(input_a[24] & input_a[5]);
  assign popcount32_d3ei_core_225 = ~(input_a[15] & input_a[15]);

  assign popcount32_d3ei_out[0] = 1'b1;
  assign popcount32_d3ei_out[1] = 1'b0;
  assign popcount32_d3ei_out[2] = 1'b0;
  assign popcount32_d3ei_out[3] = 1'b1;
  assign popcount32_d3ei_out[4] = 1'b1;
  assign popcount32_d3ei_out[5] = 1'b0;
endmodule