// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.78789
// WCE=15.0
// EP=0.890185%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_734b(input [24:0] input_a, output [4:0] popcount25_734b_out);
  wire popcount25_734b_core_027;
  wire popcount25_734b_core_028;
  wire popcount25_734b_core_029;
  wire popcount25_734b_core_030;
  wire popcount25_734b_core_032;
  wire popcount25_734b_core_033;
  wire popcount25_734b_core_035;
  wire popcount25_734b_core_036;
  wire popcount25_734b_core_037;
  wire popcount25_734b_core_038;
  wire popcount25_734b_core_041;
  wire popcount25_734b_core_043;
  wire popcount25_734b_core_044;
  wire popcount25_734b_core_045;
  wire popcount25_734b_core_051;
  wire popcount25_734b_core_052;
  wire popcount25_734b_core_054;
  wire popcount25_734b_core_055;
  wire popcount25_734b_core_057;
  wire popcount25_734b_core_058;
  wire popcount25_734b_core_059;
  wire popcount25_734b_core_061;
  wire popcount25_734b_core_062;
  wire popcount25_734b_core_064;
  wire popcount25_734b_core_065;
  wire popcount25_734b_core_066;
  wire popcount25_734b_core_069;
  wire popcount25_734b_core_070;
  wire popcount25_734b_core_073;
  wire popcount25_734b_core_075;
  wire popcount25_734b_core_076;
  wire popcount25_734b_core_077;
  wire popcount25_734b_core_078;
  wire popcount25_734b_core_080;
  wire popcount25_734b_core_081;
  wire popcount25_734b_core_083;
  wire popcount25_734b_core_085;
  wire popcount25_734b_core_086;
  wire popcount25_734b_core_090;
  wire popcount25_734b_core_091_not;
  wire popcount25_734b_core_092_not;
  wire popcount25_734b_core_094;
  wire popcount25_734b_core_099;
  wire popcount25_734b_core_100;
  wire popcount25_734b_core_101;
  wire popcount25_734b_core_102;
  wire popcount25_734b_core_103;
  wire popcount25_734b_core_104;
  wire popcount25_734b_core_105;
  wire popcount25_734b_core_107;
  wire popcount25_734b_core_108;
  wire popcount25_734b_core_109;
  wire popcount25_734b_core_110;
  wire popcount25_734b_core_112;
  wire popcount25_734b_core_115;
  wire popcount25_734b_core_116;
  wire popcount25_734b_core_118;
  wire popcount25_734b_core_120_not;
  wire popcount25_734b_core_123;
  wire popcount25_734b_core_125;
  wire popcount25_734b_core_126;
  wire popcount25_734b_core_127;
  wire popcount25_734b_core_128;
  wire popcount25_734b_core_129;
  wire popcount25_734b_core_130;
  wire popcount25_734b_core_131;
  wire popcount25_734b_core_133;
  wire popcount25_734b_core_135;
  wire popcount25_734b_core_137;
  wire popcount25_734b_core_139;
  wire popcount25_734b_core_141;
  wire popcount25_734b_core_142;
  wire popcount25_734b_core_143;
  wire popcount25_734b_core_144_not;
  wire popcount25_734b_core_148;
  wire popcount25_734b_core_149;
  wire popcount25_734b_core_150;
  wire popcount25_734b_core_152;
  wire popcount25_734b_core_153;
  wire popcount25_734b_core_156;
  wire popcount25_734b_core_157;
  wire popcount25_734b_core_158;
  wire popcount25_734b_core_160;
  wire popcount25_734b_core_162;
  wire popcount25_734b_core_165;
  wire popcount25_734b_core_166;
  wire popcount25_734b_core_167;
  wire popcount25_734b_core_168;
  wire popcount25_734b_core_169;
  wire popcount25_734b_core_170;
  wire popcount25_734b_core_171;
  wire popcount25_734b_core_172;
  wire popcount25_734b_core_173;
  wire popcount25_734b_core_174;
  wire popcount25_734b_core_175;
  wire popcount25_734b_core_176;
  wire popcount25_734b_core_178_not;
  wire popcount25_734b_core_179;
  wire popcount25_734b_core_182;
  wire popcount25_734b_core_183;

  assign popcount25_734b_core_027 = ~(input_a[20] & input_a[21]);
  assign popcount25_734b_core_028 = ~(input_a[7] ^ input_a[22]);
  assign popcount25_734b_core_029 = ~input_a[7];
  assign popcount25_734b_core_030 = ~(input_a[10] ^ input_a[2]);
  assign popcount25_734b_core_032 = ~(input_a[12] ^ input_a[16]);
  assign popcount25_734b_core_033 = input_a[11] & input_a[16];
  assign popcount25_734b_core_035 = ~input_a[21];
  assign popcount25_734b_core_036 = ~(input_a[24] & input_a[14]);
  assign popcount25_734b_core_037 = ~(input_a[15] & input_a[7]);
  assign popcount25_734b_core_038 = input_a[10] | input_a[2];
  assign popcount25_734b_core_041 = input_a[11] | input_a[11];
  assign popcount25_734b_core_043 = ~(input_a[14] ^ input_a[3]);
  assign popcount25_734b_core_044 = ~(input_a[4] ^ input_a[2]);
  assign popcount25_734b_core_045 = input_a[24] & input_a[14];
  assign popcount25_734b_core_051 = ~(input_a[8] | input_a[14]);
  assign popcount25_734b_core_052 = input_a[23] & input_a[7];
  assign popcount25_734b_core_054 = ~(input_a[15] & input_a[16]);
  assign popcount25_734b_core_055 = ~input_a[1];
  assign popcount25_734b_core_057 = input_a[1] & input_a[11];
  assign popcount25_734b_core_058 = input_a[15] | input_a[15];
  assign popcount25_734b_core_059 = input_a[13] | input_a[7];
  assign popcount25_734b_core_061 = input_a[7] | input_a[14];
  assign popcount25_734b_core_062 = input_a[8] | input_a[1];
  assign popcount25_734b_core_064 = input_a[11] ^ input_a[1];
  assign popcount25_734b_core_065 = ~input_a[1];
  assign popcount25_734b_core_066 = ~(input_a[11] | input_a[4]);
  assign popcount25_734b_core_069 = ~input_a[6];
  assign popcount25_734b_core_070 = input_a[15] | input_a[18];
  assign popcount25_734b_core_073 = ~input_a[18];
  assign popcount25_734b_core_075 = ~input_a[23];
  assign popcount25_734b_core_076 = ~(input_a[10] & input_a[18]);
  assign popcount25_734b_core_077 = ~(input_a[21] | input_a[19]);
  assign popcount25_734b_core_078 = ~(input_a[7] | input_a[11]);
  assign popcount25_734b_core_080 = input_a[16] & input_a[11];
  assign popcount25_734b_core_081 = ~(input_a[22] & input_a[10]);
  assign popcount25_734b_core_083 = ~input_a[22];
  assign popcount25_734b_core_085 = input_a[13] & input_a[8];
  assign popcount25_734b_core_086 = ~(input_a[21] | input_a[20]);
  assign popcount25_734b_core_090 = input_a[4] | input_a[12];
  assign popcount25_734b_core_091_not = ~input_a[7];
  assign popcount25_734b_core_092_not = ~input_a[1];
  assign popcount25_734b_core_094 = input_a[22] ^ input_a[0];
  assign popcount25_734b_core_099 = ~(input_a[13] ^ input_a[6]);
  assign popcount25_734b_core_100 = ~(input_a[3] & input_a[2]);
  assign popcount25_734b_core_101 = ~input_a[2];
  assign popcount25_734b_core_102 = ~(input_a[14] ^ input_a[5]);
  assign popcount25_734b_core_103 = input_a[3] & input_a[3];
  assign popcount25_734b_core_104 = ~(input_a[16] | input_a[23]);
  assign popcount25_734b_core_105 = input_a[0] & input_a[5];
  assign popcount25_734b_core_107 = input_a[18] | input_a[14];
  assign popcount25_734b_core_108 = input_a[23] | input_a[19];
  assign popcount25_734b_core_109 = ~(input_a[23] | input_a[10]);
  assign popcount25_734b_core_110 = ~input_a[2];
  assign popcount25_734b_core_112 = input_a[11] | input_a[1];
  assign popcount25_734b_core_115 = input_a[15] ^ input_a[0];
  assign popcount25_734b_core_116 = ~input_a[12];
  assign popcount25_734b_core_118 = input_a[20] ^ input_a[21];
  assign popcount25_734b_core_120_not = ~input_a[23];
  assign popcount25_734b_core_123 = ~(input_a[16] | input_a[24]);
  assign popcount25_734b_core_125 = ~(input_a[18] ^ input_a[8]);
  assign popcount25_734b_core_126 = ~(input_a[19] & input_a[3]);
  assign popcount25_734b_core_127 = input_a[16] & input_a[9];
  assign popcount25_734b_core_128 = input_a[22] ^ input_a[12];
  assign popcount25_734b_core_129 = ~(input_a[10] & input_a[1]);
  assign popcount25_734b_core_130 = ~(input_a[5] & input_a[5]);
  assign popcount25_734b_core_131 = input_a[24] & input_a[3];
  assign popcount25_734b_core_133 = ~(input_a[20] | input_a[15]);
  assign popcount25_734b_core_135 = ~input_a[6];
  assign popcount25_734b_core_137 = ~input_a[23];
  assign popcount25_734b_core_139 = ~(input_a[2] ^ input_a[21]);
  assign popcount25_734b_core_141 = input_a[3] & input_a[1];
  assign popcount25_734b_core_142 = input_a[3] & input_a[22];
  assign popcount25_734b_core_143 = input_a[14] & input_a[9];
  assign popcount25_734b_core_144_not = ~input_a[24];
  assign popcount25_734b_core_148 = ~(input_a[0] ^ input_a[12]);
  assign popcount25_734b_core_149 = ~input_a[22];
  assign popcount25_734b_core_150 = input_a[8] & input_a[2];
  assign popcount25_734b_core_152 = input_a[1] | input_a[16];
  assign popcount25_734b_core_153 = ~input_a[21];
  assign popcount25_734b_core_156 = ~(input_a[15] & input_a[23]);
  assign popcount25_734b_core_157 = input_a[22] | input_a[10];
  assign popcount25_734b_core_158 = ~input_a[22];
  assign popcount25_734b_core_160 = input_a[20] | input_a[14];
  assign popcount25_734b_core_162 = input_a[10] & input_a[4];
  assign popcount25_734b_core_165 = ~(input_a[4] | input_a[24]);
  assign popcount25_734b_core_166 = ~(input_a[24] & input_a[19]);
  assign popcount25_734b_core_167 = input_a[21] & input_a[16];
  assign popcount25_734b_core_168 = ~(input_a[10] & input_a[13]);
  assign popcount25_734b_core_169 = input_a[17] & input_a[18];
  assign popcount25_734b_core_170 = ~input_a[0];
  assign popcount25_734b_core_171 = input_a[23] | input_a[18];
  assign popcount25_734b_core_172 = ~(input_a[17] & input_a[6]);
  assign popcount25_734b_core_173 = input_a[10] & input_a[11];
  assign popcount25_734b_core_174 = ~(input_a[14] | input_a[11]);
  assign popcount25_734b_core_175 = ~(input_a[12] | input_a[0]);
  assign popcount25_734b_core_176 = ~(input_a[12] | input_a[13]);
  assign popcount25_734b_core_178_not = ~input_a[20];
  assign popcount25_734b_core_179 = input_a[12] | input_a[16];
  assign popcount25_734b_core_182 = ~(input_a[12] ^ input_a[7]);
  assign popcount25_734b_core_183 = ~(input_a[11] & input_a[6]);

  assign popcount25_734b_out[0] = input_a[20];
  assign popcount25_734b_out[1] = 1'b0;
  assign popcount25_734b_out[2] = input_a[0];
  assign popcount25_734b_out[3] = 1'b1;
  assign popcount25_734b_out[4] = 1'b0;
endmodule