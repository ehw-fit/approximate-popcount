// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.87753
// WCE=20.0
// EP=0.891571%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_yo1u(input [35:0] input_a, output [5:0] popcount36_yo1u_out);
  wire popcount36_yo1u_core_039;
  wire popcount36_yo1u_core_040;
  wire popcount36_yo1u_core_041_not;
  wire popcount36_yo1u_core_042;
  wire popcount36_yo1u_core_047;
  wire popcount36_yo1u_core_048;
  wire popcount36_yo1u_core_050;
  wire popcount36_yo1u_core_053;
  wire popcount36_yo1u_core_054;
  wire popcount36_yo1u_core_055;
  wire popcount36_yo1u_core_057;
  wire popcount36_yo1u_core_059;
  wire popcount36_yo1u_core_060;
  wire popcount36_yo1u_core_061;
  wire popcount36_yo1u_core_062;
  wire popcount36_yo1u_core_068;
  wire popcount36_yo1u_core_070;
  wire popcount36_yo1u_core_071;
  wire popcount36_yo1u_core_073;
  wire popcount36_yo1u_core_074;
  wire popcount36_yo1u_core_076;
  wire popcount36_yo1u_core_077;
  wire popcount36_yo1u_core_078;
  wire popcount36_yo1u_core_079;
  wire popcount36_yo1u_core_080;
  wire popcount36_yo1u_core_081;
  wire popcount36_yo1u_core_082;
  wire popcount36_yo1u_core_083;
  wire popcount36_yo1u_core_084;
  wire popcount36_yo1u_core_085;
  wire popcount36_yo1u_core_086;
  wire popcount36_yo1u_core_089;
  wire popcount36_yo1u_core_092;
  wire popcount36_yo1u_core_094;
  wire popcount36_yo1u_core_095_not;
  wire popcount36_yo1u_core_096;
  wire popcount36_yo1u_core_099;
  wire popcount36_yo1u_core_100;
  wire popcount36_yo1u_core_101;
  wire popcount36_yo1u_core_102;
  wire popcount36_yo1u_core_104;
  wire popcount36_yo1u_core_105;
  wire popcount36_yo1u_core_106;
  wire popcount36_yo1u_core_108;
  wire popcount36_yo1u_core_109;
  wire popcount36_yo1u_core_110;
  wire popcount36_yo1u_core_111;
  wire popcount36_yo1u_core_115;
  wire popcount36_yo1u_core_118;
  wire popcount36_yo1u_core_120;
  wire popcount36_yo1u_core_121;
  wire popcount36_yo1u_core_122;
  wire popcount36_yo1u_core_125;
  wire popcount36_yo1u_core_126;
  wire popcount36_yo1u_core_130;
  wire popcount36_yo1u_core_131;
  wire popcount36_yo1u_core_136;
  wire popcount36_yo1u_core_137;
  wire popcount36_yo1u_core_138;
  wire popcount36_yo1u_core_140;
  wire popcount36_yo1u_core_141_not;
  wire popcount36_yo1u_core_142_not;
  wire popcount36_yo1u_core_147;
  wire popcount36_yo1u_core_148;
  wire popcount36_yo1u_core_149;
  wire popcount36_yo1u_core_152;
  wire popcount36_yo1u_core_154;
  wire popcount36_yo1u_core_156;
  wire popcount36_yo1u_core_157;
  wire popcount36_yo1u_core_159;
  wire popcount36_yo1u_core_160;
  wire popcount36_yo1u_core_161;
  wire popcount36_yo1u_core_163;
  wire popcount36_yo1u_core_165;
  wire popcount36_yo1u_core_166;
  wire popcount36_yo1u_core_168;
  wire popcount36_yo1u_core_170;
  wire popcount36_yo1u_core_171;
  wire popcount36_yo1u_core_172;
  wire popcount36_yo1u_core_174;
  wire popcount36_yo1u_core_175;
  wire popcount36_yo1u_core_176;
  wire popcount36_yo1u_core_177;
  wire popcount36_yo1u_core_178;
  wire popcount36_yo1u_core_180;
  wire popcount36_yo1u_core_183;
  wire popcount36_yo1u_core_184;
  wire popcount36_yo1u_core_185;
  wire popcount36_yo1u_core_189;
  wire popcount36_yo1u_core_190;
  wire popcount36_yo1u_core_194;
  wire popcount36_yo1u_core_195;
  wire popcount36_yo1u_core_196;
  wire popcount36_yo1u_core_197;
  wire popcount36_yo1u_core_198;
  wire popcount36_yo1u_core_199;
  wire popcount36_yo1u_core_201;
  wire popcount36_yo1u_core_202;
  wire popcount36_yo1u_core_203;
  wire popcount36_yo1u_core_205;
  wire popcount36_yo1u_core_207;
  wire popcount36_yo1u_core_209;
  wire popcount36_yo1u_core_210;
  wire popcount36_yo1u_core_211;
  wire popcount36_yo1u_core_213;
  wire popcount36_yo1u_core_214;
  wire popcount36_yo1u_core_215;
  wire popcount36_yo1u_core_216;
  wire popcount36_yo1u_core_218;
  wire popcount36_yo1u_core_219_not;
  wire popcount36_yo1u_core_220;
  wire popcount36_yo1u_core_222;
  wire popcount36_yo1u_core_223;
  wire popcount36_yo1u_core_224;
  wire popcount36_yo1u_core_227;
  wire popcount36_yo1u_core_229;
  wire popcount36_yo1u_core_231;
  wire popcount36_yo1u_core_232;
  wire popcount36_yo1u_core_233;
  wire popcount36_yo1u_core_234;
  wire popcount36_yo1u_core_236;
  wire popcount36_yo1u_core_240;
  wire popcount36_yo1u_core_241;
  wire popcount36_yo1u_core_242;
  wire popcount36_yo1u_core_244;
  wire popcount36_yo1u_core_245;
  wire popcount36_yo1u_core_247;
  wire popcount36_yo1u_core_249;
  wire popcount36_yo1u_core_250;
  wire popcount36_yo1u_core_253;
  wire popcount36_yo1u_core_254;
  wire popcount36_yo1u_core_255;
  wire popcount36_yo1u_core_257;
  wire popcount36_yo1u_core_258;
  wire popcount36_yo1u_core_259;
  wire popcount36_yo1u_core_260;
  wire popcount36_yo1u_core_261;
  wire popcount36_yo1u_core_262;
  wire popcount36_yo1u_core_265;
  wire popcount36_yo1u_core_266;
  wire popcount36_yo1u_core_268;
  wire popcount36_yo1u_core_269;
  wire popcount36_yo1u_core_270;
  wire popcount36_yo1u_core_271;
  wire popcount36_yo1u_core_274;

  assign popcount36_yo1u_core_039 = input_a[16] ^ input_a[23];
  assign popcount36_yo1u_core_040 = input_a[27] ^ input_a[19];
  assign popcount36_yo1u_core_041_not = ~input_a[26];
  assign popcount36_yo1u_core_042 = ~input_a[26];
  assign popcount36_yo1u_core_047 = ~(input_a[13] | input_a[30]);
  assign popcount36_yo1u_core_048 = input_a[15] ^ input_a[16];
  assign popcount36_yo1u_core_050 = ~(input_a[6] & input_a[27]);
  assign popcount36_yo1u_core_053 = ~(input_a[24] | input_a[7]);
  assign popcount36_yo1u_core_054 = ~(input_a[11] | input_a[26]);
  assign popcount36_yo1u_core_055 = input_a[26] | input_a[9];
  assign popcount36_yo1u_core_057 = input_a[33] & input_a[12];
  assign popcount36_yo1u_core_059 = input_a[13] | input_a[30];
  assign popcount36_yo1u_core_060 = input_a[11] & input_a[2];
  assign popcount36_yo1u_core_061 = ~(input_a[15] | input_a[12]);
  assign popcount36_yo1u_core_062 = ~(input_a[26] & input_a[16]);
  assign popcount36_yo1u_core_068 = input_a[3] | input_a[33];
  assign popcount36_yo1u_core_070 = input_a[21] ^ input_a[18];
  assign popcount36_yo1u_core_071 = ~(input_a[13] | input_a[23]);
  assign popcount36_yo1u_core_073 = ~(input_a[24] & input_a[30]);
  assign popcount36_yo1u_core_074 = ~(input_a[5] & input_a[7]);
  assign popcount36_yo1u_core_076 = ~input_a[4];
  assign popcount36_yo1u_core_077 = ~(input_a[14] ^ input_a[3]);
  assign popcount36_yo1u_core_078 = ~(input_a[35] | input_a[3]);
  assign popcount36_yo1u_core_079 = ~(input_a[17] ^ input_a[2]);
  assign popcount36_yo1u_core_080 = input_a[14] | input_a[24];
  assign popcount36_yo1u_core_081 = input_a[35] & input_a[14];
  assign popcount36_yo1u_core_082 = input_a[8] & input_a[31];
  assign popcount36_yo1u_core_083 = input_a[27] & input_a[8];
  assign popcount36_yo1u_core_084 = ~(input_a[0] & input_a[16]);
  assign popcount36_yo1u_core_085 = ~(input_a[9] ^ input_a[15]);
  assign popcount36_yo1u_core_086 = ~(input_a[2] | input_a[25]);
  assign popcount36_yo1u_core_089 = ~(input_a[15] & input_a[34]);
  assign popcount36_yo1u_core_092 = input_a[7] & input_a[16];
  assign popcount36_yo1u_core_094 = input_a[26] ^ input_a[24];
  assign popcount36_yo1u_core_095_not = ~input_a[31];
  assign popcount36_yo1u_core_096 = ~(input_a[14] | input_a[28]);
  assign popcount36_yo1u_core_099 = ~input_a[6];
  assign popcount36_yo1u_core_100 = ~(input_a[21] & input_a[9]);
  assign popcount36_yo1u_core_101 = input_a[20] | input_a[26];
  assign popcount36_yo1u_core_102 = ~input_a[2];
  assign popcount36_yo1u_core_104 = input_a[16] ^ input_a[1];
  assign popcount36_yo1u_core_105 = input_a[22] & input_a[27];
  assign popcount36_yo1u_core_106 = ~(input_a[21] | input_a[7]);
  assign popcount36_yo1u_core_108 = input_a[29] | input_a[8];
  assign popcount36_yo1u_core_109 = input_a[19] & input_a[22];
  assign popcount36_yo1u_core_110 = input_a[16] ^ input_a[12];
  assign popcount36_yo1u_core_111 = ~(input_a[26] ^ input_a[2]);
  assign popcount36_yo1u_core_115 = ~input_a[0];
  assign popcount36_yo1u_core_118 = ~(input_a[0] ^ input_a[32]);
  assign popcount36_yo1u_core_120 = input_a[35] ^ input_a[19];
  assign popcount36_yo1u_core_121 = input_a[18] ^ input_a[12];
  assign popcount36_yo1u_core_122 = ~(input_a[3] | input_a[18]);
  assign popcount36_yo1u_core_125 = ~(input_a[6] & input_a[2]);
  assign popcount36_yo1u_core_126 = input_a[27] & input_a[14];
  assign popcount36_yo1u_core_130 = ~input_a[21];
  assign popcount36_yo1u_core_131 = ~(input_a[1] & input_a[18]);
  assign popcount36_yo1u_core_136 = ~(input_a[9] | input_a[11]);
  assign popcount36_yo1u_core_137 = ~(input_a[34] ^ input_a[12]);
  assign popcount36_yo1u_core_138 = input_a[14] & input_a[34];
  assign popcount36_yo1u_core_140 = input_a[2] ^ input_a[24];
  assign popcount36_yo1u_core_141_not = ~input_a[20];
  assign popcount36_yo1u_core_142_not = ~input_a[14];
  assign popcount36_yo1u_core_147 = ~(input_a[26] ^ input_a[25]);
  assign popcount36_yo1u_core_148 = input_a[11] & input_a[4];
  assign popcount36_yo1u_core_149 = ~(input_a[29] & input_a[27]);
  assign popcount36_yo1u_core_152 = ~input_a[4];
  assign popcount36_yo1u_core_154 = input_a[28] | input_a[7];
  assign popcount36_yo1u_core_156 = ~(input_a[4] | input_a[25]);
  assign popcount36_yo1u_core_157 = ~input_a[1];
  assign popcount36_yo1u_core_159 = ~input_a[30];
  assign popcount36_yo1u_core_160 = input_a[3] ^ input_a[11];
  assign popcount36_yo1u_core_161 = input_a[9] ^ input_a[35];
  assign popcount36_yo1u_core_163 = ~(input_a[28] & input_a[16]);
  assign popcount36_yo1u_core_165 = input_a[17] & input_a[34];
  assign popcount36_yo1u_core_166 = input_a[9] | input_a[33];
  assign popcount36_yo1u_core_168 = input_a[5] | input_a[27];
  assign popcount36_yo1u_core_170 = ~(input_a[21] & input_a[23]);
  assign popcount36_yo1u_core_171 = ~(input_a[12] | input_a[31]);
  assign popcount36_yo1u_core_172 = ~(input_a[13] ^ input_a[20]);
  assign popcount36_yo1u_core_174 = ~(input_a[31] ^ input_a[4]);
  assign popcount36_yo1u_core_175 = ~(input_a[10] ^ input_a[33]);
  assign popcount36_yo1u_core_176 = ~(input_a[32] | input_a[26]);
  assign popcount36_yo1u_core_177 = ~input_a[6];
  assign popcount36_yo1u_core_178 = ~(input_a[29] & input_a[24]);
  assign popcount36_yo1u_core_180 = ~(input_a[7] | input_a[4]);
  assign popcount36_yo1u_core_183 = ~input_a[24];
  assign popcount36_yo1u_core_184 = ~(input_a[12] & input_a[4]);
  assign popcount36_yo1u_core_185 = input_a[2] | input_a[34];
  assign popcount36_yo1u_core_189 = input_a[24] | input_a[0];
  assign popcount36_yo1u_core_190 = input_a[21] | input_a[5];
  assign popcount36_yo1u_core_194 = ~(input_a[2] ^ input_a[3]);
  assign popcount36_yo1u_core_195 = ~input_a[22];
  assign popcount36_yo1u_core_196 = ~(input_a[29] | input_a[19]);
  assign popcount36_yo1u_core_197 = ~input_a[25];
  assign popcount36_yo1u_core_198 = ~(input_a[22] ^ input_a[14]);
  assign popcount36_yo1u_core_199 = ~(input_a[5] & input_a[10]);
  assign popcount36_yo1u_core_201 = ~(input_a[8] | input_a[18]);
  assign popcount36_yo1u_core_202 = input_a[32] ^ input_a[1];
  assign popcount36_yo1u_core_203 = ~(input_a[6] ^ input_a[30]);
  assign popcount36_yo1u_core_205 = input_a[6] ^ input_a[21];
  assign popcount36_yo1u_core_207 = ~(input_a[4] ^ input_a[35]);
  assign popcount36_yo1u_core_209 = ~input_a[33];
  assign popcount36_yo1u_core_210 = input_a[20] | input_a[3];
  assign popcount36_yo1u_core_211 = ~(input_a[4] | input_a[10]);
  assign popcount36_yo1u_core_213 = ~(input_a[0] & input_a[27]);
  assign popcount36_yo1u_core_214 = input_a[29] | input_a[27];
  assign popcount36_yo1u_core_215 = input_a[33] | input_a[3];
  assign popcount36_yo1u_core_216 = ~(input_a[1] | input_a[25]);
  assign popcount36_yo1u_core_218 = input_a[1] ^ input_a[22];
  assign popcount36_yo1u_core_219_not = ~input_a[32];
  assign popcount36_yo1u_core_220 = ~(input_a[34] | input_a[26]);
  assign popcount36_yo1u_core_222 = ~(input_a[22] & input_a[32]);
  assign popcount36_yo1u_core_223 = ~(input_a[35] & input_a[27]);
  assign popcount36_yo1u_core_224 = ~(input_a[14] & input_a[3]);
  assign popcount36_yo1u_core_227 = ~(input_a[4] | input_a[10]);
  assign popcount36_yo1u_core_229 = input_a[21] | input_a[34];
  assign popcount36_yo1u_core_231 = input_a[5] | input_a[24];
  assign popcount36_yo1u_core_232 = ~(input_a[10] ^ input_a[3]);
  assign popcount36_yo1u_core_233 = input_a[21] | input_a[15];
  assign popcount36_yo1u_core_234 = ~(input_a[1] ^ input_a[3]);
  assign popcount36_yo1u_core_236 = ~(input_a[18] ^ input_a[18]);
  assign popcount36_yo1u_core_240 = input_a[17] ^ input_a[27];
  assign popcount36_yo1u_core_241 = input_a[14] ^ input_a[23];
  assign popcount36_yo1u_core_242 = ~input_a[18];
  assign popcount36_yo1u_core_244 = ~(input_a[24] ^ input_a[10]);
  assign popcount36_yo1u_core_245 = ~(input_a[27] & input_a[1]);
  assign popcount36_yo1u_core_247 = ~(input_a[17] & input_a[23]);
  assign popcount36_yo1u_core_249 = ~input_a[24];
  assign popcount36_yo1u_core_250 = input_a[34] | input_a[14];
  assign popcount36_yo1u_core_253 = input_a[7] ^ input_a[19];
  assign popcount36_yo1u_core_254 = ~(input_a[4] ^ input_a[6]);
  assign popcount36_yo1u_core_255 = input_a[17] & input_a[13];
  assign popcount36_yo1u_core_257 = ~input_a[6];
  assign popcount36_yo1u_core_258 = ~(input_a[29] | input_a[8]);
  assign popcount36_yo1u_core_259 = ~(input_a[21] & input_a[34]);
  assign popcount36_yo1u_core_260 = ~input_a[25];
  assign popcount36_yo1u_core_261 = input_a[13] & input_a[1];
  assign popcount36_yo1u_core_262 = input_a[29] & input_a[20];
  assign popcount36_yo1u_core_265 = ~input_a[29];
  assign popcount36_yo1u_core_266 = ~(input_a[13] ^ input_a[27]);
  assign popcount36_yo1u_core_268 = ~(input_a[4] & input_a[30]);
  assign popcount36_yo1u_core_269 = ~(input_a[15] ^ input_a[2]);
  assign popcount36_yo1u_core_270 = ~(input_a[8] & input_a[3]);
  assign popcount36_yo1u_core_271 = input_a[5] | input_a[5];
  assign popcount36_yo1u_core_274 = ~input_a[11];

  assign popcount36_yo1u_out[0] = input_a[0];
  assign popcount36_yo1u_out[1] = input_a[35];
  assign popcount36_yo1u_out[2] = input_a[33];
  assign popcount36_yo1u_out[3] = 1'b0;
  assign popcount36_yo1u_out[4] = 1'b1;
  assign popcount36_yo1u_out[5] = 1'b0;
endmodule