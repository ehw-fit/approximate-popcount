// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.41636
// WCE=28.0
// EP=0.953641%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_rrns(input [35:0] input_a, output [5:0] popcount36_rrns_out);
  wire popcount36_rrns_core_038;
  wire popcount36_rrns_core_039;
  wire popcount36_rrns_core_040;
  wire popcount36_rrns_core_041;
  wire popcount36_rrns_core_043;
  wire popcount36_rrns_core_044;
  wire popcount36_rrns_core_045;
  wire popcount36_rrns_core_046;
  wire popcount36_rrns_core_049;
  wire popcount36_rrns_core_050;
  wire popcount36_rrns_core_051;
  wire popcount36_rrns_core_052;
  wire popcount36_rrns_core_053;
  wire popcount36_rrns_core_054;
  wire popcount36_rrns_core_055;
  wire popcount36_rrns_core_056;
  wire popcount36_rrns_core_058;
  wire popcount36_rrns_core_059;
  wire popcount36_rrns_core_060;
  wire popcount36_rrns_core_061;
  wire popcount36_rrns_core_063;
  wire popcount36_rrns_core_065;
  wire popcount36_rrns_core_066;
  wire popcount36_rrns_core_067;
  wire popcount36_rrns_core_068;
  wire popcount36_rrns_core_070;
  wire popcount36_rrns_core_071;
  wire popcount36_rrns_core_074;
  wire popcount36_rrns_core_077_not;
  wire popcount36_rrns_core_079_not;
  wire popcount36_rrns_core_081;
  wire popcount36_rrns_core_082;
  wire popcount36_rrns_core_084;
  wire popcount36_rrns_core_086;
  wire popcount36_rrns_core_087;
  wire popcount36_rrns_core_088;
  wire popcount36_rrns_core_091;
  wire popcount36_rrns_core_092;
  wire popcount36_rrns_core_093;
  wire popcount36_rrns_core_095_not;
  wire popcount36_rrns_core_096;
  wire popcount36_rrns_core_098;
  wire popcount36_rrns_core_099;
  wire popcount36_rrns_core_101;
  wire popcount36_rrns_core_102_not;
  wire popcount36_rrns_core_104;
  wire popcount36_rrns_core_105;
  wire popcount36_rrns_core_106;
  wire popcount36_rrns_core_107;
  wire popcount36_rrns_core_108;
  wire popcount36_rrns_core_109;
  wire popcount36_rrns_core_113;
  wire popcount36_rrns_core_115;
  wire popcount36_rrns_core_116;
  wire popcount36_rrns_core_117;
  wire popcount36_rrns_core_118;
  wire popcount36_rrns_core_119;
  wire popcount36_rrns_core_121;
  wire popcount36_rrns_core_122;
  wire popcount36_rrns_core_123;
  wire popcount36_rrns_core_125;
  wire popcount36_rrns_core_126;
  wire popcount36_rrns_core_128;
  wire popcount36_rrns_core_129;
  wire popcount36_rrns_core_131;
  wire popcount36_rrns_core_135_not;
  wire popcount36_rrns_core_138;
  wire popcount36_rrns_core_140;
  wire popcount36_rrns_core_141;
  wire popcount36_rrns_core_143;
  wire popcount36_rrns_core_145;
  wire popcount36_rrns_core_147_not;
  wire popcount36_rrns_core_148;
  wire popcount36_rrns_core_151;
  wire popcount36_rrns_core_152;
  wire popcount36_rrns_core_154;
  wire popcount36_rrns_core_158;
  wire popcount36_rrns_core_159;
  wire popcount36_rrns_core_161;
  wire popcount36_rrns_core_162;
  wire popcount36_rrns_core_163;
  wire popcount36_rrns_core_164;
  wire popcount36_rrns_core_166;
  wire popcount36_rrns_core_168;
  wire popcount36_rrns_core_169;
  wire popcount36_rrns_core_170;
  wire popcount36_rrns_core_171;
  wire popcount36_rrns_core_172;
  wire popcount36_rrns_core_173;
  wire popcount36_rrns_core_174;
  wire popcount36_rrns_core_175;
  wire popcount36_rrns_core_176;
  wire popcount36_rrns_core_177;
  wire popcount36_rrns_core_180;
  wire popcount36_rrns_core_182;
  wire popcount36_rrns_core_183;
  wire popcount36_rrns_core_184;
  wire popcount36_rrns_core_185;
  wire popcount36_rrns_core_186;
  wire popcount36_rrns_core_187;
  wire popcount36_rrns_core_188;
  wire popcount36_rrns_core_190;
  wire popcount36_rrns_core_192;
  wire popcount36_rrns_core_194;
  wire popcount36_rrns_core_195;
  wire popcount36_rrns_core_197;
  wire popcount36_rrns_core_198;
  wire popcount36_rrns_core_199;
  wire popcount36_rrns_core_200;
  wire popcount36_rrns_core_201;
  wire popcount36_rrns_core_203;
  wire popcount36_rrns_core_205;
  wire popcount36_rrns_core_206;
  wire popcount36_rrns_core_207;
  wire popcount36_rrns_core_208;
  wire popcount36_rrns_core_209;
  wire popcount36_rrns_core_211;
  wire popcount36_rrns_core_215;
  wire popcount36_rrns_core_217;
  wire popcount36_rrns_core_218;
  wire popcount36_rrns_core_219;
  wire popcount36_rrns_core_220;
  wire popcount36_rrns_core_221;
  wire popcount36_rrns_core_222;
  wire popcount36_rrns_core_223;
  wire popcount36_rrns_core_224;
  wire popcount36_rrns_core_225;
  wire popcount36_rrns_core_226;
  wire popcount36_rrns_core_227;
  wire popcount36_rrns_core_228;
  wire popcount36_rrns_core_229;
  wire popcount36_rrns_core_230;
  wire popcount36_rrns_core_231;
  wire popcount36_rrns_core_232;
  wire popcount36_rrns_core_233;
  wire popcount36_rrns_core_234;
  wire popcount36_rrns_core_235;
  wire popcount36_rrns_core_236;
  wire popcount36_rrns_core_237;
  wire popcount36_rrns_core_240;
  wire popcount36_rrns_core_241;
  wire popcount36_rrns_core_243;
  wire popcount36_rrns_core_244;
  wire popcount36_rrns_core_245;
  wire popcount36_rrns_core_247;
  wire popcount36_rrns_core_250;
  wire popcount36_rrns_core_253;
  wire popcount36_rrns_core_255;
  wire popcount36_rrns_core_256;
  wire popcount36_rrns_core_257;
  wire popcount36_rrns_core_259;
  wire popcount36_rrns_core_260;
  wire popcount36_rrns_core_261;
  wire popcount36_rrns_core_262;
  wire popcount36_rrns_core_264;
  wire popcount36_rrns_core_265;
  wire popcount36_rrns_core_266;
  wire popcount36_rrns_core_267_not;
  wire popcount36_rrns_core_268;
  wire popcount36_rrns_core_269;
  wire popcount36_rrns_core_270;
  wire popcount36_rrns_core_272;
  wire popcount36_rrns_core_273;
  wire popcount36_rrns_core_274;
  wire popcount36_rrns_core_275;
  wire popcount36_rrns_core_276;

  assign popcount36_rrns_core_038 = input_a[27] | input_a[25];
  assign popcount36_rrns_core_039 = ~input_a[3];
  assign popcount36_rrns_core_040 = ~(input_a[0] ^ input_a[0]);
  assign popcount36_rrns_core_041 = ~(input_a[3] & input_a[4]);
  assign popcount36_rrns_core_043 = ~(input_a[4] ^ input_a[34]);
  assign popcount36_rrns_core_044 = input_a[31] ^ input_a[19];
  assign popcount36_rrns_core_045 = ~input_a[12];
  assign popcount36_rrns_core_046 = input_a[9] | input_a[3];
  assign popcount36_rrns_core_049 = input_a[24] & input_a[17];
  assign popcount36_rrns_core_050 = ~(input_a[16] ^ input_a[17]);
  assign popcount36_rrns_core_051 = input_a[0] & input_a[12];
  assign popcount36_rrns_core_052 = input_a[6] & input_a[11];
  assign popcount36_rrns_core_053 = input_a[35] & input_a[7];
  assign popcount36_rrns_core_054 = ~(input_a[32] & input_a[20]);
  assign popcount36_rrns_core_055 = input_a[11] ^ input_a[23];
  assign popcount36_rrns_core_056 = ~(input_a[22] & input_a[16]);
  assign popcount36_rrns_core_058 = input_a[1] ^ input_a[16];
  assign popcount36_rrns_core_059 = ~(input_a[12] | input_a[19]);
  assign popcount36_rrns_core_060 = ~(input_a[20] ^ input_a[14]);
  assign popcount36_rrns_core_061 = input_a[16] | input_a[20];
  assign popcount36_rrns_core_063 = input_a[18] & input_a[15];
  assign popcount36_rrns_core_065 = ~(input_a[33] ^ input_a[35]);
  assign popcount36_rrns_core_066 = ~(input_a[5] & input_a[1]);
  assign popcount36_rrns_core_067 = input_a[11] | input_a[34];
  assign popcount36_rrns_core_068 = input_a[33] ^ input_a[5];
  assign popcount36_rrns_core_070 = input_a[23] ^ input_a[11];
  assign popcount36_rrns_core_071 = ~input_a[27];
  assign popcount36_rrns_core_074 = ~(input_a[21] ^ input_a[7]);
  assign popcount36_rrns_core_077_not = ~input_a[13];
  assign popcount36_rrns_core_079_not = ~input_a[15];
  assign popcount36_rrns_core_081 = ~input_a[9];
  assign popcount36_rrns_core_082 = ~(input_a[9] ^ input_a[4]);
  assign popcount36_rrns_core_084 = ~(input_a[31] & input_a[1]);
  assign popcount36_rrns_core_086 = ~input_a[2];
  assign popcount36_rrns_core_087 = ~(input_a[9] & input_a[12]);
  assign popcount36_rrns_core_088 = input_a[0] ^ input_a[6];
  assign popcount36_rrns_core_091 = input_a[20] ^ input_a[23];
  assign popcount36_rrns_core_092 = ~(input_a[8] | input_a[32]);
  assign popcount36_rrns_core_093 = input_a[35] ^ input_a[16];
  assign popcount36_rrns_core_095_not = ~input_a[21];
  assign popcount36_rrns_core_096 = ~(input_a[27] & input_a[33]);
  assign popcount36_rrns_core_098 = input_a[21] ^ input_a[14];
  assign popcount36_rrns_core_099 = ~input_a[22];
  assign popcount36_rrns_core_101 = ~(input_a[31] ^ input_a[3]);
  assign popcount36_rrns_core_102_not = ~input_a[16];
  assign popcount36_rrns_core_104 = ~(input_a[35] ^ input_a[22]);
  assign popcount36_rrns_core_105 = ~(input_a[34] ^ input_a[6]);
  assign popcount36_rrns_core_106 = input_a[14] & input_a[25];
  assign popcount36_rrns_core_107 = ~(input_a[16] ^ input_a[18]);
  assign popcount36_rrns_core_108 = ~(input_a[11] ^ input_a[35]);
  assign popcount36_rrns_core_109 = ~(input_a[28] & input_a[30]);
  assign popcount36_rrns_core_113 = ~(input_a[24] ^ input_a[0]);
  assign popcount36_rrns_core_115 = ~input_a[15];
  assign popcount36_rrns_core_116 = input_a[28] ^ input_a[16];
  assign popcount36_rrns_core_117 = ~input_a[11];
  assign popcount36_rrns_core_118 = input_a[24] & input_a[28];
  assign popcount36_rrns_core_119 = ~input_a[6];
  assign popcount36_rrns_core_121 = input_a[4] & input_a[23];
  assign popcount36_rrns_core_122 = input_a[17] & input_a[12];
  assign popcount36_rrns_core_123 = input_a[12] | input_a[13];
  assign popcount36_rrns_core_125 = ~input_a[8];
  assign popcount36_rrns_core_126 = ~(input_a[21] | input_a[21]);
  assign popcount36_rrns_core_128 = input_a[21] ^ input_a[7];
  assign popcount36_rrns_core_129 = input_a[1] | input_a[12];
  assign popcount36_rrns_core_131 = ~(input_a[28] ^ input_a[15]);
  assign popcount36_rrns_core_135_not = ~input_a[29];
  assign popcount36_rrns_core_138 = ~(input_a[29] ^ input_a[4]);
  assign popcount36_rrns_core_140 = ~input_a[6];
  assign popcount36_rrns_core_141 = ~(input_a[24] ^ input_a[3]);
  assign popcount36_rrns_core_143 = input_a[21] & input_a[6];
  assign popcount36_rrns_core_145 = ~input_a[34];
  assign popcount36_rrns_core_147_not = ~input_a[30];
  assign popcount36_rrns_core_148 = input_a[7] & input_a[31];
  assign popcount36_rrns_core_151 = ~(input_a[16] | input_a[6]);
  assign popcount36_rrns_core_152 = input_a[2] | input_a[19];
  assign popcount36_rrns_core_154 = ~(input_a[14] & input_a[12]);
  assign popcount36_rrns_core_158 = ~(input_a[1] ^ input_a[35]);
  assign popcount36_rrns_core_159 = input_a[33] | input_a[19];
  assign popcount36_rrns_core_161 = ~(input_a[7] & input_a[9]);
  assign popcount36_rrns_core_162 = ~input_a[7];
  assign popcount36_rrns_core_163 = ~(input_a[4] ^ input_a[10]);
  assign popcount36_rrns_core_164 = ~(input_a[21] | input_a[25]);
  assign popcount36_rrns_core_166 = input_a[7] | input_a[29];
  assign popcount36_rrns_core_168 = ~(input_a[31] ^ input_a[11]);
  assign popcount36_rrns_core_169 = ~input_a[15];
  assign popcount36_rrns_core_170 = ~(input_a[3] ^ input_a[18]);
  assign popcount36_rrns_core_171 = ~(input_a[26] ^ input_a[14]);
  assign popcount36_rrns_core_172 = ~(input_a[32] & input_a[19]);
  assign popcount36_rrns_core_173 = input_a[19] & input_a[31];
  assign popcount36_rrns_core_174 = ~(input_a[16] & input_a[25]);
  assign popcount36_rrns_core_175 = ~input_a[33];
  assign popcount36_rrns_core_176 = ~(input_a[1] & input_a[18]);
  assign popcount36_rrns_core_177 = ~(input_a[18] & input_a[12]);
  assign popcount36_rrns_core_180 = ~(input_a[12] ^ input_a[5]);
  assign popcount36_rrns_core_182 = ~(input_a[10] & input_a[33]);
  assign popcount36_rrns_core_183 = ~input_a[27];
  assign popcount36_rrns_core_184 = input_a[20] | input_a[1];
  assign popcount36_rrns_core_185 = input_a[19] ^ input_a[0];
  assign popcount36_rrns_core_186 = ~input_a[6];
  assign popcount36_rrns_core_187 = input_a[18] | input_a[8];
  assign popcount36_rrns_core_188 = ~(input_a[7] ^ input_a[8]);
  assign popcount36_rrns_core_190 = input_a[31] | input_a[11];
  assign popcount36_rrns_core_192 = input_a[0] ^ input_a[24];
  assign popcount36_rrns_core_194 = ~input_a[34];
  assign popcount36_rrns_core_195 = ~(input_a[14] | input_a[25]);
  assign popcount36_rrns_core_197 = input_a[18] & input_a[1];
  assign popcount36_rrns_core_198 = input_a[12] ^ input_a[8];
  assign popcount36_rrns_core_199 = ~input_a[35];
  assign popcount36_rrns_core_200 = ~(input_a[17] ^ input_a[28]);
  assign popcount36_rrns_core_201 = ~(input_a[16] & input_a[20]);
  assign popcount36_rrns_core_203 = input_a[24] & input_a[2];
  assign popcount36_rrns_core_205 = input_a[24] ^ input_a[34];
  assign popcount36_rrns_core_206 = input_a[20] & input_a[23];
  assign popcount36_rrns_core_207 = input_a[27] | input_a[22];
  assign popcount36_rrns_core_208 = input_a[33] & input_a[27];
  assign popcount36_rrns_core_209 = input_a[23] ^ input_a[34];
  assign popcount36_rrns_core_211 = input_a[7] | input_a[1];
  assign popcount36_rrns_core_215 = ~(input_a[33] & input_a[11]);
  assign popcount36_rrns_core_217 = input_a[19] & input_a[23];
  assign popcount36_rrns_core_218 = input_a[15] | input_a[12];
  assign popcount36_rrns_core_219 = ~(input_a[8] | input_a[33]);
  assign popcount36_rrns_core_220 = input_a[13] ^ input_a[7];
  assign popcount36_rrns_core_221 = input_a[16] ^ input_a[11];
  assign popcount36_rrns_core_222 = input_a[11] | input_a[33];
  assign popcount36_rrns_core_223 = ~(input_a[32] | input_a[2]);
  assign popcount36_rrns_core_224 = input_a[18] ^ input_a[27];
  assign popcount36_rrns_core_225 = input_a[28] | input_a[17];
  assign popcount36_rrns_core_226 = ~input_a[22];
  assign popcount36_rrns_core_227 = input_a[27] | input_a[4];
  assign popcount36_rrns_core_228 = ~input_a[34];
  assign popcount36_rrns_core_229 = input_a[7] | input_a[13];
  assign popcount36_rrns_core_230 = input_a[19] | input_a[1];
  assign popcount36_rrns_core_231 = input_a[15] & input_a[15];
  assign popcount36_rrns_core_232 = input_a[17] ^ input_a[2];
  assign popcount36_rrns_core_233 = ~(input_a[19] ^ input_a[29]);
  assign popcount36_rrns_core_234 = ~input_a[33];
  assign popcount36_rrns_core_235 = ~(input_a[15] ^ input_a[12]);
  assign popcount36_rrns_core_236 = ~input_a[13];
  assign popcount36_rrns_core_237 = ~input_a[20];
  assign popcount36_rrns_core_240 = input_a[4] | input_a[34];
  assign popcount36_rrns_core_241 = ~input_a[20];
  assign popcount36_rrns_core_243 = ~(input_a[3] & input_a[25]);
  assign popcount36_rrns_core_244 = input_a[9] ^ input_a[35];
  assign popcount36_rrns_core_245 = ~(input_a[16] & input_a[32]);
  assign popcount36_rrns_core_247 = ~input_a[31];
  assign popcount36_rrns_core_250 = ~(input_a[20] ^ input_a[10]);
  assign popcount36_rrns_core_253 = input_a[17] & input_a[33];
  assign popcount36_rrns_core_255 = ~(input_a[28] ^ input_a[10]);
  assign popcount36_rrns_core_256 = ~input_a[6];
  assign popcount36_rrns_core_257 = ~(input_a[1] & input_a[31]);
  assign popcount36_rrns_core_259 = input_a[34] & input_a[5];
  assign popcount36_rrns_core_260 = ~(input_a[9] ^ input_a[11]);
  assign popcount36_rrns_core_261 = ~(input_a[23] ^ input_a[27]);
  assign popcount36_rrns_core_262 = input_a[22] ^ input_a[24];
  assign popcount36_rrns_core_264 = input_a[28] ^ input_a[33];
  assign popcount36_rrns_core_265 = input_a[26] & input_a[33];
  assign popcount36_rrns_core_266 = ~(input_a[10] ^ input_a[22]);
  assign popcount36_rrns_core_267_not = ~input_a[34];
  assign popcount36_rrns_core_268 = input_a[32] | input_a[12];
  assign popcount36_rrns_core_269 = ~(input_a[5] ^ input_a[9]);
  assign popcount36_rrns_core_270 = ~input_a[21];
  assign popcount36_rrns_core_272 = ~input_a[0];
  assign popcount36_rrns_core_273 = ~(input_a[21] ^ input_a[20]);
  assign popcount36_rrns_core_274 = ~(input_a[17] | input_a[12]);
  assign popcount36_rrns_core_275 = ~(input_a[0] | input_a[18]);
  assign popcount36_rrns_core_276 = input_a[20] ^ input_a[0];

  assign popcount36_rrns_out[0] = 1'b1;
  assign popcount36_rrns_out[1] = input_a[17];
  assign popcount36_rrns_out[2] = input_a[15];
  assign popcount36_rrns_out[3] = input_a[26];
  assign popcount36_rrns_out[4] = 1'b1;
  assign popcount36_rrns_out[5] = 1'b0;
endmodule