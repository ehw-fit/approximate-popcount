// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.02935
// WCE=26.0
// EP=0.9628%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_wbjs(input [22:0] input_a, output [4:0] popcount23_wbjs_out);
  wire popcount23_wbjs_core_026;
  wire popcount23_wbjs_core_027;
  wire popcount23_wbjs_core_030;
  wire popcount23_wbjs_core_031;
  wire popcount23_wbjs_core_034;
  wire popcount23_wbjs_core_035;
  wire popcount23_wbjs_core_036;
  wire popcount23_wbjs_core_037;
  wire popcount23_wbjs_core_038;
  wire popcount23_wbjs_core_040;
  wire popcount23_wbjs_core_042;
  wire popcount23_wbjs_core_043_not;
  wire popcount23_wbjs_core_044;
  wire popcount23_wbjs_core_045;
  wire popcount23_wbjs_core_046;
  wire popcount23_wbjs_core_049;
  wire popcount23_wbjs_core_050;
  wire popcount23_wbjs_core_052;
  wire popcount23_wbjs_core_053;
  wire popcount23_wbjs_core_055;
  wire popcount23_wbjs_core_056;
  wire popcount23_wbjs_core_058;
  wire popcount23_wbjs_core_060;
  wire popcount23_wbjs_core_061;
  wire popcount23_wbjs_core_062;
  wire popcount23_wbjs_core_063;
  wire popcount23_wbjs_core_064;
  wire popcount23_wbjs_core_065;
  wire popcount23_wbjs_core_066;
  wire popcount23_wbjs_core_069;
  wire popcount23_wbjs_core_070;
  wire popcount23_wbjs_core_074;
  wire popcount23_wbjs_core_075_not;
  wire popcount23_wbjs_core_076;
  wire popcount23_wbjs_core_077;
  wire popcount23_wbjs_core_079;
  wire popcount23_wbjs_core_081;
  wire popcount23_wbjs_core_082;
  wire popcount23_wbjs_core_083;
  wire popcount23_wbjs_core_084;
  wire popcount23_wbjs_core_085;
  wire popcount23_wbjs_core_086;
  wire popcount23_wbjs_core_088;
  wire popcount23_wbjs_core_089;
  wire popcount23_wbjs_core_091;
  wire popcount23_wbjs_core_092;
  wire popcount23_wbjs_core_093;
  wire popcount23_wbjs_core_095;
  wire popcount23_wbjs_core_098;
  wire popcount23_wbjs_core_100;
  wire popcount23_wbjs_core_101;
  wire popcount23_wbjs_core_103;
  wire popcount23_wbjs_core_104;
  wire popcount23_wbjs_core_105;
  wire popcount23_wbjs_core_107;
  wire popcount23_wbjs_core_113;
  wire popcount23_wbjs_core_114;
  wire popcount23_wbjs_core_115;
  wire popcount23_wbjs_core_116;
  wire popcount23_wbjs_core_117_not;
  wire popcount23_wbjs_core_118;
  wire popcount23_wbjs_core_119;
  wire popcount23_wbjs_core_122;
  wire popcount23_wbjs_core_123;
  wire popcount23_wbjs_core_128;
  wire popcount23_wbjs_core_131;
  wire popcount23_wbjs_core_132;
  wire popcount23_wbjs_core_133;
  wire popcount23_wbjs_core_134;
  wire popcount23_wbjs_core_135;
  wire popcount23_wbjs_core_137_not;
  wire popcount23_wbjs_core_138;
  wire popcount23_wbjs_core_140_not;
  wire popcount23_wbjs_core_142;
  wire popcount23_wbjs_core_143;
  wire popcount23_wbjs_core_145;
  wire popcount23_wbjs_core_146;
  wire popcount23_wbjs_core_147;
  wire popcount23_wbjs_core_148;
  wire popcount23_wbjs_core_152;
  wire popcount23_wbjs_core_153;
  wire popcount23_wbjs_core_155;
  wire popcount23_wbjs_core_157;
  wire popcount23_wbjs_core_159;
  wire popcount23_wbjs_core_160;
  wire popcount23_wbjs_core_161;
  wire popcount23_wbjs_core_164;
  wire popcount23_wbjs_core_166;
  wire popcount23_wbjs_core_167;
  wire popcount23_wbjs_core_168_not;

  assign popcount23_wbjs_core_026 = ~(input_a[19] | input_a[12]);
  assign popcount23_wbjs_core_027 = input_a[8] & input_a[1];
  assign popcount23_wbjs_core_030 = input_a[20] & input_a[14];
  assign popcount23_wbjs_core_031 = ~(input_a[3] ^ input_a[21]);
  assign popcount23_wbjs_core_034 = ~(input_a[11] & input_a[15]);
  assign popcount23_wbjs_core_035 = ~input_a[0];
  assign popcount23_wbjs_core_036 = input_a[7] ^ input_a[21];
  assign popcount23_wbjs_core_037 = input_a[20] | input_a[18];
  assign popcount23_wbjs_core_038 = ~input_a[9];
  assign popcount23_wbjs_core_040 = ~(input_a[19] ^ input_a[2]);
  assign popcount23_wbjs_core_042 = input_a[6] | input_a[11];
  assign popcount23_wbjs_core_043_not = ~input_a[7];
  assign popcount23_wbjs_core_044 = input_a[21] & input_a[2];
  assign popcount23_wbjs_core_045 = ~(input_a[1] & input_a[6]);
  assign popcount23_wbjs_core_046 = ~(input_a[13] ^ input_a[17]);
  assign popcount23_wbjs_core_049 = ~(input_a[20] & input_a[6]);
  assign popcount23_wbjs_core_050 = input_a[11] | input_a[20];
  assign popcount23_wbjs_core_052 = ~(input_a[21] ^ input_a[11]);
  assign popcount23_wbjs_core_053 = ~(input_a[7] ^ input_a[8]);
  assign popcount23_wbjs_core_055 = ~input_a[4];
  assign popcount23_wbjs_core_056 = ~(input_a[19] | input_a[20]);
  assign popcount23_wbjs_core_058 = ~(input_a[20] ^ input_a[21]);
  assign popcount23_wbjs_core_060 = input_a[2] & input_a[22];
  assign popcount23_wbjs_core_061 = input_a[21] | input_a[3];
  assign popcount23_wbjs_core_062 = input_a[7] & input_a[3];
  assign popcount23_wbjs_core_063 = ~(input_a[18] ^ input_a[9]);
  assign popcount23_wbjs_core_064 = ~input_a[15];
  assign popcount23_wbjs_core_065 = ~(input_a[5] ^ input_a[19]);
  assign popcount23_wbjs_core_066 = ~input_a[16];
  assign popcount23_wbjs_core_069 = ~input_a[20];
  assign popcount23_wbjs_core_070 = ~(input_a[17] & input_a[4]);
  assign popcount23_wbjs_core_074 = ~input_a[14];
  assign popcount23_wbjs_core_075_not = ~input_a[3];
  assign popcount23_wbjs_core_076 = input_a[10] | input_a[22];
  assign popcount23_wbjs_core_077 = ~(input_a[18] | input_a[22]);
  assign popcount23_wbjs_core_079 = input_a[19] ^ input_a[16];
  assign popcount23_wbjs_core_081 = input_a[6] ^ input_a[1];
  assign popcount23_wbjs_core_082 = ~input_a[7];
  assign popcount23_wbjs_core_083 = input_a[8] | input_a[22];
  assign popcount23_wbjs_core_084 = ~(input_a[8] & input_a[5]);
  assign popcount23_wbjs_core_085 = input_a[6] | input_a[10];
  assign popcount23_wbjs_core_086 = ~(input_a[4] ^ input_a[17]);
  assign popcount23_wbjs_core_088 = ~(input_a[10] | input_a[7]);
  assign popcount23_wbjs_core_089 = input_a[12] & input_a[10];
  assign popcount23_wbjs_core_091 = ~(input_a[11] & input_a[0]);
  assign popcount23_wbjs_core_092 = ~(input_a[19] | input_a[3]);
  assign popcount23_wbjs_core_093 = ~(input_a[6] & input_a[9]);
  assign popcount23_wbjs_core_095 = ~(input_a[2] ^ input_a[0]);
  assign popcount23_wbjs_core_098 = ~input_a[1];
  assign popcount23_wbjs_core_100 = ~input_a[18];
  assign popcount23_wbjs_core_101 = input_a[22] | input_a[5];
  assign popcount23_wbjs_core_103 = ~input_a[22];
  assign popcount23_wbjs_core_104 = ~(input_a[8] ^ input_a[12]);
  assign popcount23_wbjs_core_105 = ~input_a[14];
  assign popcount23_wbjs_core_107 = input_a[16] ^ input_a[15];
  assign popcount23_wbjs_core_113 = ~(input_a[5] & input_a[6]);
  assign popcount23_wbjs_core_114 = input_a[14] | input_a[12];
  assign popcount23_wbjs_core_115 = ~(input_a[13] & input_a[10]);
  assign popcount23_wbjs_core_116 = input_a[19] & input_a[13];
  assign popcount23_wbjs_core_117_not = ~input_a[9];
  assign popcount23_wbjs_core_118 = input_a[21] ^ input_a[20];
  assign popcount23_wbjs_core_119 = ~(input_a[13] | input_a[21]);
  assign popcount23_wbjs_core_122 = input_a[14] ^ input_a[8];
  assign popcount23_wbjs_core_123 = ~input_a[8];
  assign popcount23_wbjs_core_128 = ~(input_a[3] ^ input_a[6]);
  assign popcount23_wbjs_core_131 = ~input_a[4];
  assign popcount23_wbjs_core_132 = ~input_a[21];
  assign popcount23_wbjs_core_133 = input_a[19] & input_a[10];
  assign popcount23_wbjs_core_134 = input_a[19] & input_a[1];
  assign popcount23_wbjs_core_135 = ~input_a[11];
  assign popcount23_wbjs_core_137_not = ~input_a[5];
  assign popcount23_wbjs_core_138 = input_a[11] | input_a[17];
  assign popcount23_wbjs_core_140_not = ~input_a[9];
  assign popcount23_wbjs_core_142 = input_a[0] & input_a[5];
  assign popcount23_wbjs_core_143 = ~(input_a[7] & input_a[14]);
  assign popcount23_wbjs_core_145 = ~(input_a[8] & input_a[7]);
  assign popcount23_wbjs_core_146 = input_a[22] | input_a[14];
  assign popcount23_wbjs_core_147 = ~(input_a[6] & input_a[8]);
  assign popcount23_wbjs_core_148 = ~(input_a[10] | input_a[19]);
  assign popcount23_wbjs_core_152 = ~input_a[19];
  assign popcount23_wbjs_core_153 = input_a[3] ^ input_a[11];
  assign popcount23_wbjs_core_155 = ~(input_a[4] | input_a[2]);
  assign popcount23_wbjs_core_157 = input_a[11] & input_a[4];
  assign popcount23_wbjs_core_159 = ~(input_a[7] ^ input_a[22]);
  assign popcount23_wbjs_core_160 = input_a[1] | input_a[22];
  assign popcount23_wbjs_core_161 = ~(input_a[0] & input_a[5]);
  assign popcount23_wbjs_core_164 = ~(input_a[13] | input_a[8]);
  assign popcount23_wbjs_core_166 = input_a[21] | input_a[2];
  assign popcount23_wbjs_core_167 = ~(input_a[9] & input_a[1]);
  assign popcount23_wbjs_core_168_not = ~input_a[12];

  assign popcount23_wbjs_out[0] = input_a[16];
  assign popcount23_wbjs_out[1] = input_a[0];
  assign popcount23_wbjs_out[2] = input_a[1];
  assign popcount23_wbjs_out[3] = input_a[5];
  assign popcount23_wbjs_out[4] = input_a[11];
endmodule