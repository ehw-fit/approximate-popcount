// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.66785
// WCE=9.0
// EP=0.905449%
// Printed PDK parameters:
//  Area=4731470.0
//  Delay=12188812.0
//  Power=259860.0

module popcount18_f88b(input [17:0] input_a, output [4:0] popcount18_f88b_out);
  wire popcount18_f88b_core_020;
  wire popcount18_f88b_core_021;
  wire popcount18_f88b_core_022;
  wire popcount18_f88b_core_023;
  wire popcount18_f88b_core_024;
  wire popcount18_f88b_core_025;
  wire popcount18_f88b_core_026;
  wire popcount18_f88b_core_027;
  wire popcount18_f88b_core_029;
  wire popcount18_f88b_core_031;
  wire popcount18_f88b_core_032;
  wire popcount18_f88b_core_033;
  wire popcount18_f88b_core_034;
  wire popcount18_f88b_core_035;
  wire popcount18_f88b_core_036;
  wire popcount18_f88b_core_037;
  wire popcount18_f88b_core_039;
  wire popcount18_f88b_core_040;
  wire popcount18_f88b_core_041;
  wire popcount18_f88b_core_042;
  wire popcount18_f88b_core_043;
  wire popcount18_f88b_core_044;
  wire popcount18_f88b_core_045;
  wire popcount18_f88b_core_047;
  wire popcount18_f88b_core_048;
  wire popcount18_f88b_core_049;
  wire popcount18_f88b_core_051;
  wire popcount18_f88b_core_052;
  wire popcount18_f88b_core_053;
  wire popcount18_f88b_core_054;
  wire popcount18_f88b_core_055;
  wire popcount18_f88b_core_056;
  wire popcount18_f88b_core_057;
  wire popcount18_f88b_core_058;
  wire popcount18_f88b_core_059;
  wire popcount18_f88b_core_060;
  wire popcount18_f88b_core_064;
  wire popcount18_f88b_core_065;
  wire popcount18_f88b_core_066;
  wire popcount18_f88b_core_067;
  wire popcount18_f88b_core_069;
  wire popcount18_f88b_core_070;
  wire popcount18_f88b_core_072;
  wire popcount18_f88b_core_073;
  wire popcount18_f88b_core_074;
  wire popcount18_f88b_core_075;
  wire popcount18_f88b_core_076;
  wire popcount18_f88b_core_077;
  wire popcount18_f88b_core_078;
  wire popcount18_f88b_core_081;
  wire popcount18_f88b_core_083;
  wire popcount18_f88b_core_084;
  wire popcount18_f88b_core_085;
  wire popcount18_f88b_core_086;
  wire popcount18_f88b_core_087;
  wire popcount18_f88b_core_088;
  wire popcount18_f88b_core_091;
  wire popcount18_f88b_core_093;
  wire popcount18_f88b_core_094;
  wire popcount18_f88b_core_095;
  wire popcount18_f88b_core_096;
  wire popcount18_f88b_core_097;
  wire popcount18_f88b_core_099;
  wire popcount18_f88b_core_100;
  wire popcount18_f88b_core_101;
  wire popcount18_f88b_core_102;
  wire popcount18_f88b_core_103;
  wire popcount18_f88b_core_104;
  wire popcount18_f88b_core_109;
  wire popcount18_f88b_core_110;
  wire popcount18_f88b_core_111;
  wire popcount18_f88b_core_112;
  wire popcount18_f88b_core_113;
  wire popcount18_f88b_core_114;
  wire popcount18_f88b_core_115;
  wire popcount18_f88b_core_116;
  wire popcount18_f88b_core_117;
  wire popcount18_f88b_core_118;
  wire popcount18_f88b_core_120;
  wire popcount18_f88b_core_123_not;
  wire popcount18_f88b_core_124;
  wire popcount18_f88b_core_125;

  assign popcount18_f88b_core_020 = ~(input_a[10] & input_a[17]);
  assign popcount18_f88b_core_021 = input_a[0] & input_a[15];
  assign popcount18_f88b_core_022 = ~(input_a[17] ^ input_a[13]);
  assign popcount18_f88b_core_023 = input_a[1] & input_a[2];
  assign popcount18_f88b_core_024 = ~popcount18_f88b_core_020;
  assign popcount18_f88b_core_025 = ~(input_a[16] & input_a[14]);
  assign popcount18_f88b_core_026 = ~(popcount18_f88b_core_021 & popcount18_f88b_core_023);
  assign popcount18_f88b_core_027 = popcount18_f88b_core_021 & popcount18_f88b_core_023;
  assign popcount18_f88b_core_029 = input_a[1] ^ input_a[17];
  assign popcount18_f88b_core_031 = ~(input_a[4] & input_a[5]);
  assign popcount18_f88b_core_032 = input_a[4] & input_a[5];
  assign popcount18_f88b_core_033 = ~(input_a[7] & input_a[8]);
  assign popcount18_f88b_core_034 = input_a[7] & input_a[8];
  assign popcount18_f88b_core_035 = input_a[6] ^ popcount18_f88b_core_033;
  assign popcount18_f88b_core_036 = input_a[12] & input_a[17];
  assign popcount18_f88b_core_037 = popcount18_f88b_core_034 | input_a[6];
  assign popcount18_f88b_core_039 = popcount18_f88b_core_031 ^ popcount18_f88b_core_035;
  assign popcount18_f88b_core_040 = popcount18_f88b_core_031 & popcount18_f88b_core_035;
  assign popcount18_f88b_core_041 = popcount18_f88b_core_032 ^ popcount18_f88b_core_037;
  assign popcount18_f88b_core_042 = popcount18_f88b_core_032 & popcount18_f88b_core_037;
  assign popcount18_f88b_core_043 = popcount18_f88b_core_041 ^ popcount18_f88b_core_040;
  assign popcount18_f88b_core_044 = input_a[6] & popcount18_f88b_core_040;
  assign popcount18_f88b_core_045 = popcount18_f88b_core_042 | popcount18_f88b_core_044;
  assign popcount18_f88b_core_047 = ~(input_a[6] | input_a[12]);
  assign popcount18_f88b_core_048 = ~input_a[0];
  assign popcount18_f88b_core_049 = popcount18_f88b_core_024 & popcount18_f88b_core_039;
  assign popcount18_f88b_core_051 = popcount18_f88b_core_026 & popcount18_f88b_core_043;
  assign popcount18_f88b_core_052 = ~(input_a[12] ^ input_a[8]);
  assign popcount18_f88b_core_053 = popcount18_f88b_core_026 & popcount18_f88b_core_049;
  assign popcount18_f88b_core_054 = popcount18_f88b_core_051 | popcount18_f88b_core_053;
  assign popcount18_f88b_core_055 = popcount18_f88b_core_027 ^ popcount18_f88b_core_045;
  assign popcount18_f88b_core_056 = popcount18_f88b_core_027 & popcount18_f88b_core_045;
  assign popcount18_f88b_core_057 = popcount18_f88b_core_055 ^ popcount18_f88b_core_054;
  assign popcount18_f88b_core_058 = popcount18_f88b_core_055 & popcount18_f88b_core_054;
  assign popcount18_f88b_core_059 = popcount18_f88b_core_056 | popcount18_f88b_core_058;
  assign popcount18_f88b_core_060 = ~(input_a[4] & input_a[5]);
  assign popcount18_f88b_core_064 = ~(input_a[13] & input_a[11]);
  assign popcount18_f88b_core_065 = input_a[0] & input_a[17];
  assign popcount18_f88b_core_066 = input_a[7] & input_a[15];
  assign popcount18_f88b_core_067 = input_a[1] | input_a[6];
  assign popcount18_f88b_core_069 = ~(input_a[8] | input_a[10]);
  assign popcount18_f88b_core_070 = ~input_a[0];
  assign popcount18_f88b_core_072 = input_a[10] ^ input_a[15];
  assign popcount18_f88b_core_073 = ~input_a[16];
  assign popcount18_f88b_core_074 = ~(input_a[6] ^ input_a[17]);
  assign popcount18_f88b_core_075 = ~(input_a[12] ^ input_a[4]);
  assign popcount18_f88b_core_076 = input_a[9] ^ input_a[5];
  assign popcount18_f88b_core_077 = ~(input_a[10] ^ input_a[14]);
  assign popcount18_f88b_core_078 = input_a[1] | input_a[10];
  assign popcount18_f88b_core_081 = ~input_a[0];
  assign popcount18_f88b_core_083 = input_a[16] & input_a[3];
  assign popcount18_f88b_core_084 = input_a[6] | input_a[15];
  assign popcount18_f88b_core_085 = input_a[11] & input_a[12];
  assign popcount18_f88b_core_086 = input_a[1] & input_a[10];
  assign popcount18_f88b_core_087 = ~(input_a[13] ^ input_a[3]);
  assign popcount18_f88b_core_088 = ~input_a[16];
  assign popcount18_f88b_core_091 = ~(input_a[13] ^ input_a[4]);
  assign popcount18_f88b_core_093 = ~(input_a[2] & input_a[11]);
  assign popcount18_f88b_core_094 = ~(input_a[2] & input_a[16]);
  assign popcount18_f88b_core_095 = ~input_a[0];
  assign popcount18_f88b_core_096 = ~input_a[12];
  assign popcount18_f88b_core_097 = ~input_a[6];
  assign popcount18_f88b_core_099 = ~input_a[6];
  assign popcount18_f88b_core_100 = input_a[4] | input_a[9];
  assign popcount18_f88b_core_101 = ~(input_a[12] | input_a[11]);
  assign popcount18_f88b_core_102 = ~(input_a[14] & input_a[0]);
  assign popcount18_f88b_core_103 = ~(input_a[10] ^ input_a[4]);
  assign popcount18_f88b_core_104 = input_a[7] & input_a[10];
  assign popcount18_f88b_core_109 = input_a[16] | input_a[10];
  assign popcount18_f88b_core_110 = input_a[17] | input_a[6];
  assign popcount18_f88b_core_111 = ~(input_a[9] | input_a[9]);
  assign popcount18_f88b_core_112 = ~input_a[2];
  assign popcount18_f88b_core_113 = ~(input_a[7] ^ input_a[12]);
  assign popcount18_f88b_core_114 = input_a[0] & input_a[6];
  assign popcount18_f88b_core_115 = ~(input_a[0] ^ input_a[2]);
  assign popcount18_f88b_core_116 = ~input_a[5];
  assign popcount18_f88b_core_117 = input_a[2] & input_a[9];
  assign popcount18_f88b_core_118 = input_a[3] | input_a[15];
  assign popcount18_f88b_core_120 = ~input_a[12];
  assign popcount18_f88b_core_123_not = ~input_a[13];
  assign popcount18_f88b_core_124 = ~(input_a[16] & input_a[3]);
  assign popcount18_f88b_core_125 = ~(input_a[4] ^ input_a[4]);

  assign popcount18_f88b_out[0] = input_a[3];
  assign popcount18_f88b_out[1] = popcount18_f88b_core_057;
  assign popcount18_f88b_out[2] = popcount18_f88b_core_057;
  assign popcount18_f88b_out[3] = 1'b0;
  assign popcount18_f88b_out[4] = popcount18_f88b_core_059;
endmodule