// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.59324
// WCE=24.0
// EP=0.929865%
// Printed PDK parameters:
//  Area=42088520.0
//  Delay=69825784.0
//  Power=1900400.0

module popcount47_cbgb(input [46:0] input_a, output [5:0] popcount47_cbgb_out);
  wire popcount47_cbgb_core_051;
  wire popcount47_cbgb_core_052;
  wire popcount47_cbgb_core_053;
  wire popcount47_cbgb_core_054;
  wire popcount47_cbgb_core_055;
  wire popcount47_cbgb_core_056;
  wire popcount47_cbgb_core_057;
  wire popcount47_cbgb_core_058;
  wire popcount47_cbgb_core_060;
  wire popcount47_cbgb_core_063_not;
  wire popcount47_cbgb_core_065;
  wire popcount47_cbgb_core_067;
  wire popcount47_cbgb_core_068;
  wire popcount47_cbgb_core_069;
  wire popcount47_cbgb_core_073;
  wire popcount47_cbgb_core_074;
  wire popcount47_cbgb_core_075;
  wire popcount47_cbgb_core_076;
  wire popcount47_cbgb_core_077;
  wire popcount47_cbgb_core_078;
  wire popcount47_cbgb_core_079;
  wire popcount47_cbgb_core_080;
  wire popcount47_cbgb_core_081;
  wire popcount47_cbgb_core_082;
  wire popcount47_cbgb_core_083;
  wire popcount47_cbgb_core_084;
  wire popcount47_cbgb_core_086;
  wire popcount47_cbgb_core_088;
  wire popcount47_cbgb_core_089;
  wire popcount47_cbgb_core_092;
  wire popcount47_cbgb_core_093;
  wire popcount47_cbgb_core_095;
  wire popcount47_cbgb_core_099;
  wire popcount47_cbgb_core_100;
  wire popcount47_cbgb_core_103;
  wire popcount47_cbgb_core_107;
  wire popcount47_cbgb_core_108;
  wire popcount47_cbgb_core_109;
  wire popcount47_cbgb_core_110;
  wire popcount47_cbgb_core_117;
  wire popcount47_cbgb_core_118;
  wire popcount47_cbgb_core_120;
  wire popcount47_cbgb_core_123;
  wire popcount47_cbgb_core_124;
  wire popcount47_cbgb_core_125;
  wire popcount47_cbgb_core_130;
  wire popcount47_cbgb_core_133;
  wire popcount47_cbgb_core_134;
  wire popcount47_cbgb_core_136;
  wire popcount47_cbgb_core_138;
  wire popcount47_cbgb_core_139;
  wire popcount47_cbgb_core_140;
  wire popcount47_cbgb_core_141;
  wire popcount47_cbgb_core_142;
  wire popcount47_cbgb_core_144;
  wire popcount47_cbgb_core_146;
  wire popcount47_cbgb_core_149_not;
  wire popcount47_cbgb_core_151;
  wire popcount47_cbgb_core_152;
  wire popcount47_cbgb_core_153;
  wire popcount47_cbgb_core_155;
  wire popcount47_cbgb_core_157;
  wire popcount47_cbgb_core_158;
  wire popcount47_cbgb_core_163;
  wire popcount47_cbgb_core_166;
  wire popcount47_cbgb_core_167;
  wire popcount47_cbgb_core_168;
  wire popcount47_cbgb_core_169;
  wire popcount47_cbgb_core_171;
  wire popcount47_cbgb_core_172;
  wire popcount47_cbgb_core_173;
  wire popcount47_cbgb_core_175;
  wire popcount47_cbgb_core_176_not;
  wire popcount47_cbgb_core_178;
  wire popcount47_cbgb_core_179;
  wire popcount47_cbgb_core_180;
  wire popcount47_cbgb_core_181;
  wire popcount47_cbgb_core_182;
  wire popcount47_cbgb_core_183;
  wire popcount47_cbgb_core_184;
  wire popcount47_cbgb_core_185;
  wire popcount47_cbgb_core_186;
  wire popcount47_cbgb_core_187;
  wire popcount47_cbgb_core_188;
  wire popcount47_cbgb_core_190;
  wire popcount47_cbgb_core_192;
  wire popcount47_cbgb_core_194;
  wire popcount47_cbgb_core_195;
  wire popcount47_cbgb_core_197;
  wire popcount47_cbgb_core_198;
  wire popcount47_cbgb_core_199;
  wire popcount47_cbgb_core_200;
  wire popcount47_cbgb_core_201;
  wire popcount47_cbgb_core_202;
  wire popcount47_cbgb_core_203;
  wire popcount47_cbgb_core_204;
  wire popcount47_cbgb_core_205;
  wire popcount47_cbgb_core_206;
  wire popcount47_cbgb_core_208;
  wire popcount47_cbgb_core_209;
  wire popcount47_cbgb_core_211;
  wire popcount47_cbgb_core_213;
  wire popcount47_cbgb_core_217;
  wire popcount47_cbgb_core_220;
  wire popcount47_cbgb_core_221;
  wire popcount47_cbgb_core_222;
  wire popcount47_cbgb_core_227;
  wire popcount47_cbgb_core_230;
  wire popcount47_cbgb_core_232;
  wire popcount47_cbgb_core_233;
  wire popcount47_cbgb_core_236;
  wire popcount47_cbgb_core_238;
  wire popcount47_cbgb_core_243;
  wire popcount47_cbgb_core_244;
  wire popcount47_cbgb_core_245;
  wire popcount47_cbgb_core_246;
  wire popcount47_cbgb_core_247_not;
  wire popcount47_cbgb_core_249;
  wire popcount47_cbgb_core_250;
  wire popcount47_cbgb_core_254;
  wire popcount47_cbgb_core_257;
  wire popcount47_cbgb_core_258;
  wire popcount47_cbgb_core_259;
  wire popcount47_cbgb_core_260;
  wire popcount47_cbgb_core_261;
  wire popcount47_cbgb_core_263;
  wire popcount47_cbgb_core_265;
  wire popcount47_cbgb_core_267;
  wire popcount47_cbgb_core_268;
  wire popcount47_cbgb_core_269;
  wire popcount47_cbgb_core_272;
  wire popcount47_cbgb_core_273;
  wire popcount47_cbgb_core_277;
  wire popcount47_cbgb_core_279;
  wire popcount47_cbgb_core_281;
  wire popcount47_cbgb_core_282;
  wire popcount47_cbgb_core_283;
  wire popcount47_cbgb_core_284;
  wire popcount47_cbgb_core_288;
  wire popcount47_cbgb_core_289;
  wire popcount47_cbgb_core_290;
  wire popcount47_cbgb_core_291;
  wire popcount47_cbgb_core_292;
  wire popcount47_cbgb_core_293;
  wire popcount47_cbgb_core_296;
  wire popcount47_cbgb_core_299;
  wire popcount47_cbgb_core_300;
  wire popcount47_cbgb_core_306_not;
  wire popcount47_cbgb_core_309;
  wire popcount47_cbgb_core_310;
  wire popcount47_cbgb_core_316;
  wire popcount47_cbgb_core_317;
  wire popcount47_cbgb_core_318;
  wire popcount47_cbgb_core_319;
  wire popcount47_cbgb_core_323;
  wire popcount47_cbgb_core_324;
  wire popcount47_cbgb_core_325;
  wire popcount47_cbgb_core_326;
  wire popcount47_cbgb_core_327;
  wire popcount47_cbgb_core_328;
  wire popcount47_cbgb_core_329;
  wire popcount47_cbgb_core_330;
  wire popcount47_cbgb_core_331_not;
  wire popcount47_cbgb_core_338;
  wire popcount47_cbgb_core_339;
  wire popcount47_cbgb_core_344;
  wire popcount47_cbgb_core_345;
  wire popcount47_cbgb_core_347;
  wire popcount47_cbgb_core_348;
  wire popcount47_cbgb_core_350;
  wire popcount47_cbgb_core_352;
  wire popcount47_cbgb_core_353;
  wire popcount47_cbgb_core_354;
  wire popcount47_cbgb_core_355;
  wire popcount47_cbgb_core_356;
  wire popcount47_cbgb_core_357;
  wire popcount47_cbgb_core_358;
  wire popcount47_cbgb_core_359;
  wire popcount47_cbgb_core_360;
  wire popcount47_cbgb_core_361;
  wire popcount47_cbgb_core_362;
  wire popcount47_cbgb_core_363;
  wire popcount47_cbgb_core_364;
  wire popcount47_cbgb_core_365;
  wire popcount47_cbgb_core_366;
  wire popcount47_cbgb_core_367;
  wire popcount47_cbgb_core_369;
  wire popcount47_cbgb_core_371;
  wire popcount47_cbgb_core_372;

  assign popcount47_cbgb_core_051 = input_a[3] | input_a[4];
  assign popcount47_cbgb_core_052 = input_a[3] & input_a[4];
  assign popcount47_cbgb_core_053 = input_a[2] & popcount47_cbgb_core_051;
  assign popcount47_cbgb_core_054 = input_a[7] & popcount47_cbgb_core_051;
  assign popcount47_cbgb_core_055 = popcount47_cbgb_core_052 | popcount47_cbgb_core_054;
  assign popcount47_cbgb_core_056 = ~(input_a[31] | input_a[41]);
  assign popcount47_cbgb_core_057 = input_a[35] | input_a[34];
  assign popcount47_cbgb_core_058 = ~(input_a[6] | input_a[24]);
  assign popcount47_cbgb_core_060 = ~input_a[8];
  assign popcount47_cbgb_core_063_not = ~input_a[43];
  assign popcount47_cbgb_core_065 = input_a[29] | input_a[24];
  assign popcount47_cbgb_core_067 = input_a[35] & input_a[13];
  assign popcount47_cbgb_core_068 = input_a[25] | input_a[32];
  assign popcount47_cbgb_core_069 = ~input_a[8];
  assign popcount47_cbgb_core_073 = input_a[9] & input_a[10];
  assign popcount47_cbgb_core_074 = ~input_a[28];
  assign popcount47_cbgb_core_075 = input_a[8] & input_a[31];
  assign popcount47_cbgb_core_076 = popcount47_cbgb_core_073 | popcount47_cbgb_core_075;
  assign popcount47_cbgb_core_077 = ~(input_a[16] & input_a[37]);
  assign popcount47_cbgb_core_078 = popcount47_cbgb_core_068 ^ input_a[36];
  assign popcount47_cbgb_core_079 = input_a[40] & input_a[11];
  assign popcount47_cbgb_core_080 = popcount47_cbgb_core_067 ^ popcount47_cbgb_core_076;
  assign popcount47_cbgb_core_081 = popcount47_cbgb_core_067 & popcount47_cbgb_core_076;
  assign popcount47_cbgb_core_082 = popcount47_cbgb_core_080 ^ popcount47_cbgb_core_079;
  assign popcount47_cbgb_core_083 = popcount47_cbgb_core_080 & popcount47_cbgb_core_079;
  assign popcount47_cbgb_core_084 = popcount47_cbgb_core_081 | popcount47_cbgb_core_083;
  assign popcount47_cbgb_core_086 = input_a[41] | input_a[40];
  assign popcount47_cbgb_core_088 = ~(input_a[40] | input_a[40]);
  assign popcount47_cbgb_core_089 = ~input_a[34];
  assign popcount47_cbgb_core_092 = popcount47_cbgb_core_055 ^ popcount47_cbgb_core_082;
  assign popcount47_cbgb_core_093 = popcount47_cbgb_core_055 & popcount47_cbgb_core_082;
  assign popcount47_cbgb_core_095 = input_a[12] | input_a[39];
  assign popcount47_cbgb_core_099 = popcount47_cbgb_core_084 ^ popcount47_cbgb_core_093;
  assign popcount47_cbgb_core_100 = popcount47_cbgb_core_084 & popcount47_cbgb_core_093;
  assign popcount47_cbgb_core_103 = input_a[32] & input_a[18];
  assign popcount47_cbgb_core_107 = ~(input_a[14] | input_a[2]);
  assign popcount47_cbgb_core_108 = input_a[46] ^ input_a[6];
  assign popcount47_cbgb_core_109 = input_a[11] ^ input_a[41];
  assign popcount47_cbgb_core_110 = input_a[9] | input_a[39];
  assign popcount47_cbgb_core_117 = input_a[20] & input_a[21];
  assign popcount47_cbgb_core_118 = ~(input_a[8] & input_a[20]);
  assign popcount47_cbgb_core_120 = ~(input_a[36] | input_a[1]);
  assign popcount47_cbgb_core_123 = input_a[6] & input_a[43];
  assign popcount47_cbgb_core_124 = ~(input_a[28] ^ input_a[21]);
  assign popcount47_cbgb_core_125 = input_a[35] ^ input_a[2];
  assign popcount47_cbgb_core_130 = input_a[37] & input_a[20];
  assign popcount47_cbgb_core_133 = input_a[30] & input_a[11];
  assign popcount47_cbgb_core_134 = input_a[39] ^ input_a[17];
  assign popcount47_cbgb_core_136 = ~(input_a[9] & input_a[4]);
  assign popcount47_cbgb_core_138 = input_a[6] | input_a[17];
  assign popcount47_cbgb_core_139 = ~input_a[40];
  assign popcount47_cbgb_core_140 = ~(input_a[30] & input_a[24]);
  assign popcount47_cbgb_core_141 = ~(input_a[34] ^ input_a[39]);
  assign popcount47_cbgb_core_142 = input_a[22] ^ input_a[6];
  assign popcount47_cbgb_core_144 = ~(input_a[24] ^ input_a[12]);
  assign popcount47_cbgb_core_146 = input_a[8] & input_a[24];
  assign popcount47_cbgb_core_149_not = ~input_a[30];
  assign popcount47_cbgb_core_151 = input_a[39] ^ input_a[34];
  assign popcount47_cbgb_core_152 = ~input_a[24];
  assign popcount47_cbgb_core_153 = ~input_a[2];
  assign popcount47_cbgb_core_155 = input_a[42] ^ input_a[37];
  assign popcount47_cbgb_core_157 = popcount47_cbgb_core_123 ^ input_a[17];
  assign popcount47_cbgb_core_158 = popcount47_cbgb_core_123 & input_a[17];
  assign popcount47_cbgb_core_163 = ~input_a[30];
  assign popcount47_cbgb_core_166 = ~(input_a[14] | input_a[32]);
  assign popcount47_cbgb_core_167 = input_a[31] ^ input_a[39];
  assign popcount47_cbgb_core_168 = input_a[9] & input_a[8];
  assign popcount47_cbgb_core_169 = input_a[21] | input_a[33];
  assign popcount47_cbgb_core_171 = ~(input_a[4] | input_a[36]);
  assign popcount47_cbgb_core_172 = input_a[25] ^ input_a[23];
  assign popcount47_cbgb_core_173 = input_a[25] & input_a[41];
  assign popcount47_cbgb_core_175 = popcount47_cbgb_core_092 & popcount47_cbgb_core_157;
  assign popcount47_cbgb_core_176_not = ~popcount47_cbgb_core_173;
  assign popcount47_cbgb_core_178 = popcount47_cbgb_core_175 | popcount47_cbgb_core_173;
  assign popcount47_cbgb_core_179 = popcount47_cbgb_core_099 ^ popcount47_cbgb_core_158;
  assign popcount47_cbgb_core_180 = popcount47_cbgb_core_099 & popcount47_cbgb_core_158;
  assign popcount47_cbgb_core_181 = popcount47_cbgb_core_179 ^ popcount47_cbgb_core_178;
  assign popcount47_cbgb_core_182 = popcount47_cbgb_core_179 & popcount47_cbgb_core_178;
  assign popcount47_cbgb_core_183 = popcount47_cbgb_core_180 | popcount47_cbgb_core_182;
  assign popcount47_cbgb_core_184 = popcount47_cbgb_core_100 ^ popcount47_cbgb_core_169;
  assign popcount47_cbgb_core_185 = popcount47_cbgb_core_100 & popcount47_cbgb_core_169;
  assign popcount47_cbgb_core_186 = popcount47_cbgb_core_184 ^ popcount47_cbgb_core_183;
  assign popcount47_cbgb_core_187 = popcount47_cbgb_core_184 & popcount47_cbgb_core_183;
  assign popcount47_cbgb_core_188 = popcount47_cbgb_core_185 | popcount47_cbgb_core_187;
  assign popcount47_cbgb_core_190 = ~input_a[28];
  assign popcount47_cbgb_core_192 = input_a[43] ^ input_a[26];
  assign popcount47_cbgb_core_194 = ~input_a[38];
  assign popcount47_cbgb_core_195 = ~(input_a[1] ^ input_a[19]);
  assign popcount47_cbgb_core_197 = ~(input_a[34] ^ input_a[16]);
  assign popcount47_cbgb_core_198 = input_a[21] ^ input_a[4];
  assign popcount47_cbgb_core_199 = ~(input_a[29] ^ input_a[32]);
  assign popcount47_cbgb_core_200 = ~(input_a[31] | input_a[5]);
  assign popcount47_cbgb_core_201 = ~(input_a[12] | input_a[45]);
  assign popcount47_cbgb_core_202 = ~(input_a[40] | input_a[1]);
  assign popcount47_cbgb_core_203 = input_a[2] ^ input_a[9];
  assign popcount47_cbgb_core_204 = input_a[31] ^ input_a[16];
  assign popcount47_cbgb_core_205 = ~(input_a[27] | input_a[11]);
  assign popcount47_cbgb_core_206 = ~(input_a[8] | input_a[40]);
  assign popcount47_cbgb_core_208 = ~input_a[28];
  assign popcount47_cbgb_core_209 = ~(input_a[42] | input_a[13]);
  assign popcount47_cbgb_core_211 = ~(input_a[29] ^ input_a[45]);
  assign popcount47_cbgb_core_213 = ~(input_a[46] ^ input_a[31]);
  assign popcount47_cbgb_core_217 = ~(input_a[12] ^ input_a[31]);
  assign popcount47_cbgb_core_220 = input_a[30] | input_a[5];
  assign popcount47_cbgb_core_221 = input_a[41] | input_a[39];
  assign popcount47_cbgb_core_222 = ~input_a[30];
  assign popcount47_cbgb_core_227 = ~input_a[12];
  assign popcount47_cbgb_core_230 = input_a[36] | input_a[22];
  assign popcount47_cbgb_core_232 = ~(input_a[33] & input_a[38]);
  assign popcount47_cbgb_core_233 = input_a[12] ^ input_a[34];
  assign popcount47_cbgb_core_236 = ~(input_a[16] & input_a[33]);
  assign popcount47_cbgb_core_238 = ~(input_a[43] | input_a[22]);
  assign popcount47_cbgb_core_243 = popcount47_cbgb_core_206 & input_a[41];
  assign popcount47_cbgb_core_244 = ~(input_a[18] & input_a[4]);
  assign popcount47_cbgb_core_245 = input_a[24] & input_a[31];
  assign popcount47_cbgb_core_246 = input_a[0] & input_a[28];
  assign popcount47_cbgb_core_247_not = ~input_a[42];
  assign popcount47_cbgb_core_249 = ~input_a[32];
  assign popcount47_cbgb_core_250 = ~(input_a[14] | input_a[14]);
  assign popcount47_cbgb_core_254 = ~input_a[6];
  assign popcount47_cbgb_core_257 = input_a[28] | input_a[41];
  assign popcount47_cbgb_core_258 = ~(input_a[22] ^ input_a[38]);
  assign popcount47_cbgb_core_259 = ~(input_a[36] | input_a[44]);
  assign popcount47_cbgb_core_260 = input_a[22] ^ input_a[32];
  assign popcount47_cbgb_core_261 = ~(input_a[36] | input_a[10]);
  assign popcount47_cbgb_core_263 = input_a[34] ^ input_a[36];
  assign popcount47_cbgb_core_265 = ~(input_a[17] & input_a[28]);
  assign popcount47_cbgb_core_267 = ~input_a[36];
  assign popcount47_cbgb_core_268 = input_a[7] ^ input_a[11];
  assign popcount47_cbgb_core_269 = ~input_a[7];
  assign popcount47_cbgb_core_272 = input_a[7] ^ input_a[9];
  assign popcount47_cbgb_core_273 = popcount47_cbgb_core_263 ^ input_a[14];
  assign popcount47_cbgb_core_277 = input_a[28] | input_a[16];
  assign popcount47_cbgb_core_279 = input_a[32] | input_a[42];
  assign popcount47_cbgb_core_281 = input_a[13] ^ input_a[30];
  assign popcount47_cbgb_core_282 = ~input_a[34];
  assign popcount47_cbgb_core_283 = input_a[27] ^ input_a[33];
  assign popcount47_cbgb_core_284 = input_a[23] | input_a[0];
  assign popcount47_cbgb_core_288 = ~(input_a[29] | input_a[34]);
  assign popcount47_cbgb_core_289 = input_a[45] ^ input_a[34];
  assign popcount47_cbgb_core_290 = input_a[45] & input_a[46];
  assign popcount47_cbgb_core_291 = input_a[44] ^ popcount47_cbgb_core_289;
  assign popcount47_cbgb_core_292 = input_a[44] & popcount47_cbgb_core_289;
  assign popcount47_cbgb_core_293 = popcount47_cbgb_core_290 | popcount47_cbgb_core_292;
  assign popcount47_cbgb_core_296 = input_a[37] & input_a[30];
  assign popcount47_cbgb_core_299 = popcount47_cbgb_core_293 ^ popcount47_cbgb_core_296;
  assign popcount47_cbgb_core_300 = popcount47_cbgb_core_293 & popcount47_cbgb_core_296;
  assign popcount47_cbgb_core_306_not = ~input_a[39];
  assign popcount47_cbgb_core_309 = input_a[22] ^ popcount47_cbgb_core_299;
  assign popcount47_cbgb_core_310 = input_a[22] & popcount47_cbgb_core_299;
  assign popcount47_cbgb_core_316 = popcount47_cbgb_core_300 | popcount47_cbgb_core_310;
  assign popcount47_cbgb_core_317 = input_a[13] | input_a[24];
  assign popcount47_cbgb_core_318 = input_a[21] & input_a[29];
  assign popcount47_cbgb_core_319 = input_a[25] | input_a[13];
  assign popcount47_cbgb_core_323 = ~(input_a[5] & input_a[7]);
  assign popcount47_cbgb_core_324 = input_a[9] & input_a[36];
  assign popcount47_cbgb_core_325 = input_a[5] & input_a[18];
  assign popcount47_cbgb_core_326 = popcount47_cbgb_core_246 | popcount47_cbgb_core_309;
  assign popcount47_cbgb_core_327 = ~(input_a[19] | input_a[18]);
  assign popcount47_cbgb_core_328 = popcount47_cbgb_core_326 | popcount47_cbgb_core_325;
  assign popcount47_cbgb_core_329 = ~(input_a[0] | input_a[10]);
  assign popcount47_cbgb_core_330 = input_a[18] ^ input_a[22];
  assign popcount47_cbgb_core_331_not = ~popcount47_cbgb_core_316;
  assign popcount47_cbgb_core_338 = input_a[26] ^ popcount47_cbgb_core_316;
  assign popcount47_cbgb_core_339 = input_a[26] & popcount47_cbgb_core_316;
  assign popcount47_cbgb_core_344 = input_a[43] | input_a[0];
  assign popcount47_cbgb_core_345 = input_a[37] ^ input_a[12];
  assign popcount47_cbgb_core_347 = ~(input_a[24] & input_a[43]);
  assign popcount47_cbgb_core_348 = popcount47_cbgb_core_176_not ^ popcount47_cbgb_core_328;
  assign popcount47_cbgb_core_350 = ~popcount47_cbgb_core_348;
  assign popcount47_cbgb_core_352 = popcount47_cbgb_core_176_not | popcount47_cbgb_core_348;
  assign popcount47_cbgb_core_353 = popcount47_cbgb_core_181 ^ popcount47_cbgb_core_331_not;
  assign popcount47_cbgb_core_354 = popcount47_cbgb_core_181 & popcount47_cbgb_core_331_not;
  assign popcount47_cbgb_core_355 = popcount47_cbgb_core_353 ^ popcount47_cbgb_core_352;
  assign popcount47_cbgb_core_356 = popcount47_cbgb_core_353 & popcount47_cbgb_core_352;
  assign popcount47_cbgb_core_357 = popcount47_cbgb_core_354 | popcount47_cbgb_core_356;
  assign popcount47_cbgb_core_358 = popcount47_cbgb_core_186 ^ popcount47_cbgb_core_338;
  assign popcount47_cbgb_core_359 = popcount47_cbgb_core_186 & popcount47_cbgb_core_338;
  assign popcount47_cbgb_core_360 = popcount47_cbgb_core_358 ^ popcount47_cbgb_core_357;
  assign popcount47_cbgb_core_361 = popcount47_cbgb_core_358 & popcount47_cbgb_core_357;
  assign popcount47_cbgb_core_362 = popcount47_cbgb_core_359 | popcount47_cbgb_core_361;
  assign popcount47_cbgb_core_363 = popcount47_cbgb_core_188 ^ popcount47_cbgb_core_339;
  assign popcount47_cbgb_core_364 = popcount47_cbgb_core_188 & popcount47_cbgb_core_339;
  assign popcount47_cbgb_core_365 = popcount47_cbgb_core_363 ^ popcount47_cbgb_core_362;
  assign popcount47_cbgb_core_366 = popcount47_cbgb_core_363 & popcount47_cbgb_core_362;
  assign popcount47_cbgb_core_367 = popcount47_cbgb_core_364 | popcount47_cbgb_core_366;
  assign popcount47_cbgb_core_369 = ~input_a[2];
  assign popcount47_cbgb_core_371 = input_a[15] | input_a[31];
  assign popcount47_cbgb_core_372 = input_a[22] | input_a[9];

  assign popcount47_cbgb_out[0] = input_a[19];
  assign popcount47_cbgb_out[1] = popcount47_cbgb_core_350;
  assign popcount47_cbgb_out[2] = popcount47_cbgb_core_355;
  assign popcount47_cbgb_out[3] = popcount47_cbgb_core_360;
  assign popcount47_cbgb_out[4] = popcount47_cbgb_core_365;
  assign popcount47_cbgb_out[5] = popcount47_cbgb_core_367;
endmodule