// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.49608
// WCE=9.0
// EP=0.792889%
// Printed PDK parameters:
//  Area=37174084.0
//  Delay=64488444.0
//  Power=1971000.0

module popcount30_dedb(input [29:0] input_a, output [4:0] popcount30_dedb_out);
  wire popcount30_dedb_core_032;
  wire popcount30_dedb_core_034_not;
  wire popcount30_dedb_core_036;
  wire popcount30_dedb_core_039;
  wire popcount30_dedb_core_040;
  wire popcount30_dedb_core_041;
  wire popcount30_dedb_core_042;
  wire popcount30_dedb_core_043;
  wire popcount30_dedb_core_044;
  wire popcount30_dedb_core_045;
  wire popcount30_dedb_core_046;
  wire popcount30_dedb_core_047;
  wire popcount30_dedb_core_049_not;
  wire popcount30_dedb_core_050;
  wire popcount30_dedb_core_051;
  wire popcount30_dedb_core_052;
  wire popcount30_dedb_core_057;
  wire popcount30_dedb_core_058;
  wire popcount30_dedb_core_059;
  wire popcount30_dedb_core_060;
  wire popcount30_dedb_core_061;
  wire popcount30_dedb_core_062;
  wire popcount30_dedb_core_064;
  wire popcount30_dedb_core_065;
  wire popcount30_dedb_core_066;
  wire popcount30_dedb_core_068;
  wire popcount30_dedb_core_069;
  wire popcount30_dedb_core_070;
  wire popcount30_dedb_core_071;
  wire popcount30_dedb_core_073;
  wire popcount30_dedb_core_074;
  wire popcount30_dedb_core_075;
  wire popcount30_dedb_core_076;
  wire popcount30_dedb_core_077;
  wire popcount30_dedb_core_078;
  wire popcount30_dedb_core_079;
  wire popcount30_dedb_core_081;
  wire popcount30_dedb_core_082;
  wire popcount30_dedb_core_083;
  wire popcount30_dedb_core_084;
  wire popcount30_dedb_core_085;
  wire popcount30_dedb_core_086;
  wire popcount30_dedb_core_088;
  wire popcount30_dedb_core_091;
  wire popcount30_dedb_core_094;
  wire popcount30_dedb_core_095;
  wire popcount30_dedb_core_096;
  wire popcount30_dedb_core_097;
  wire popcount30_dedb_core_099;
  wire popcount30_dedb_core_101;
  wire popcount30_dedb_core_102;
  wire popcount30_dedb_core_104;
  wire popcount30_dedb_core_105;
  wire popcount30_dedb_core_106;
  wire popcount30_dedb_core_108;
  wire popcount30_dedb_core_110;
  wire popcount30_dedb_core_111;
  wire popcount30_dedb_core_112;
  wire popcount30_dedb_core_113;
  wire popcount30_dedb_core_114;
  wire popcount30_dedb_core_115;
  wire popcount30_dedb_core_116;
  wire popcount30_dedb_core_117;
  wire popcount30_dedb_core_118;
  wire popcount30_dedb_core_119;
  wire popcount30_dedb_core_120;
  wire popcount30_dedb_core_121;
  wire popcount30_dedb_core_123;
  wire popcount30_dedb_core_125;
  wire popcount30_dedb_core_128;
  wire popcount30_dedb_core_130;
  wire popcount30_dedb_core_131;
  wire popcount30_dedb_core_132;
  wire popcount30_dedb_core_133;
  wire popcount30_dedb_core_134;
  wire popcount30_dedb_core_135;
  wire popcount30_dedb_core_137;
  wire popcount30_dedb_core_139;
  wire popcount30_dedb_core_142;
  wire popcount30_dedb_core_143;
  wire popcount30_dedb_core_144;
  wire popcount30_dedb_core_145;
  wire popcount30_dedb_core_146;
  wire popcount30_dedb_core_148;
  wire popcount30_dedb_core_150;
  wire popcount30_dedb_core_151;
  wire popcount30_dedb_core_152;
  wire popcount30_dedb_core_153;
  wire popcount30_dedb_core_154;
  wire popcount30_dedb_core_156;
  wire popcount30_dedb_core_157;
  wire popcount30_dedb_core_158;
  wire popcount30_dedb_core_160;
  wire popcount30_dedb_core_161;
  wire popcount30_dedb_core_163;
  wire popcount30_dedb_core_165;
  wire popcount30_dedb_core_167;
  wire popcount30_dedb_core_168;
  wire popcount30_dedb_core_169;
  wire popcount30_dedb_core_173;
  wire popcount30_dedb_core_175;
  wire popcount30_dedb_core_176;
  wire popcount30_dedb_core_177;
  wire popcount30_dedb_core_178;
  wire popcount30_dedb_core_179;
  wire popcount30_dedb_core_180;
  wire popcount30_dedb_core_181;
  wire popcount30_dedb_core_182;
  wire popcount30_dedb_core_183;
  wire popcount30_dedb_core_184;
  wire popcount30_dedb_core_185;
  wire popcount30_dedb_core_186;
  wire popcount30_dedb_core_188;
  wire popcount30_dedb_core_193;
  wire popcount30_dedb_core_194;
  wire popcount30_dedb_core_195;
  wire popcount30_dedb_core_196;
  wire popcount30_dedb_core_197;
  wire popcount30_dedb_core_198;
  wire popcount30_dedb_core_199;
  wire popcount30_dedb_core_200;
  wire popcount30_dedb_core_201;
  wire popcount30_dedb_core_202;
  wire popcount30_dedb_core_203;
  wire popcount30_dedb_core_204;
  wire popcount30_dedb_core_205;
  wire popcount30_dedb_core_206;
  wire popcount30_dedb_core_207;
  wire popcount30_dedb_core_208;
  wire popcount30_dedb_core_213;

  assign popcount30_dedb_core_032 = ~(input_a[9] | input_a[16]);
  assign popcount30_dedb_core_034_not = ~input_a[19];
  assign popcount30_dedb_core_036 = input_a[14] | input_a[23];
  assign popcount30_dedb_core_039 = input_a[3] & input_a[4];
  assign popcount30_dedb_core_040 = input_a[22] & input_a[16];
  assign popcount30_dedb_core_041 = input_a[27] & input_a[28];
  assign popcount30_dedb_core_042 = input_a[9] ^ input_a[29];
  assign popcount30_dedb_core_043 = input_a[18] & input_a[2];
  assign popcount30_dedb_core_044 = popcount30_dedb_core_039 ^ popcount30_dedb_core_041;
  assign popcount30_dedb_core_045 = popcount30_dedb_core_039 & popcount30_dedb_core_041;
  assign popcount30_dedb_core_046 = popcount30_dedb_core_044 | popcount30_dedb_core_043;
  assign popcount30_dedb_core_047 = ~(input_a[9] ^ input_a[24]);
  assign popcount30_dedb_core_049_not = ~input_a[6];
  assign popcount30_dedb_core_050 = ~(input_a[26] | input_a[5]);
  assign popcount30_dedb_core_051 = popcount30_dedb_core_036 ^ popcount30_dedb_core_046;
  assign popcount30_dedb_core_052 = popcount30_dedb_core_036 & popcount30_dedb_core_046;
  assign popcount30_dedb_core_057 = input_a[10] | input_a[4];
  assign popcount30_dedb_core_058 = popcount30_dedb_core_045 | popcount30_dedb_core_052;
  assign popcount30_dedb_core_059 = ~input_a[13];
  assign popcount30_dedb_core_060 = ~(input_a[27] | input_a[7]);
  assign popcount30_dedb_core_061 = input_a[26] | input_a[3];
  assign popcount30_dedb_core_062 = input_a[24] ^ input_a[22];
  assign popcount30_dedb_core_064 = input_a[9] ^ input_a[24];
  assign popcount30_dedb_core_065 = ~input_a[9];
  assign popcount30_dedb_core_066 = ~input_a[1];
  assign popcount30_dedb_core_068 = ~(input_a[10] ^ input_a[4]);
  assign popcount30_dedb_core_069 = input_a[0] | input_a[26];
  assign popcount30_dedb_core_070 = input_a[21] ^ input_a[23];
  assign popcount30_dedb_core_071 = ~(input_a[17] | input_a[29]);
  assign popcount30_dedb_core_073 = input_a[5] & input_a[8];
  assign popcount30_dedb_core_074 = input_a[6] & input_a[9];
  assign popcount30_dedb_core_075 = input_a[24] & input_a[25];
  assign popcount30_dedb_core_076 = ~(input_a[9] ^ input_a[2]);
  assign popcount30_dedb_core_077 = ~(input_a[2] | input_a[11]);
  assign popcount30_dedb_core_078 = popcount30_dedb_core_073 | input_a[24];
  assign popcount30_dedb_core_079 = ~input_a[12];
  assign popcount30_dedb_core_081 = ~(input_a[17] & input_a[17]);
  assign popcount30_dedb_core_082 = input_a[3] & input_a[26];
  assign popcount30_dedb_core_083 = input_a[21] & input_a[19];
  assign popcount30_dedb_core_084 = ~(input_a[24] & input_a[23]);
  assign popcount30_dedb_core_085 = ~(popcount30_dedb_core_069 & popcount30_dedb_core_078);
  assign popcount30_dedb_core_086 = popcount30_dedb_core_069 & popcount30_dedb_core_078;
  assign popcount30_dedb_core_088 = input_a[26] | input_a[23];
  assign popcount30_dedb_core_091 = input_a[9] | input_a[5];
  assign popcount30_dedb_core_094 = input_a[4] | input_a[21];
  assign popcount30_dedb_core_095 = ~(input_a[17] & input_a[15]);
  assign popcount30_dedb_core_096 = ~(input_a[8] ^ input_a[10]);
  assign popcount30_dedb_core_097 = popcount30_dedb_core_051 ^ popcount30_dedb_core_085;
  assign popcount30_dedb_core_099 = ~popcount30_dedb_core_097;
  assign popcount30_dedb_core_101 = popcount30_dedb_core_051 | popcount30_dedb_core_097;
  assign popcount30_dedb_core_102 = popcount30_dedb_core_058 ^ popcount30_dedb_core_086;
  assign popcount30_dedb_core_104 = popcount30_dedb_core_102 ^ popcount30_dedb_core_101;
  assign popcount30_dedb_core_105 = popcount30_dedb_core_102 & popcount30_dedb_core_101;
  assign popcount30_dedb_core_106 = popcount30_dedb_core_058 | popcount30_dedb_core_105;
  assign popcount30_dedb_core_108 = ~(input_a[2] | input_a[20]);
  assign popcount30_dedb_core_110 = ~input_a[8];
  assign popcount30_dedb_core_111 = input_a[24] & input_a[20];
  assign popcount30_dedb_core_112 = ~input_a[8];
  assign popcount30_dedb_core_113 = input_a[10] & input_a[17];
  assign popcount30_dedb_core_114 = input_a[13] & input_a[5];
  assign popcount30_dedb_core_115 = input_a[11] & input_a[6];
  assign popcount30_dedb_core_116 = popcount30_dedb_core_113 | popcount30_dedb_core_115;
  assign popcount30_dedb_core_117 = ~(input_a[29] ^ input_a[25]);
  assign popcount30_dedb_core_118 = ~(input_a[23] ^ input_a[20]);
  assign popcount30_dedb_core_119 = input_a[13] & input_a[20];
  assign popcount30_dedb_core_120 = ~(input_a[8] ^ input_a[6]);
  assign popcount30_dedb_core_121 = input_a[13] | input_a[6];
  assign popcount30_dedb_core_123 = ~(input_a[23] | input_a[29]);
  assign popcount30_dedb_core_125 = ~(input_a[22] | input_a[26]);
  assign popcount30_dedb_core_128 = input_a[5] & input_a[11];
  assign popcount30_dedb_core_130 = ~input_a[5];
  assign popcount30_dedb_core_131 = popcount30_dedb_core_116 ^ popcount30_dedb_core_119;
  assign popcount30_dedb_core_132 = popcount30_dedb_core_116 & popcount30_dedb_core_119;
  assign popcount30_dedb_core_133 = popcount30_dedb_core_131 ^ input_a[25];
  assign popcount30_dedb_core_134 = popcount30_dedb_core_131 & input_a[25];
  assign popcount30_dedb_core_135 = popcount30_dedb_core_132 | popcount30_dedb_core_134;
  assign popcount30_dedb_core_137 = input_a[14] | input_a[1];
  assign popcount30_dedb_core_139 = input_a[28] | input_a[19];
  assign popcount30_dedb_core_142 = input_a[19] & input_a[9];
  assign popcount30_dedb_core_143 = input_a[8] | input_a[13];
  assign popcount30_dedb_core_144 = ~(input_a[13] | input_a[12]);
  assign popcount30_dedb_core_145 = input_a[22] & input_a[16];
  assign popcount30_dedb_core_146 = input_a[2] & input_a[12];
  assign popcount30_dedb_core_148 = input_a[14] | input_a[23];
  assign popcount30_dedb_core_150 = ~(input_a[18] & input_a[20]);
  assign popcount30_dedb_core_151 = ~(input_a[14] ^ input_a[9]);
  assign popcount30_dedb_core_152 = input_a[28] ^ input_a[14];
  assign popcount30_dedb_core_153 = input_a[17] | input_a[17];
  assign popcount30_dedb_core_154 = ~(input_a[20] ^ input_a[2]);
  assign popcount30_dedb_core_156 = input_a[17] | input_a[12];
  assign popcount30_dedb_core_157 = ~(input_a[26] & input_a[8]);
  assign popcount30_dedb_core_158 = input_a[9] & input_a[5];
  assign popcount30_dedb_core_160 = ~input_a[15];
  assign popcount30_dedb_core_161 = ~(input_a[26] & input_a[19]);
  assign popcount30_dedb_core_163 = input_a[7] | input_a[29];
  assign popcount30_dedb_core_165 = ~popcount30_dedb_core_142;
  assign popcount30_dedb_core_167 = popcount30_dedb_core_165 ^ popcount30_dedb_core_145;
  assign popcount30_dedb_core_168 = input_a[22] & popcount30_dedb_core_145;
  assign popcount30_dedb_core_169 = popcount30_dedb_core_142 | popcount30_dedb_core_168;
  assign popcount30_dedb_core_173 = input_a[6] | input_a[0];
  assign popcount30_dedb_core_175 = input_a[13] & input_a[5];
  assign popcount30_dedb_core_176 = input_a[12] & popcount30_dedb_core_163;
  assign popcount30_dedb_core_177 = popcount30_dedb_core_133 ^ popcount30_dedb_core_167;
  assign popcount30_dedb_core_178 = popcount30_dedb_core_133 & popcount30_dedb_core_167;
  assign popcount30_dedb_core_179 = popcount30_dedb_core_177 ^ popcount30_dedb_core_176;
  assign popcount30_dedb_core_180 = popcount30_dedb_core_177 & popcount30_dedb_core_176;
  assign popcount30_dedb_core_181 = popcount30_dedb_core_178 | popcount30_dedb_core_180;
  assign popcount30_dedb_core_182 = popcount30_dedb_core_135 ^ popcount30_dedb_core_169;
  assign popcount30_dedb_core_183 = popcount30_dedb_core_135 & popcount30_dedb_core_169;
  assign popcount30_dedb_core_184 = popcount30_dedb_core_182 ^ popcount30_dedb_core_181;
  assign popcount30_dedb_core_185 = popcount30_dedb_core_182 & popcount30_dedb_core_181;
  assign popcount30_dedb_core_186 = popcount30_dedb_core_183 | popcount30_dedb_core_185;
  assign popcount30_dedb_core_188 = ~(input_a[0] & input_a[18]);
  assign popcount30_dedb_core_193 = input_a[21] & input_a[1];
  assign popcount30_dedb_core_194 = popcount30_dedb_core_099 ^ popcount30_dedb_core_179;
  assign popcount30_dedb_core_195 = popcount30_dedb_core_099 & popcount30_dedb_core_179;
  assign popcount30_dedb_core_196 = popcount30_dedb_core_194 ^ popcount30_dedb_core_193;
  assign popcount30_dedb_core_197 = popcount30_dedb_core_194 & popcount30_dedb_core_193;
  assign popcount30_dedb_core_198 = popcount30_dedb_core_195 | popcount30_dedb_core_197;
  assign popcount30_dedb_core_199 = popcount30_dedb_core_104 ^ popcount30_dedb_core_184;
  assign popcount30_dedb_core_200 = popcount30_dedb_core_104 & popcount30_dedb_core_184;
  assign popcount30_dedb_core_201 = popcount30_dedb_core_199 ^ popcount30_dedb_core_198;
  assign popcount30_dedb_core_202 = popcount30_dedb_core_199 & popcount30_dedb_core_198;
  assign popcount30_dedb_core_203 = popcount30_dedb_core_200 | popcount30_dedb_core_202;
  assign popcount30_dedb_core_204 = popcount30_dedb_core_106 ^ popcount30_dedb_core_186;
  assign popcount30_dedb_core_205 = popcount30_dedb_core_106 & popcount30_dedb_core_186;
  assign popcount30_dedb_core_206 = popcount30_dedb_core_204 ^ popcount30_dedb_core_203;
  assign popcount30_dedb_core_207 = popcount30_dedb_core_204 & popcount30_dedb_core_203;
  assign popcount30_dedb_core_208 = popcount30_dedb_core_205 | popcount30_dedb_core_207;
  assign popcount30_dedb_core_213 = ~(input_a[9] & input_a[1]);

  assign popcount30_dedb_out[0] = popcount30_dedb_core_206;
  assign popcount30_dedb_out[1] = popcount30_dedb_core_196;
  assign popcount30_dedb_out[2] = popcount30_dedb_core_201;
  assign popcount30_dedb_out[3] = popcount30_dedb_core_206;
  assign popcount30_dedb_out[4] = popcount30_dedb_core_208;
endmodule