// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.55409
// WCE=14.0
// EP=0.8831%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_jxwu(input [24:0] input_a, output [4:0] popcount25_jxwu_out);
  wire popcount25_jxwu_core_027;
  wire popcount25_jxwu_core_030;
  wire popcount25_jxwu_core_032;
  wire popcount25_jxwu_core_033;
  wire popcount25_jxwu_core_034;
  wire popcount25_jxwu_core_035;
  wire popcount25_jxwu_core_036;
  wire popcount25_jxwu_core_039;
  wire popcount25_jxwu_core_040;
  wire popcount25_jxwu_core_041;
  wire popcount25_jxwu_core_045;
  wire popcount25_jxwu_core_047;
  wire popcount25_jxwu_core_049;
  wire popcount25_jxwu_core_050;
  wire popcount25_jxwu_core_054;
  wire popcount25_jxwu_core_057;
  wire popcount25_jxwu_core_058;
  wire popcount25_jxwu_core_060;
  wire popcount25_jxwu_core_061;
  wire popcount25_jxwu_core_065;
  wire popcount25_jxwu_core_066;
  wire popcount25_jxwu_core_068;
  wire popcount25_jxwu_core_070;
  wire popcount25_jxwu_core_072;
  wire popcount25_jxwu_core_075;
  wire popcount25_jxwu_core_076;
  wire popcount25_jxwu_core_077;
  wire popcount25_jxwu_core_080_not;
  wire popcount25_jxwu_core_081;
  wire popcount25_jxwu_core_082;
  wire popcount25_jxwu_core_083;
  wire popcount25_jxwu_core_086;
  wire popcount25_jxwu_core_087;
  wire popcount25_jxwu_core_088;
  wire popcount25_jxwu_core_089;
  wire popcount25_jxwu_core_093;
  wire popcount25_jxwu_core_098_not;
  wire popcount25_jxwu_core_099;
  wire popcount25_jxwu_core_100;
  wire popcount25_jxwu_core_102;
  wire popcount25_jxwu_core_103_not;
  wire popcount25_jxwu_core_104;
  wire popcount25_jxwu_core_106;
  wire popcount25_jxwu_core_107;
  wire popcount25_jxwu_core_109;
  wire popcount25_jxwu_core_110;
  wire popcount25_jxwu_core_111;
  wire popcount25_jxwu_core_113;
  wire popcount25_jxwu_core_116;
  wire popcount25_jxwu_core_117;
  wire popcount25_jxwu_core_119;
  wire popcount25_jxwu_core_121;
  wire popcount25_jxwu_core_122;
  wire popcount25_jxwu_core_123;
  wire popcount25_jxwu_core_125;
  wire popcount25_jxwu_core_126;
  wire popcount25_jxwu_core_128;
  wire popcount25_jxwu_core_129_not;
  wire popcount25_jxwu_core_130;
  wire popcount25_jxwu_core_132;
  wire popcount25_jxwu_core_135;
  wire popcount25_jxwu_core_136;
  wire popcount25_jxwu_core_137;
  wire popcount25_jxwu_core_138;
  wire popcount25_jxwu_core_139;
  wire popcount25_jxwu_core_141;
  wire popcount25_jxwu_core_145;
  wire popcount25_jxwu_core_147;
  wire popcount25_jxwu_core_148;
  wire popcount25_jxwu_core_150;
  wire popcount25_jxwu_core_152;
  wire popcount25_jxwu_core_153;
  wire popcount25_jxwu_core_157;
  wire popcount25_jxwu_core_159;
  wire popcount25_jxwu_core_160;
  wire popcount25_jxwu_core_163;
  wire popcount25_jxwu_core_164;
  wire popcount25_jxwu_core_165;
  wire popcount25_jxwu_core_166;
  wire popcount25_jxwu_core_170;
  wire popcount25_jxwu_core_171;
  wire popcount25_jxwu_core_174;
  wire popcount25_jxwu_core_176;
  wire popcount25_jxwu_core_178;
  wire popcount25_jxwu_core_179;
  wire popcount25_jxwu_core_180;
  wire popcount25_jxwu_core_181;
  wire popcount25_jxwu_core_182;
  wire popcount25_jxwu_core_183;

  assign popcount25_jxwu_core_027 = ~(input_a[20] | input_a[3]);
  assign popcount25_jxwu_core_030 = input_a[3] | input_a[21];
  assign popcount25_jxwu_core_032 = ~(input_a[7] & input_a[22]);
  assign popcount25_jxwu_core_033 = input_a[6] | input_a[4];
  assign popcount25_jxwu_core_034 = ~(input_a[7] & input_a[11]);
  assign popcount25_jxwu_core_035 = ~(input_a[21] ^ input_a[14]);
  assign popcount25_jxwu_core_036 = ~input_a[23];
  assign popcount25_jxwu_core_039 = input_a[21] & input_a[4];
  assign popcount25_jxwu_core_040 = ~(input_a[3] | input_a[17]);
  assign popcount25_jxwu_core_041 = input_a[3] & input_a[6];
  assign popcount25_jxwu_core_045 = ~input_a[16];
  assign popcount25_jxwu_core_047 = input_a[21] | input_a[21];
  assign popcount25_jxwu_core_049 = input_a[5] & input_a[15];
  assign popcount25_jxwu_core_050 = input_a[4] | input_a[8];
  assign popcount25_jxwu_core_054 = ~(input_a[11] ^ input_a[10]);
  assign popcount25_jxwu_core_057 = input_a[7] ^ input_a[21];
  assign popcount25_jxwu_core_058 = input_a[22] ^ input_a[4];
  assign popcount25_jxwu_core_060 = input_a[13] | input_a[22];
  assign popcount25_jxwu_core_061 = input_a[6] | input_a[22];
  assign popcount25_jxwu_core_065 = ~(input_a[19] ^ input_a[13]);
  assign popcount25_jxwu_core_066 = input_a[2] | input_a[1];
  assign popcount25_jxwu_core_068 = ~(input_a[17] | input_a[13]);
  assign popcount25_jxwu_core_070 = ~(input_a[16] | input_a[24]);
  assign popcount25_jxwu_core_072 = input_a[24] | input_a[2];
  assign popcount25_jxwu_core_075 = input_a[11] | input_a[12];
  assign popcount25_jxwu_core_076 = ~(input_a[10] & input_a[5]);
  assign popcount25_jxwu_core_077 = input_a[7] | input_a[8];
  assign popcount25_jxwu_core_080_not = ~input_a[8];
  assign popcount25_jxwu_core_081 = input_a[0] & input_a[7];
  assign popcount25_jxwu_core_082 = ~(input_a[4] | input_a[21]);
  assign popcount25_jxwu_core_083 = ~(input_a[11] ^ input_a[18]);
  assign popcount25_jxwu_core_086 = ~(input_a[9] & input_a[0]);
  assign popcount25_jxwu_core_087 = input_a[4] ^ input_a[22];
  assign popcount25_jxwu_core_088 = ~(input_a[1] & input_a[14]);
  assign popcount25_jxwu_core_089 = ~input_a[3];
  assign popcount25_jxwu_core_093 = input_a[3] | input_a[15];
  assign popcount25_jxwu_core_098_not = ~input_a[8];
  assign popcount25_jxwu_core_099 = ~(input_a[18] | input_a[12]);
  assign popcount25_jxwu_core_100 = input_a[14] | input_a[0];
  assign popcount25_jxwu_core_102 = ~(input_a[5] ^ input_a[21]);
  assign popcount25_jxwu_core_103_not = ~input_a[19];
  assign popcount25_jxwu_core_104 = ~(input_a[2] | input_a[12]);
  assign popcount25_jxwu_core_106 = ~input_a[15];
  assign popcount25_jxwu_core_107 = input_a[2] | input_a[17];
  assign popcount25_jxwu_core_109 = ~input_a[1];
  assign popcount25_jxwu_core_110 = input_a[1] & input_a[19];
  assign popcount25_jxwu_core_111 = ~input_a[15];
  assign popcount25_jxwu_core_113 = ~(input_a[14] | input_a[10]);
  assign popcount25_jxwu_core_116 = input_a[6] ^ input_a[9];
  assign popcount25_jxwu_core_117 = input_a[4] ^ input_a[19];
  assign popcount25_jxwu_core_119 = ~(input_a[14] | input_a[1]);
  assign popcount25_jxwu_core_121 = input_a[12] & input_a[23];
  assign popcount25_jxwu_core_122 = ~input_a[13];
  assign popcount25_jxwu_core_123 = input_a[3] | input_a[10];
  assign popcount25_jxwu_core_125 = input_a[11] ^ input_a[2];
  assign popcount25_jxwu_core_126 = ~input_a[16];
  assign popcount25_jxwu_core_128 = input_a[0] & input_a[17];
  assign popcount25_jxwu_core_129_not = ~input_a[13];
  assign popcount25_jxwu_core_130 = input_a[7] | input_a[18];
  assign popcount25_jxwu_core_132 = ~input_a[17];
  assign popcount25_jxwu_core_135 = input_a[16] | input_a[24];
  assign popcount25_jxwu_core_136 = input_a[10] & input_a[17];
  assign popcount25_jxwu_core_137 = ~(input_a[3] | input_a[24]);
  assign popcount25_jxwu_core_138 = input_a[21] | input_a[23];
  assign popcount25_jxwu_core_139 = ~(input_a[24] | input_a[18]);
  assign popcount25_jxwu_core_141 = ~(input_a[14] | input_a[23]);
  assign popcount25_jxwu_core_145 = ~(input_a[6] | input_a[22]);
  assign popcount25_jxwu_core_147 = ~input_a[19];
  assign popcount25_jxwu_core_148 = input_a[2] & input_a[7];
  assign popcount25_jxwu_core_150 = input_a[15] ^ input_a[3];
  assign popcount25_jxwu_core_152 = ~input_a[18];
  assign popcount25_jxwu_core_153 = input_a[17] ^ input_a[24];
  assign popcount25_jxwu_core_157 = input_a[13] ^ input_a[13];
  assign popcount25_jxwu_core_159 = input_a[22] & input_a[6];
  assign popcount25_jxwu_core_160 = ~input_a[18];
  assign popcount25_jxwu_core_163 = input_a[11] & input_a[14];
  assign popcount25_jxwu_core_164 = input_a[4] ^ input_a[23];
  assign popcount25_jxwu_core_165 = ~(input_a[8] ^ input_a[9]);
  assign popcount25_jxwu_core_166 = input_a[23] | input_a[17];
  assign popcount25_jxwu_core_170 = ~(input_a[20] | input_a[13]);
  assign popcount25_jxwu_core_171 = input_a[17] & input_a[3];
  assign popcount25_jxwu_core_174 = input_a[4] & input_a[12];
  assign popcount25_jxwu_core_176 = ~input_a[6];
  assign popcount25_jxwu_core_178 = ~input_a[10];
  assign popcount25_jxwu_core_179 = input_a[14] | input_a[12];
  assign popcount25_jxwu_core_180 = ~(input_a[23] | input_a[9]);
  assign popcount25_jxwu_core_181 = ~(input_a[24] & input_a[1]);
  assign popcount25_jxwu_core_182 = ~(input_a[6] | input_a[21]);
  assign popcount25_jxwu_core_183 = ~(input_a[10] & input_a[20]);

  assign popcount25_jxwu_out[0] = input_a[17];
  assign popcount25_jxwu_out[1] = 1'b1;
  assign popcount25_jxwu_out[2] = 1'b0;
  assign popcount25_jxwu_out[3] = 1'b1;
  assign popcount25_jxwu_out[4] = 1'b0;
endmodule