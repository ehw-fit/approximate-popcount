// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.50742
// WCE=20.0
// EP=0.992607%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_59hv(input [22:0] input_a, output [4:0] popcount23_59hv_out);
  wire popcount23_59hv_core_026;
  wire popcount23_59hv_core_027;
  wire popcount23_59hv_core_029;
  wire popcount23_59hv_core_031;
  wire popcount23_59hv_core_032;
  wire popcount23_59hv_core_035;
  wire popcount23_59hv_core_036_not;
  wire popcount23_59hv_core_039;
  wire popcount23_59hv_core_044;
  wire popcount23_59hv_core_046;
  wire popcount23_59hv_core_047;
  wire popcount23_59hv_core_048;
  wire popcount23_59hv_core_050;
  wire popcount23_59hv_core_052;
  wire popcount23_59hv_core_053;
  wire popcount23_59hv_core_054;
  wire popcount23_59hv_core_055;
  wire popcount23_59hv_core_057;
  wire popcount23_59hv_core_059;
  wire popcount23_59hv_core_062;
  wire popcount23_59hv_core_063;
  wire popcount23_59hv_core_064;
  wire popcount23_59hv_core_065;
  wire popcount23_59hv_core_066;
  wire popcount23_59hv_core_067;
  wire popcount23_59hv_core_070;
  wire popcount23_59hv_core_071;
  wire popcount23_59hv_core_073;
  wire popcount23_59hv_core_074;
  wire popcount23_59hv_core_076;
  wire popcount23_59hv_core_078;
  wire popcount23_59hv_core_079;
  wire popcount23_59hv_core_080;
  wire popcount23_59hv_core_083;
  wire popcount23_59hv_core_084;
  wire popcount23_59hv_core_085;
  wire popcount23_59hv_core_086;
  wire popcount23_59hv_core_088;
  wire popcount23_59hv_core_089;
  wire popcount23_59hv_core_090;
  wire popcount23_59hv_core_092;
  wire popcount23_59hv_core_093;
  wire popcount23_59hv_core_094_not;
  wire popcount23_59hv_core_095;
  wire popcount23_59hv_core_097;
  wire popcount23_59hv_core_098;
  wire popcount23_59hv_core_099;
  wire popcount23_59hv_core_100;
  wire popcount23_59hv_core_102;
  wire popcount23_59hv_core_103;
  wire popcount23_59hv_core_104;
  wire popcount23_59hv_core_106;
  wire popcount23_59hv_core_107;
  wire popcount23_59hv_core_108;
  wire popcount23_59hv_core_109;
  wire popcount23_59hv_core_110;
  wire popcount23_59hv_core_115;
  wire popcount23_59hv_core_117;
  wire popcount23_59hv_core_120;
  wire popcount23_59hv_core_121;
  wire popcount23_59hv_core_123;
  wire popcount23_59hv_core_124;
  wire popcount23_59hv_core_125;
  wire popcount23_59hv_core_127;
  wire popcount23_59hv_core_128;
  wire popcount23_59hv_core_129;
  wire popcount23_59hv_core_130;
  wire popcount23_59hv_core_131;
  wire popcount23_59hv_core_132;
  wire popcount23_59hv_core_134;
  wire popcount23_59hv_core_136;
  wire popcount23_59hv_core_137;
  wire popcount23_59hv_core_138;
  wire popcount23_59hv_core_143;
  wire popcount23_59hv_core_145;
  wire popcount23_59hv_core_149;
  wire popcount23_59hv_core_150;
  wire popcount23_59hv_core_152;
  wire popcount23_59hv_core_155;
  wire popcount23_59hv_core_157;
  wire popcount23_59hv_core_158;
  wire popcount23_59hv_core_159;
  wire popcount23_59hv_core_161_not;
  wire popcount23_59hv_core_164;
  wire popcount23_59hv_core_165;
  wire popcount23_59hv_core_166;
  wire popcount23_59hv_core_167;

  assign popcount23_59hv_core_026 = input_a[1] | input_a[8];
  assign popcount23_59hv_core_027 = input_a[2] | input_a[15];
  assign popcount23_59hv_core_029 = ~(input_a[6] | input_a[3]);
  assign popcount23_59hv_core_031 = ~(input_a[21] ^ input_a[3]);
  assign popcount23_59hv_core_032 = input_a[18] | input_a[16];
  assign popcount23_59hv_core_035 = input_a[18] ^ input_a[7];
  assign popcount23_59hv_core_036_not = ~input_a[5];
  assign popcount23_59hv_core_039 = ~input_a[11];
  assign popcount23_59hv_core_044 = input_a[11] & input_a[14];
  assign popcount23_59hv_core_046 = ~(input_a[14] & input_a[10]);
  assign popcount23_59hv_core_047 = ~(input_a[12] ^ input_a[7]);
  assign popcount23_59hv_core_048 = input_a[10] & input_a[10];
  assign popcount23_59hv_core_050 = input_a[17] | input_a[1];
  assign popcount23_59hv_core_052 = ~(input_a[17] | input_a[9]);
  assign popcount23_59hv_core_053 = ~input_a[13];
  assign popcount23_59hv_core_054 = ~(input_a[9] | input_a[11]);
  assign popcount23_59hv_core_055 = ~input_a[9];
  assign popcount23_59hv_core_057 = ~(input_a[20] ^ input_a[12]);
  assign popcount23_59hv_core_059 = input_a[0] & input_a[6];
  assign popcount23_59hv_core_062 = ~(input_a[19] | input_a[10]);
  assign popcount23_59hv_core_063 = ~(input_a[6] & input_a[6]);
  assign popcount23_59hv_core_064 = input_a[14] & input_a[2];
  assign popcount23_59hv_core_065 = input_a[11] | input_a[9];
  assign popcount23_59hv_core_066 = ~(input_a[9] | input_a[14]);
  assign popcount23_59hv_core_067 = input_a[11] | input_a[17];
  assign popcount23_59hv_core_070 = ~(input_a[21] & input_a[11]);
  assign popcount23_59hv_core_071 = ~(input_a[9] & input_a[2]);
  assign popcount23_59hv_core_073 = ~(input_a[8] ^ input_a[21]);
  assign popcount23_59hv_core_074 = ~(input_a[18] ^ input_a[22]);
  assign popcount23_59hv_core_076 = ~(input_a[16] ^ input_a[20]);
  assign popcount23_59hv_core_078 = input_a[20] & input_a[13];
  assign popcount23_59hv_core_079 = ~input_a[6];
  assign popcount23_59hv_core_080 = input_a[22] | input_a[11];
  assign popcount23_59hv_core_083 = input_a[15] & input_a[17];
  assign popcount23_59hv_core_084 = ~(input_a[22] | input_a[0]);
  assign popcount23_59hv_core_085 = ~(input_a[9] ^ input_a[9]);
  assign popcount23_59hv_core_086 = input_a[3] | input_a[10];
  assign popcount23_59hv_core_088 = ~(input_a[19] ^ input_a[18]);
  assign popcount23_59hv_core_089 = ~(input_a[21] & input_a[11]);
  assign popcount23_59hv_core_090 = input_a[0] ^ input_a[3];
  assign popcount23_59hv_core_092 = input_a[0] | input_a[2];
  assign popcount23_59hv_core_093 = ~input_a[6];
  assign popcount23_59hv_core_094_not = ~input_a[18];
  assign popcount23_59hv_core_095 = ~(input_a[17] & input_a[20]);
  assign popcount23_59hv_core_097 = ~(input_a[9] | input_a[15]);
  assign popcount23_59hv_core_098 = input_a[4] ^ input_a[8];
  assign popcount23_59hv_core_099 = ~input_a[13];
  assign popcount23_59hv_core_100 = input_a[20] | input_a[4];
  assign popcount23_59hv_core_102 = input_a[20] | input_a[16];
  assign popcount23_59hv_core_103 = input_a[14] ^ input_a[2];
  assign popcount23_59hv_core_104 = input_a[2] & input_a[6];
  assign popcount23_59hv_core_106 = input_a[15] | input_a[20];
  assign popcount23_59hv_core_107 = ~(input_a[18] ^ input_a[8]);
  assign popcount23_59hv_core_108 = ~(input_a[13] | input_a[11]);
  assign popcount23_59hv_core_109 = ~(input_a[4] ^ input_a[6]);
  assign popcount23_59hv_core_110 = input_a[19] & input_a[20];
  assign popcount23_59hv_core_115 = input_a[16] ^ input_a[22];
  assign popcount23_59hv_core_117 = input_a[6] & input_a[18];
  assign popcount23_59hv_core_120 = ~(input_a[6] | input_a[6]);
  assign popcount23_59hv_core_121 = input_a[9] ^ input_a[15];
  assign popcount23_59hv_core_123 = input_a[20] | input_a[2];
  assign popcount23_59hv_core_124 = ~(input_a[3] | input_a[2]);
  assign popcount23_59hv_core_125 = ~(input_a[9] | input_a[20]);
  assign popcount23_59hv_core_127 = ~input_a[7];
  assign popcount23_59hv_core_128 = input_a[18] | input_a[19];
  assign popcount23_59hv_core_129 = input_a[0] & input_a[9];
  assign popcount23_59hv_core_130 = input_a[1] | input_a[10];
  assign popcount23_59hv_core_131 = input_a[2] & input_a[1];
  assign popcount23_59hv_core_132 = input_a[1] ^ input_a[13];
  assign popcount23_59hv_core_134 = input_a[21] ^ input_a[20];
  assign popcount23_59hv_core_136 = ~input_a[15];
  assign popcount23_59hv_core_137 = input_a[2] & input_a[14];
  assign popcount23_59hv_core_138 = ~(input_a[10] ^ input_a[12]);
  assign popcount23_59hv_core_143 = ~(input_a[22] & input_a[17]);
  assign popcount23_59hv_core_145 = input_a[17] & input_a[20];
  assign popcount23_59hv_core_149 = ~input_a[8];
  assign popcount23_59hv_core_150 = input_a[18] ^ input_a[1];
  assign popcount23_59hv_core_152 = ~(input_a[21] | input_a[4]);
  assign popcount23_59hv_core_155 = ~(input_a[20] & input_a[16]);
  assign popcount23_59hv_core_157 = ~input_a[22];
  assign popcount23_59hv_core_158 = input_a[18] ^ input_a[12];
  assign popcount23_59hv_core_159 = input_a[17] | input_a[0];
  assign popcount23_59hv_core_161_not = ~input_a[12];
  assign popcount23_59hv_core_164 = ~input_a[4];
  assign popcount23_59hv_core_165 = ~(input_a[20] | input_a[14]);
  assign popcount23_59hv_core_166 = ~(input_a[18] ^ input_a[8]);
  assign popcount23_59hv_core_167 = ~(input_a[11] | input_a[0]);

  assign popcount23_59hv_out[0] = input_a[15];
  assign popcount23_59hv_out[1] = input_a[10];
  assign popcount23_59hv_out[2] = input_a[10];
  assign popcount23_59hv_out[3] = 1'b0;
  assign popcount23_59hv_out[4] = input_a[9];
endmodule