// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.2392
// WCE=16.0
// EP=0.86005%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount32_ckmq(input [31:0] input_a, output [5:0] popcount32_ckmq_out);
  wire popcount32_ckmq_core_034;
  wire popcount32_ckmq_core_035;
  wire popcount32_ckmq_core_036;
  wire popcount32_ckmq_core_038;
  wire popcount32_ckmq_core_039;
  wire popcount32_ckmq_core_040_not;
  wire popcount32_ckmq_core_042;
  wire popcount32_ckmq_core_043;
  wire popcount32_ckmq_core_044;
  wire popcount32_ckmq_core_045;
  wire popcount32_ckmq_core_046;
  wire popcount32_ckmq_core_047;
  wire popcount32_ckmq_core_048;
  wire popcount32_ckmq_core_049_not;
  wire popcount32_ckmq_core_051;
  wire popcount32_ckmq_core_053;
  wire popcount32_ckmq_core_054;
  wire popcount32_ckmq_core_055;
  wire popcount32_ckmq_core_056;
  wire popcount32_ckmq_core_057_not;
  wire popcount32_ckmq_core_058;
  wire popcount32_ckmq_core_060;
  wire popcount32_ckmq_core_061;
  wire popcount32_ckmq_core_062;
  wire popcount32_ckmq_core_063;
  wire popcount32_ckmq_core_064;
  wire popcount32_ckmq_core_066;
  wire popcount32_ckmq_core_068;
  wire popcount32_ckmq_core_069;
  wire popcount32_ckmq_core_071;
  wire popcount32_ckmq_core_073;
  wire popcount32_ckmq_core_074;
  wire popcount32_ckmq_core_075;
  wire popcount32_ckmq_core_076;
  wire popcount32_ckmq_core_078;
  wire popcount32_ckmq_core_080;
  wire popcount32_ckmq_core_081;
  wire popcount32_ckmq_core_082;
  wire popcount32_ckmq_core_083;
  wire popcount32_ckmq_core_084;
  wire popcount32_ckmq_core_085_not;
  wire popcount32_ckmq_core_087;
  wire popcount32_ckmq_core_088;
  wire popcount32_ckmq_core_089;
  wire popcount32_ckmq_core_090;
  wire popcount32_ckmq_core_091;
  wire popcount32_ckmq_core_092;
  wire popcount32_ckmq_core_093;
  wire popcount32_ckmq_core_094;
  wire popcount32_ckmq_core_096;
  wire popcount32_ckmq_core_097;
  wire popcount32_ckmq_core_098;
  wire popcount32_ckmq_core_100;
  wire popcount32_ckmq_core_101;
  wire popcount32_ckmq_core_102;
  wire popcount32_ckmq_core_103;
  wire popcount32_ckmq_core_104;
  wire popcount32_ckmq_core_105_not;
  wire popcount32_ckmq_core_108;
  wire popcount32_ckmq_core_110;
  wire popcount32_ckmq_core_112_not;
  wire popcount32_ckmq_core_116;
  wire popcount32_ckmq_core_117;
  wire popcount32_ckmq_core_118;
  wire popcount32_ckmq_core_120;
  wire popcount32_ckmq_core_121;
  wire popcount32_ckmq_core_124;
  wire popcount32_ckmq_core_127;
  wire popcount32_ckmq_core_129;
  wire popcount32_ckmq_core_130;
  wire popcount32_ckmq_core_131;
  wire popcount32_ckmq_core_132;
  wire popcount32_ckmq_core_133;
  wire popcount32_ckmq_core_134;
  wire popcount32_ckmq_core_135;
  wire popcount32_ckmq_core_137;
  wire popcount32_ckmq_core_138;
  wire popcount32_ckmq_core_139;
  wire popcount32_ckmq_core_141;
  wire popcount32_ckmq_core_142;
  wire popcount32_ckmq_core_144;
  wire popcount32_ckmq_core_145;
  wire popcount32_ckmq_core_146;
  wire popcount32_ckmq_core_148;
  wire popcount32_ckmq_core_149;
  wire popcount32_ckmq_core_150;
  wire popcount32_ckmq_core_151;
  wire popcount32_ckmq_core_152;
  wire popcount32_ckmq_core_155;
  wire popcount32_ckmq_core_156;
  wire popcount32_ckmq_core_157;
  wire popcount32_ckmq_core_158;
  wire popcount32_ckmq_core_160;
  wire popcount32_ckmq_core_161;
  wire popcount32_ckmq_core_162;
  wire popcount32_ckmq_core_165;
  wire popcount32_ckmq_core_168;
  wire popcount32_ckmq_core_169;
  wire popcount32_ckmq_core_173;
  wire popcount32_ckmq_core_174;
  wire popcount32_ckmq_core_176;
  wire popcount32_ckmq_core_177;
  wire popcount32_ckmq_core_178;
  wire popcount32_ckmq_core_179;
  wire popcount32_ckmq_core_180;
  wire popcount32_ckmq_core_181;
  wire popcount32_ckmq_core_182;
  wire popcount32_ckmq_core_185_not;
  wire popcount32_ckmq_core_189;
  wire popcount32_ckmq_core_190;
  wire popcount32_ckmq_core_191;
  wire popcount32_ckmq_core_192;
  wire popcount32_ckmq_core_193;
  wire popcount32_ckmq_core_195;
  wire popcount32_ckmq_core_196;
  wire popcount32_ckmq_core_197;
  wire popcount32_ckmq_core_198;
  wire popcount32_ckmq_core_199;
  wire popcount32_ckmq_core_203;
  wire popcount32_ckmq_core_205;
  wire popcount32_ckmq_core_206;
  wire popcount32_ckmq_core_207;
  wire popcount32_ckmq_core_209;
  wire popcount32_ckmq_core_210;
  wire popcount32_ckmq_core_211;
  wire popcount32_ckmq_core_213;
  wire popcount32_ckmq_core_214;
  wire popcount32_ckmq_core_215;
  wire popcount32_ckmq_core_219;
  wire popcount32_ckmq_core_220;
  wire popcount32_ckmq_core_223_not;
  wire popcount32_ckmq_core_224;

  assign popcount32_ckmq_core_034 = input_a[6] & input_a[19];
  assign popcount32_ckmq_core_035 = input_a[29] ^ input_a[3];
  assign popcount32_ckmq_core_036 = ~input_a[29];
  assign popcount32_ckmq_core_038 = input_a[9] & input_a[24];
  assign popcount32_ckmq_core_039 = ~input_a[24];
  assign popcount32_ckmq_core_040_not = ~input_a[8];
  assign popcount32_ckmq_core_042 = ~(input_a[9] ^ input_a[12]);
  assign popcount32_ckmq_core_043 = ~input_a[3];
  assign popcount32_ckmq_core_044 = ~(input_a[18] ^ input_a[30]);
  assign popcount32_ckmq_core_045 = input_a[25] ^ input_a[16];
  assign popcount32_ckmq_core_046 = input_a[2] ^ input_a[9];
  assign popcount32_ckmq_core_047 = ~(input_a[29] & input_a[7]);
  assign popcount32_ckmq_core_048 = ~(input_a[27] & input_a[13]);
  assign popcount32_ckmq_core_049_not = ~input_a[9];
  assign popcount32_ckmq_core_051 = ~input_a[0];
  assign popcount32_ckmq_core_053 = ~(input_a[15] ^ input_a[0]);
  assign popcount32_ckmq_core_054 = input_a[9] | input_a[16];
  assign popcount32_ckmq_core_055 = ~(input_a[9] ^ input_a[12]);
  assign popcount32_ckmq_core_056 = ~(input_a[22] | input_a[8]);
  assign popcount32_ckmq_core_057_not = ~input_a[5];
  assign popcount32_ckmq_core_058 = ~(input_a[16] ^ input_a[23]);
  assign popcount32_ckmq_core_060 = ~input_a[29];
  assign popcount32_ckmq_core_061 = input_a[23] | input_a[16];
  assign popcount32_ckmq_core_062 = ~(input_a[7] & input_a[4]);
  assign popcount32_ckmq_core_063 = ~input_a[6];
  assign popcount32_ckmq_core_064 = ~input_a[25];
  assign popcount32_ckmq_core_066 = input_a[26] & input_a[17];
  assign popcount32_ckmq_core_068 = ~(input_a[2] & input_a[9]);
  assign popcount32_ckmq_core_069 = ~(input_a[18] ^ input_a[31]);
  assign popcount32_ckmq_core_071 = input_a[24] | input_a[2];
  assign popcount32_ckmq_core_073 = input_a[20] ^ input_a[19];
  assign popcount32_ckmq_core_074 = ~input_a[6];
  assign popcount32_ckmq_core_075 = ~(input_a[5] & input_a[10]);
  assign popcount32_ckmq_core_076 = input_a[0] | input_a[7];
  assign popcount32_ckmq_core_078 = ~input_a[13];
  assign popcount32_ckmq_core_080 = input_a[1] | input_a[5];
  assign popcount32_ckmq_core_081 = ~(input_a[19] & input_a[9]);
  assign popcount32_ckmq_core_082 = ~(input_a[21] & input_a[27]);
  assign popcount32_ckmq_core_083 = input_a[7] & input_a[10];
  assign popcount32_ckmq_core_084 = ~input_a[24];
  assign popcount32_ckmq_core_085_not = ~input_a[16];
  assign popcount32_ckmq_core_087 = input_a[28] ^ input_a[20];
  assign popcount32_ckmq_core_088 = ~(input_a[10] ^ input_a[4]);
  assign popcount32_ckmq_core_089 = ~(input_a[4] | input_a[0]);
  assign popcount32_ckmq_core_090 = ~(input_a[23] ^ input_a[15]);
  assign popcount32_ckmq_core_091 = ~(input_a[29] ^ input_a[28]);
  assign popcount32_ckmq_core_092 = ~(input_a[5] & input_a[22]);
  assign popcount32_ckmq_core_093 = ~(input_a[15] ^ input_a[0]);
  assign popcount32_ckmq_core_094 = input_a[22] | input_a[6];
  assign popcount32_ckmq_core_096 = ~(input_a[21] & input_a[28]);
  assign popcount32_ckmq_core_097 = ~(input_a[1] & input_a[1]);
  assign popcount32_ckmq_core_098 = ~(input_a[5] | input_a[13]);
  assign popcount32_ckmq_core_100 = input_a[2] ^ input_a[16];
  assign popcount32_ckmq_core_101 = ~(input_a[14] ^ input_a[26]);
  assign popcount32_ckmq_core_102 = ~(input_a[12] & input_a[11]);
  assign popcount32_ckmq_core_103 = ~(input_a[29] & input_a[1]);
  assign popcount32_ckmq_core_104 = ~(input_a[30] ^ input_a[22]);
  assign popcount32_ckmq_core_105_not = ~input_a[5];
  assign popcount32_ckmq_core_108 = input_a[25] ^ input_a[24];
  assign popcount32_ckmq_core_110 = ~(input_a[27] ^ input_a[14]);
  assign popcount32_ckmq_core_112_not = ~input_a[30];
  assign popcount32_ckmq_core_116 = ~(input_a[9] ^ input_a[26]);
  assign popcount32_ckmq_core_117 = ~input_a[30];
  assign popcount32_ckmq_core_118 = ~(input_a[14] & input_a[10]);
  assign popcount32_ckmq_core_120 = ~(input_a[30] & input_a[3]);
  assign popcount32_ckmq_core_121 = ~(input_a[18] | input_a[8]);
  assign popcount32_ckmq_core_124 = ~(input_a[1] ^ input_a[12]);
  assign popcount32_ckmq_core_127 = ~(input_a[5] | input_a[10]);
  assign popcount32_ckmq_core_129 = ~(input_a[10] & input_a[1]);
  assign popcount32_ckmq_core_130 = input_a[9] | input_a[25];
  assign popcount32_ckmq_core_131 = ~(input_a[4] & input_a[8]);
  assign popcount32_ckmq_core_132 = input_a[10] ^ input_a[27];
  assign popcount32_ckmq_core_133 = ~(input_a[31] ^ input_a[16]);
  assign popcount32_ckmq_core_134 = input_a[14] & input_a[29];
  assign popcount32_ckmq_core_135 = ~(input_a[0] ^ input_a[2]);
  assign popcount32_ckmq_core_137 = ~(input_a[10] | input_a[23]);
  assign popcount32_ckmq_core_138 = ~(input_a[29] | input_a[14]);
  assign popcount32_ckmq_core_139 = ~(input_a[0] ^ input_a[30]);
  assign popcount32_ckmq_core_141 = input_a[24] ^ input_a[25];
  assign popcount32_ckmq_core_142 = input_a[11] & input_a[2];
  assign popcount32_ckmq_core_144 = input_a[29] | input_a[8];
  assign popcount32_ckmq_core_145 = ~(input_a[25] | input_a[20]);
  assign popcount32_ckmq_core_146 = ~(input_a[12] | input_a[16]);
  assign popcount32_ckmq_core_148 = input_a[14] & input_a[5];
  assign popcount32_ckmq_core_149 = ~(input_a[14] | input_a[1]);
  assign popcount32_ckmq_core_150 = input_a[1] ^ input_a[24];
  assign popcount32_ckmq_core_151 = ~(input_a[18] | input_a[2]);
  assign popcount32_ckmq_core_152 = ~(input_a[7] & input_a[15]);
  assign popcount32_ckmq_core_155 = ~(input_a[26] | input_a[18]);
  assign popcount32_ckmq_core_156 = input_a[0] ^ input_a[16];
  assign popcount32_ckmq_core_157 = input_a[26] ^ input_a[13];
  assign popcount32_ckmq_core_158 = ~(input_a[30] & input_a[28]);
  assign popcount32_ckmq_core_160 = input_a[27] ^ input_a[27];
  assign popcount32_ckmq_core_161 = input_a[11] ^ input_a[22];
  assign popcount32_ckmq_core_162 = input_a[27] ^ input_a[20];
  assign popcount32_ckmq_core_165 = ~(input_a[25] & input_a[26]);
  assign popcount32_ckmq_core_168 = ~(input_a[10] | input_a[13]);
  assign popcount32_ckmq_core_169 = input_a[12] & input_a[16];
  assign popcount32_ckmq_core_173 = ~(input_a[24] ^ input_a[15]);
  assign popcount32_ckmq_core_174 = input_a[12] ^ input_a[3];
  assign popcount32_ckmq_core_176 = ~(input_a[14] ^ input_a[0]);
  assign popcount32_ckmq_core_177 = ~(input_a[27] & input_a[1]);
  assign popcount32_ckmq_core_178 = input_a[31] ^ input_a[30];
  assign popcount32_ckmq_core_179 = input_a[18] ^ input_a[30];
  assign popcount32_ckmq_core_180 = input_a[14] ^ input_a[10];
  assign popcount32_ckmq_core_181 = ~(input_a[24] | input_a[22]);
  assign popcount32_ckmq_core_182 = input_a[19] | input_a[6];
  assign popcount32_ckmq_core_185_not = ~input_a[12];
  assign popcount32_ckmq_core_189 = input_a[14] & input_a[4];
  assign popcount32_ckmq_core_190 = ~input_a[12];
  assign popcount32_ckmq_core_191 = input_a[26] & input_a[16];
  assign popcount32_ckmq_core_192 = input_a[29] | input_a[6];
  assign popcount32_ckmq_core_193 = input_a[31] & input_a[26];
  assign popcount32_ckmq_core_195 = ~(input_a[14] ^ input_a[6]);
  assign popcount32_ckmq_core_196 = input_a[24] | input_a[22];
  assign popcount32_ckmq_core_197 = ~(input_a[14] ^ input_a[7]);
  assign popcount32_ckmq_core_198 = ~(input_a[13] ^ input_a[2]);
  assign popcount32_ckmq_core_199 = input_a[14] | input_a[13];
  assign popcount32_ckmq_core_203 = ~(input_a[10] & input_a[14]);
  assign popcount32_ckmq_core_205 = ~(input_a[1] & input_a[16]);
  assign popcount32_ckmq_core_206 = ~(input_a[17] ^ input_a[3]);
  assign popcount32_ckmq_core_207 = ~(input_a[16] | input_a[21]);
  assign popcount32_ckmq_core_209 = ~(input_a[11] & input_a[24]);
  assign popcount32_ckmq_core_210 = ~(input_a[23] | input_a[30]);
  assign popcount32_ckmq_core_211 = ~input_a[10];
  assign popcount32_ckmq_core_213 = input_a[11] & input_a[21];
  assign popcount32_ckmq_core_214 = ~input_a[25];
  assign popcount32_ckmq_core_215 = ~(input_a[0] ^ input_a[13]);
  assign popcount32_ckmq_core_219 = input_a[24] & input_a[6];
  assign popcount32_ckmq_core_220 = input_a[25] | input_a[9];
  assign popcount32_ckmq_core_223_not = ~input_a[28];
  assign popcount32_ckmq_core_224 = ~(input_a[27] ^ input_a[2]);

  assign popcount32_ckmq_out[0] = input_a[0];
  assign popcount32_ckmq_out[1] = popcount32_ckmq_core_211;
  assign popcount32_ckmq_out[2] = popcount32_ckmq_core_211;
  assign popcount32_ckmq_out[3] = popcount32_ckmq_core_211;
  assign popcount32_ckmq_out[4] = input_a[10];
  assign popcount32_ckmq_out[5] = 1'b0;
endmodule