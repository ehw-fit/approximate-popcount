// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.04597
// WCE=18.0
// EP=0.903956%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_j87r(input [31:0] input_a, output [5:0] popcount32_j87r_out);
  wire popcount32_j87r_core_034;
  wire popcount32_j87r_core_035;
  wire popcount32_j87r_core_036;
  wire popcount32_j87r_core_038;
  wire popcount32_j87r_core_039;
  wire popcount32_j87r_core_042;
  wire popcount32_j87r_core_044;
  wire popcount32_j87r_core_047;
  wire popcount32_j87r_core_050;
  wire popcount32_j87r_core_051;
  wire popcount32_j87r_core_052;
  wire popcount32_j87r_core_053;
  wire popcount32_j87r_core_055;
  wire popcount32_j87r_core_056;
  wire popcount32_j87r_core_057;
  wire popcount32_j87r_core_058;
  wire popcount32_j87r_core_060;
  wire popcount32_j87r_core_061;
  wire popcount32_j87r_core_062;
  wire popcount32_j87r_core_063;
  wire popcount32_j87r_core_064;
  wire popcount32_j87r_core_065;
  wire popcount32_j87r_core_066;
  wire popcount32_j87r_core_068;
  wire popcount32_j87r_core_069;
  wire popcount32_j87r_core_071_not;
  wire popcount32_j87r_core_072;
  wire popcount32_j87r_core_074;
  wire popcount32_j87r_core_075;
  wire popcount32_j87r_core_076;
  wire popcount32_j87r_core_077;
  wire popcount32_j87r_core_078;
  wire popcount32_j87r_core_079;
  wire popcount32_j87r_core_081;
  wire popcount32_j87r_core_082;
  wire popcount32_j87r_core_083;
  wire popcount32_j87r_core_086;
  wire popcount32_j87r_core_087;
  wire popcount32_j87r_core_088;
  wire popcount32_j87r_core_089;
  wire popcount32_j87r_core_090;
  wire popcount32_j87r_core_092;
  wire popcount32_j87r_core_096;
  wire popcount32_j87r_core_097;
  wire popcount32_j87r_core_099;
  wire popcount32_j87r_core_100;
  wire popcount32_j87r_core_101;
  wire popcount32_j87r_core_103;
  wire popcount32_j87r_core_104;
  wire popcount32_j87r_core_105;
  wire popcount32_j87r_core_106;
  wire popcount32_j87r_core_107;
  wire popcount32_j87r_core_108;
  wire popcount32_j87r_core_109;
  wire popcount32_j87r_core_116;
  wire popcount32_j87r_core_117;
  wire popcount32_j87r_core_118;
  wire popcount32_j87r_core_120;
  wire popcount32_j87r_core_121;
  wire popcount32_j87r_core_122;
  wire popcount32_j87r_core_123;
  wire popcount32_j87r_core_125;
  wire popcount32_j87r_core_126;
  wire popcount32_j87r_core_127;
  wire popcount32_j87r_core_128;
  wire popcount32_j87r_core_129;
  wire popcount32_j87r_core_130;
  wire popcount32_j87r_core_132;
  wire popcount32_j87r_core_133;
  wire popcount32_j87r_core_135;
  wire popcount32_j87r_core_137;
  wire popcount32_j87r_core_140;
  wire popcount32_j87r_core_142;
  wire popcount32_j87r_core_144;
  wire popcount32_j87r_core_145;
  wire popcount32_j87r_core_146;
  wire popcount32_j87r_core_147;
  wire popcount32_j87r_core_149;
  wire popcount32_j87r_core_151;
  wire popcount32_j87r_core_152;
  wire popcount32_j87r_core_154;
  wire popcount32_j87r_core_155;
  wire popcount32_j87r_core_156_not;
  wire popcount32_j87r_core_157;
  wire popcount32_j87r_core_158;
  wire popcount32_j87r_core_159;
  wire popcount32_j87r_core_161;
  wire popcount32_j87r_core_163;
  wire popcount32_j87r_core_166;
  wire popcount32_j87r_core_169;
  wire popcount32_j87r_core_170_not;
  wire popcount32_j87r_core_171;
  wire popcount32_j87r_core_172;
  wire popcount32_j87r_core_173;
  wire popcount32_j87r_core_174;
  wire popcount32_j87r_core_175;
  wire popcount32_j87r_core_178;
  wire popcount32_j87r_core_180;
  wire popcount32_j87r_core_181;
  wire popcount32_j87r_core_182;
  wire popcount32_j87r_core_183;
  wire popcount32_j87r_core_185;
  wire popcount32_j87r_core_187;
  wire popcount32_j87r_core_192;
  wire popcount32_j87r_core_195;
  wire popcount32_j87r_core_196;
  wire popcount32_j87r_core_197;
  wire popcount32_j87r_core_199;
  wire popcount32_j87r_core_201;
  wire popcount32_j87r_core_203;
  wire popcount32_j87r_core_205;
  wire popcount32_j87r_core_206;
  wire popcount32_j87r_core_207;
  wire popcount32_j87r_core_208;
  wire popcount32_j87r_core_209;
  wire popcount32_j87r_core_210;
  wire popcount32_j87r_core_215;
  wire popcount32_j87r_core_217;
  wire popcount32_j87r_core_219;
  wire popcount32_j87r_core_223_not;
  wire popcount32_j87r_core_224;
  wire popcount32_j87r_core_225;

  assign popcount32_j87r_core_034 = ~(input_a[12] ^ input_a[27]);
  assign popcount32_j87r_core_035 = ~(input_a[20] ^ input_a[31]);
  assign popcount32_j87r_core_036 = input_a[7] | input_a[21];
  assign popcount32_j87r_core_038 = ~(input_a[13] ^ input_a[10]);
  assign popcount32_j87r_core_039 = ~(input_a[10] | input_a[21]);
  assign popcount32_j87r_core_042 = ~input_a[1];
  assign popcount32_j87r_core_044 = ~input_a[3];
  assign popcount32_j87r_core_047 = input_a[7] ^ input_a[13];
  assign popcount32_j87r_core_050 = input_a[14] ^ input_a[24];
  assign popcount32_j87r_core_051 = input_a[14] | input_a[31];
  assign popcount32_j87r_core_052 = ~(input_a[29] & input_a[6]);
  assign popcount32_j87r_core_053 = input_a[25] & input_a[25];
  assign popcount32_j87r_core_055 = ~(input_a[31] & input_a[11]);
  assign popcount32_j87r_core_056 = ~(input_a[18] ^ input_a[30]);
  assign popcount32_j87r_core_057 = ~(input_a[18] | input_a[25]);
  assign popcount32_j87r_core_058 = ~input_a[15];
  assign popcount32_j87r_core_060 = ~(input_a[29] & input_a[22]);
  assign popcount32_j87r_core_061 = ~(input_a[7] | input_a[25]);
  assign popcount32_j87r_core_062 = input_a[12] ^ input_a[13];
  assign popcount32_j87r_core_063 = ~(input_a[28] & input_a[16]);
  assign popcount32_j87r_core_064 = ~(input_a[18] & input_a[11]);
  assign popcount32_j87r_core_065 = input_a[16] & input_a[10];
  assign popcount32_j87r_core_066 = input_a[19] | input_a[17];
  assign popcount32_j87r_core_068 = input_a[24] | input_a[7];
  assign popcount32_j87r_core_069 = input_a[16] | input_a[12];
  assign popcount32_j87r_core_071_not = ~input_a[27];
  assign popcount32_j87r_core_072 = ~(input_a[31] | input_a[28]);
  assign popcount32_j87r_core_074 = input_a[30] ^ input_a[1];
  assign popcount32_j87r_core_075 = input_a[13] | input_a[7];
  assign popcount32_j87r_core_076 = input_a[26] & input_a[13];
  assign popcount32_j87r_core_077 = input_a[1] | input_a[3];
  assign popcount32_j87r_core_078 = ~input_a[0];
  assign popcount32_j87r_core_079 = ~(input_a[27] & input_a[14]);
  assign popcount32_j87r_core_081 = ~(input_a[12] | input_a[24]);
  assign popcount32_j87r_core_082 = input_a[17] ^ input_a[27];
  assign popcount32_j87r_core_083 = input_a[18] | input_a[12];
  assign popcount32_j87r_core_086 = input_a[8] | input_a[2];
  assign popcount32_j87r_core_087 = input_a[5] & input_a[19];
  assign popcount32_j87r_core_088 = input_a[24] ^ input_a[16];
  assign popcount32_j87r_core_089 = ~input_a[7];
  assign popcount32_j87r_core_090 = ~input_a[13];
  assign popcount32_j87r_core_092 = ~(input_a[12] & input_a[26]);
  assign popcount32_j87r_core_096 = input_a[6] | input_a[21];
  assign popcount32_j87r_core_097 = ~input_a[6];
  assign popcount32_j87r_core_099 = input_a[17] | input_a[15];
  assign popcount32_j87r_core_100 = ~(input_a[20] | input_a[2]);
  assign popcount32_j87r_core_101 = input_a[26] & input_a[2];
  assign popcount32_j87r_core_103 = input_a[26] ^ input_a[19];
  assign popcount32_j87r_core_104 = ~(input_a[28] | input_a[23]);
  assign popcount32_j87r_core_105 = ~input_a[31];
  assign popcount32_j87r_core_106 = input_a[24] ^ input_a[21];
  assign popcount32_j87r_core_107 = input_a[0] ^ input_a[26];
  assign popcount32_j87r_core_108 = ~(input_a[1] ^ input_a[0]);
  assign popcount32_j87r_core_109 = input_a[24] | input_a[14];
  assign popcount32_j87r_core_116 = ~(input_a[9] | input_a[0]);
  assign popcount32_j87r_core_117 = input_a[21] & input_a[2];
  assign popcount32_j87r_core_118 = input_a[30] ^ input_a[10];
  assign popcount32_j87r_core_120 = ~(input_a[23] ^ input_a[1]);
  assign popcount32_j87r_core_121 = input_a[26] | input_a[5];
  assign popcount32_j87r_core_122 = ~(input_a[29] ^ input_a[4]);
  assign popcount32_j87r_core_123 = ~input_a[28];
  assign popcount32_j87r_core_125 = input_a[8] ^ input_a[2];
  assign popcount32_j87r_core_126 = ~(input_a[14] & input_a[4]);
  assign popcount32_j87r_core_127 = ~(input_a[2] & input_a[10]);
  assign popcount32_j87r_core_128 = ~(input_a[11] | input_a[21]);
  assign popcount32_j87r_core_129 = ~input_a[26];
  assign popcount32_j87r_core_130 = input_a[29] & input_a[11];
  assign popcount32_j87r_core_132 = input_a[18] & input_a[24];
  assign popcount32_j87r_core_133 = ~(input_a[12] ^ input_a[7]);
  assign popcount32_j87r_core_135 = ~(input_a[24] | input_a[15]);
  assign popcount32_j87r_core_137 = ~input_a[31];
  assign popcount32_j87r_core_140 = ~input_a[12];
  assign popcount32_j87r_core_142 = input_a[23] | input_a[31];
  assign popcount32_j87r_core_144 = input_a[13] & input_a[25];
  assign popcount32_j87r_core_145 = input_a[29] & input_a[10];
  assign popcount32_j87r_core_146 = input_a[17] | input_a[0];
  assign popcount32_j87r_core_147 = input_a[3] | input_a[22];
  assign popcount32_j87r_core_149 = input_a[14] | input_a[23];
  assign popcount32_j87r_core_151 = ~input_a[22];
  assign popcount32_j87r_core_152 = input_a[8] | input_a[14];
  assign popcount32_j87r_core_154 = ~(input_a[28] | input_a[12]);
  assign popcount32_j87r_core_155 = input_a[14] & input_a[10];
  assign popcount32_j87r_core_156_not = ~input_a[9];
  assign popcount32_j87r_core_157 = ~input_a[4];
  assign popcount32_j87r_core_158 = ~(input_a[29] ^ input_a[22]);
  assign popcount32_j87r_core_159 = ~(input_a[9] ^ input_a[19]);
  assign popcount32_j87r_core_161 = ~(input_a[18] & input_a[25]);
  assign popcount32_j87r_core_163 = ~(input_a[13] & input_a[24]);
  assign popcount32_j87r_core_166 = ~(input_a[8] & input_a[21]);
  assign popcount32_j87r_core_169 = input_a[31] ^ input_a[13];
  assign popcount32_j87r_core_170_not = ~input_a[3];
  assign popcount32_j87r_core_171 = input_a[8] & input_a[0];
  assign popcount32_j87r_core_172 = input_a[26] & input_a[27];
  assign popcount32_j87r_core_173 = input_a[18] ^ input_a[19];
  assign popcount32_j87r_core_174 = ~input_a[30];
  assign popcount32_j87r_core_175 = input_a[4] | input_a[7];
  assign popcount32_j87r_core_178 = ~(input_a[3] | input_a[22]);
  assign popcount32_j87r_core_180 = ~(input_a[5] | input_a[23]);
  assign popcount32_j87r_core_181 = input_a[27] ^ input_a[13];
  assign popcount32_j87r_core_182 = ~(input_a[14] | input_a[12]);
  assign popcount32_j87r_core_183 = ~input_a[14];
  assign popcount32_j87r_core_185 = input_a[26] | input_a[14];
  assign popcount32_j87r_core_187 = input_a[26] | input_a[27];
  assign popcount32_j87r_core_192 = ~input_a[16];
  assign popcount32_j87r_core_195 = ~(input_a[22] ^ input_a[27]);
  assign popcount32_j87r_core_196 = ~input_a[27];
  assign popcount32_j87r_core_197 = input_a[10] ^ input_a[28];
  assign popcount32_j87r_core_199 = input_a[30] ^ input_a[4];
  assign popcount32_j87r_core_201 = input_a[9] | input_a[19];
  assign popcount32_j87r_core_203 = input_a[29] ^ input_a[11];
  assign popcount32_j87r_core_205 = ~(input_a[20] & input_a[11]);
  assign popcount32_j87r_core_206 = ~(input_a[10] | input_a[7]);
  assign popcount32_j87r_core_207 = ~input_a[6];
  assign popcount32_j87r_core_208 = ~(input_a[1] ^ input_a[26]);
  assign popcount32_j87r_core_209 = ~(input_a[22] & input_a[11]);
  assign popcount32_j87r_core_210 = ~(input_a[10] | input_a[4]);
  assign popcount32_j87r_core_215 = input_a[11] & input_a[25];
  assign popcount32_j87r_core_217 = ~input_a[9];
  assign popcount32_j87r_core_219 = ~(input_a[6] ^ input_a[5]);
  assign popcount32_j87r_core_223_not = ~input_a[1];
  assign popcount32_j87r_core_224 = input_a[5] | input_a[27];
  assign popcount32_j87r_core_225 = ~(input_a[7] & input_a[2]);

  assign popcount32_j87r_out[0] = input_a[13];
  assign popcount32_j87r_out[1] = input_a[14];
  assign popcount32_j87r_out[2] = 1'b1;
  assign popcount32_j87r_out[3] = 1'b1;
  assign popcount32_j87r_out[4] = 1'b0;
  assign popcount32_j87r_out[5] = 1'b0;
endmodule