// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.58979
// WCE=34.0
// EP=0.910004%
// Printed PDK parameters:
//  Area=53491792.0
//  Delay=65343904.0
//  Power=2957500.0

module popcount36_2ba4(input [35:0] input_a, output [5:0] popcount36_2ba4_out);
  wire popcount36_2ba4_core_038;
  wire popcount36_2ba4_core_039;
  wire popcount36_2ba4_core_040;
  wire popcount36_2ba4_core_041;
  wire popcount36_2ba4_core_042;
  wire popcount36_2ba4_core_043;
  wire popcount36_2ba4_core_044;
  wire popcount36_2ba4_core_046;
  wire popcount36_2ba4_core_048;
  wire popcount36_2ba4_core_050;
  wire popcount36_2ba4_core_051;
  wire popcount36_2ba4_core_052;
  wire popcount36_2ba4_core_053;
  wire popcount36_2ba4_core_054;
  wire popcount36_2ba4_core_056;
  wire popcount36_2ba4_core_057;
  wire popcount36_2ba4_core_058;
  wire popcount36_2ba4_core_061;
  wire popcount36_2ba4_core_062;
  wire popcount36_2ba4_core_066;
  wire popcount36_2ba4_core_067;
  wire popcount36_2ba4_core_068;
  wire popcount36_2ba4_core_069;
  wire popcount36_2ba4_core_070;
  wire popcount36_2ba4_core_071;
  wire popcount36_2ba4_core_072;
  wire popcount36_2ba4_core_081;
  wire popcount36_2ba4_core_082;
  wire popcount36_2ba4_core_083;
  wire popcount36_2ba4_core_084;
  wire popcount36_2ba4_core_086;
  wire popcount36_2ba4_core_087;
  wire popcount36_2ba4_core_088;
  wire popcount36_2ba4_core_089;
  wire popcount36_2ba4_core_090;
  wire popcount36_2ba4_core_091;
  wire popcount36_2ba4_core_092;
  wire popcount36_2ba4_core_093;
  wire popcount36_2ba4_core_096;
  wire popcount36_2ba4_core_099_not;
  wire popcount36_2ba4_core_101;
  wire popcount36_2ba4_core_102;
  wire popcount36_2ba4_core_103;
  wire popcount36_2ba4_core_104;
  wire popcount36_2ba4_core_105;
  wire popcount36_2ba4_core_106;
  wire popcount36_2ba4_core_110;
  wire popcount36_2ba4_core_111;
  wire popcount36_2ba4_core_115;
  wire popcount36_2ba4_core_116;
  wire popcount36_2ba4_core_117;
  wire popcount36_2ba4_core_118;
  wire popcount36_2ba4_core_119;
  wire popcount36_2ba4_core_124;
  wire popcount36_2ba4_core_125;
  wire popcount36_2ba4_core_128;
  wire popcount36_2ba4_core_129;
  wire popcount36_2ba4_core_131;
  wire popcount36_2ba4_core_132;
  wire popcount36_2ba4_core_136;
  wire popcount36_2ba4_core_137;
  wire popcount36_2ba4_core_144;
  wire popcount36_2ba4_core_145;
  wire popcount36_2ba4_core_146;
  wire popcount36_2ba4_core_147;
  wire popcount36_2ba4_core_148;
  wire popcount36_2ba4_core_149;
  wire popcount36_2ba4_core_150;
  wire popcount36_2ba4_core_151;
  wire popcount36_2ba4_core_152;
  wire popcount36_2ba4_core_153;
  wire popcount36_2ba4_core_154_not;
  wire popcount36_2ba4_core_155;
  wire popcount36_2ba4_core_156;
  wire popcount36_2ba4_core_157;
  wire popcount36_2ba4_core_158;
  wire popcount36_2ba4_core_159;
  wire popcount36_2ba4_core_160;
  wire popcount36_2ba4_core_161;
  wire popcount36_2ba4_core_162;
  wire popcount36_2ba4_core_163;
  wire popcount36_2ba4_core_164;
  wire popcount36_2ba4_core_165;
  wire popcount36_2ba4_core_166;
  wire popcount36_2ba4_core_167;
  wire popcount36_2ba4_core_168;
  wire popcount36_2ba4_core_169;
  wire popcount36_2ba4_core_170;
  wire popcount36_2ba4_core_173;
  wire popcount36_2ba4_core_174;
  wire popcount36_2ba4_core_176;
  wire popcount36_2ba4_core_177;
  wire popcount36_2ba4_core_186;
  wire popcount36_2ba4_core_187;
  wire popcount36_2ba4_core_188;
  wire popcount36_2ba4_core_189;
  wire popcount36_2ba4_core_190;
  wire popcount36_2ba4_core_191;
  wire popcount36_2ba4_core_192;
  wire popcount36_2ba4_core_193;
  wire popcount36_2ba4_core_194;
  wire popcount36_2ba4_core_197;
  wire popcount36_2ba4_core_198;
  wire popcount36_2ba4_core_199;
  wire popcount36_2ba4_core_200;
  wire popcount36_2ba4_core_201;
  wire popcount36_2ba4_core_202;
  wire popcount36_2ba4_core_203;
  wire popcount36_2ba4_core_204;
  wire popcount36_2ba4_core_205;
  wire popcount36_2ba4_core_207;
  wire popcount36_2ba4_core_208;
  wire popcount36_2ba4_core_209;
  wire popcount36_2ba4_core_212;
  wire popcount36_2ba4_core_213;
  wire popcount36_2ba4_core_214;
  wire popcount36_2ba4_core_215;
  wire popcount36_2ba4_core_216;
  wire popcount36_2ba4_core_217;
  wire popcount36_2ba4_core_218;
  wire popcount36_2ba4_core_219;
  wire popcount36_2ba4_core_220;
  wire popcount36_2ba4_core_221;
  wire popcount36_2ba4_core_223;
  wire popcount36_2ba4_core_224;
  wire popcount36_2ba4_core_226;
  wire popcount36_2ba4_core_227;
  wire popcount36_2ba4_core_228;
  wire popcount36_2ba4_core_229;
  wire popcount36_2ba4_core_230;
  wire popcount36_2ba4_core_231;
  wire popcount36_2ba4_core_232;
  wire popcount36_2ba4_core_233;
  wire popcount36_2ba4_core_234;
  wire popcount36_2ba4_core_235;
  wire popcount36_2ba4_core_236;
  wire popcount36_2ba4_core_237;
  wire popcount36_2ba4_core_238;
  wire popcount36_2ba4_core_239;
  wire popcount36_2ba4_core_240;
  wire popcount36_2ba4_core_241;
  wire popcount36_2ba4_core_242;
  wire popcount36_2ba4_core_243;
  wire popcount36_2ba4_core_244;
  wire popcount36_2ba4_core_247;
  wire popcount36_2ba4_core_248;
  wire popcount36_2ba4_core_250;
  wire popcount36_2ba4_core_257;
  wire popcount36_2ba4_core_258;
  wire popcount36_2ba4_core_259;
  wire popcount36_2ba4_core_260;
  wire popcount36_2ba4_core_261;
  wire popcount36_2ba4_core_262;
  wire popcount36_2ba4_core_263;
  wire popcount36_2ba4_core_264;
  wire popcount36_2ba4_core_265;
  wire popcount36_2ba4_core_266;
  wire popcount36_2ba4_core_267;
  wire popcount36_2ba4_core_268;
  wire popcount36_2ba4_core_269;
  wire popcount36_2ba4_core_270;
  wire popcount36_2ba4_core_271;
  wire popcount36_2ba4_core_274;
  wire popcount36_2ba4_core_275;

  assign popcount36_2ba4_core_038 = input_a[32] ^ input_a[1];
  assign popcount36_2ba4_core_039 = input_a[0] & input_a[7];
  assign popcount36_2ba4_core_040 = input_a[2] ^ input_a[3];
  assign popcount36_2ba4_core_041 = input_a[2] & input_a[3];
  assign popcount36_2ba4_core_042 = popcount36_2ba4_core_038 | popcount36_2ba4_core_040;
  assign popcount36_2ba4_core_043 = ~popcount36_2ba4_core_038;
  assign popcount36_2ba4_core_044 = popcount36_2ba4_core_039 ^ popcount36_2ba4_core_041;
  assign popcount36_2ba4_core_046 = popcount36_2ba4_core_044 ^ popcount36_2ba4_core_043;
  assign popcount36_2ba4_core_048 = popcount36_2ba4_core_039 | input_a[18];
  assign popcount36_2ba4_core_050 = input_a[10] & input_a[5];
  assign popcount36_2ba4_core_051 = ~input_a[7];
  assign popcount36_2ba4_core_052 = input_a[7] & input_a[8];
  assign popcount36_2ba4_core_053 = input_a[13] ^ input_a[27];
  assign popcount36_2ba4_core_054 = input_a[22] & popcount36_2ba4_core_051;
  assign popcount36_2ba4_core_056 = popcount36_2ba4_core_052 & popcount36_2ba4_core_054;
  assign popcount36_2ba4_core_057 = input_a[24] ^ popcount36_2ba4_core_053;
  assign popcount36_2ba4_core_058 = input_a[5] & popcount36_2ba4_core_053;
  assign popcount36_2ba4_core_061 = input_a[32] ^ input_a[24];
  assign popcount36_2ba4_core_062 = input_a[32] ^ input_a[13];
  assign popcount36_2ba4_core_066 = popcount36_2ba4_core_042 ^ popcount36_2ba4_core_057;
  assign popcount36_2ba4_core_067 = input_a[33] & input_a[31];
  assign popcount36_2ba4_core_068 = ~(popcount36_2ba4_core_046 | input_a[25]);
  assign popcount36_2ba4_core_069 = popcount36_2ba4_core_046 & input_a[1];
  assign popcount36_2ba4_core_070 = popcount36_2ba4_core_068 & popcount36_2ba4_core_067;
  assign popcount36_2ba4_core_071 = input_a[20] & popcount36_2ba4_core_067;
  assign popcount36_2ba4_core_072 = popcount36_2ba4_core_069 | popcount36_2ba4_core_071;
  assign popcount36_2ba4_core_081 = input_a[8] & input_a[10];
  assign popcount36_2ba4_core_082 = input_a[35] ^ input_a[12];
  assign popcount36_2ba4_core_083 = input_a[21] & input_a[12];
  assign popcount36_2ba4_core_084 = ~input_a[30];
  assign popcount36_2ba4_core_086 = popcount36_2ba4_core_081 ^ input_a[25];
  assign popcount36_2ba4_core_087 = popcount36_2ba4_core_081 & popcount36_2ba4_core_083;
  assign popcount36_2ba4_core_088 = popcount36_2ba4_core_086 ^ input_a[33];
  assign popcount36_2ba4_core_089 = popcount36_2ba4_core_086 & input_a[31];
  assign popcount36_2ba4_core_090 = popcount36_2ba4_core_087 | input_a[16];
  assign popcount36_2ba4_core_091 = input_a[31] ^ input_a[14];
  assign popcount36_2ba4_core_092 = input_a[13] & input_a[14];
  assign popcount36_2ba4_core_093 = input_a[13] ^ input_a[17];
  assign popcount36_2ba4_core_096 = input_a[32] & input_a[18];
  assign popcount36_2ba4_core_099_not = ~popcount36_2ba4_core_091;
  assign popcount36_2ba4_core_101 = popcount36_2ba4_core_092 ^ input_a[27];
  assign popcount36_2ba4_core_102 = popcount36_2ba4_core_092 | input_a[27];
  assign popcount36_2ba4_core_103 = popcount36_2ba4_core_101 ^ popcount36_2ba4_core_091;
  assign popcount36_2ba4_core_104 = input_a[13] & input_a[19];
  assign popcount36_2ba4_core_105 = input_a[21] | popcount36_2ba4_core_104;
  assign popcount36_2ba4_core_106 = input_a[17] ^ popcount36_2ba4_core_105;
  assign popcount36_2ba4_core_110 = popcount36_2ba4_core_088 ^ popcount36_2ba4_core_103;
  assign popcount36_2ba4_core_111 = popcount36_2ba4_core_088 & input_a[18];
  assign popcount36_2ba4_core_115 = popcount36_2ba4_core_090 ^ popcount36_2ba4_core_106;
  assign popcount36_2ba4_core_116 = popcount36_2ba4_core_090 & popcount36_2ba4_core_106;
  assign popcount36_2ba4_core_117 = popcount36_2ba4_core_115 ^ popcount36_2ba4_core_111;
  assign popcount36_2ba4_core_118 = popcount36_2ba4_core_115 & popcount36_2ba4_core_111;
  assign popcount36_2ba4_core_119 = popcount36_2ba4_core_116 | popcount36_2ba4_core_118;
  assign popcount36_2ba4_core_124 = popcount36_2ba4_core_070 ^ input_a[34];
  assign popcount36_2ba4_core_125 = input_a[22] & input_a[34];
  assign popcount36_2ba4_core_128 = popcount36_2ba4_core_125 | input_a[11];
  assign popcount36_2ba4_core_129 = popcount36_2ba4_core_072 ^ popcount36_2ba4_core_117;
  assign popcount36_2ba4_core_131 = popcount36_2ba4_core_129 ^ popcount36_2ba4_core_128;
  assign popcount36_2ba4_core_132 = popcount36_2ba4_core_129 & popcount36_2ba4_core_128;
  assign popcount36_2ba4_core_136 = ~(popcount36_2ba4_core_119 & popcount36_2ba4_core_132);
  assign popcount36_2ba4_core_137 = popcount36_2ba4_core_119 & popcount36_2ba4_core_132;
  assign popcount36_2ba4_core_144 = input_a[8] ^ input_a[19];
  assign popcount36_2ba4_core_145 = ~(input_a[14] & input_a[27]);
  assign popcount36_2ba4_core_146 = input_a[20] ^ input_a[21];
  assign popcount36_2ba4_core_147 = input_a[24] & input_a[21];
  assign popcount36_2ba4_core_148 = input_a[21] ^ input_a[22];
  assign popcount36_2ba4_core_149 = ~(input_a[23] | popcount36_2ba4_core_146);
  assign popcount36_2ba4_core_150 = input_a[9] ^ popcount36_2ba4_core_147;
  assign popcount36_2ba4_core_151 = popcount36_2ba4_core_145 & input_a[19];
  assign popcount36_2ba4_core_152 = popcount36_2ba4_core_150 & input_a[29];
  assign popcount36_2ba4_core_153 = ~(input_a[26] | popcount36_2ba4_core_149);
  assign popcount36_2ba4_core_154_not = ~popcount36_2ba4_core_153;
  assign popcount36_2ba4_core_155 = input_a[22] ^ input_a[23];
  assign popcount36_2ba4_core_156 = input_a[12] & input_a[34];
  assign popcount36_2ba4_core_157 = input_a[25] | input_a[6];
  assign popcount36_2ba4_core_158 = input_a[25] & input_a[34];
  assign popcount36_2ba4_core_159 = input_a[24] ^ input_a[5];
  assign popcount36_2ba4_core_160 = input_a[24] & input_a[30];
  assign popcount36_2ba4_core_161 = popcount36_2ba4_core_158 ^ input_a[16];
  assign popcount36_2ba4_core_162 = popcount36_2ba4_core_158 & popcount36_2ba4_core_160;
  assign popcount36_2ba4_core_163 = input_a[28] ^ popcount36_2ba4_core_159;
  assign popcount36_2ba4_core_164 = input_a[22] & popcount36_2ba4_core_159;
  assign popcount36_2ba4_core_165 = popcount36_2ba4_core_156 ^ popcount36_2ba4_core_161;
  assign popcount36_2ba4_core_166 = ~(popcount36_2ba4_core_156 | input_a[20]);
  assign popcount36_2ba4_core_167 = input_a[35] ^ popcount36_2ba4_core_164;
  assign popcount36_2ba4_core_168 = ~(popcount36_2ba4_core_165 ^ popcount36_2ba4_core_164);
  assign popcount36_2ba4_core_169 = input_a[27] | popcount36_2ba4_core_168;
  assign popcount36_2ba4_core_170 = ~(popcount36_2ba4_core_162 ^ input_a[30]);
  assign popcount36_2ba4_core_173 = input_a[32] & popcount36_2ba4_core_163;
  assign popcount36_2ba4_core_174 = input_a[12] & popcount36_2ba4_core_167;
  assign popcount36_2ba4_core_176 = popcount36_2ba4_core_174 ^ popcount36_2ba4_core_173;
  assign popcount36_2ba4_core_177 = popcount36_2ba4_core_174 & popcount36_2ba4_core_173;
  assign popcount36_2ba4_core_186 = ~(input_a[27] | input_a[28]);
  assign popcount36_2ba4_core_187 = input_a[27] & input_a[9];
  assign popcount36_2ba4_core_188 = input_a[5] ^ input_a[5];
  assign popcount36_2ba4_core_189 = input_a[16] & input_a[30];
  assign popcount36_2ba4_core_190 = popcount36_2ba4_core_186 ^ popcount36_2ba4_core_188;
  assign popcount36_2ba4_core_191 = popcount36_2ba4_core_186 & popcount36_2ba4_core_188;
  assign popcount36_2ba4_core_192 = popcount36_2ba4_core_187 ^ input_a[24];
  assign popcount36_2ba4_core_193 = popcount36_2ba4_core_187 & popcount36_2ba4_core_189;
  assign popcount36_2ba4_core_194 = popcount36_2ba4_core_192 ^ popcount36_2ba4_core_191;
  assign popcount36_2ba4_core_197 = input_a[31] ^ input_a[33];
  assign popcount36_2ba4_core_198 = input_a[33] & input_a[32];
  assign popcount36_2ba4_core_199 = input_a[34] ^ input_a[35];
  assign popcount36_2ba4_core_200 = input_a[34] & input_a[35];
  assign popcount36_2ba4_core_201 = ~(input_a[33] ^ input_a[14]);
  assign popcount36_2ba4_core_202 = input_a[33] & popcount36_2ba4_core_199;
  assign popcount36_2ba4_core_203 = popcount36_2ba4_core_200 & popcount36_2ba4_core_202;
  assign popcount36_2ba4_core_204 = popcount36_2ba4_core_200 & popcount36_2ba4_core_202;
  assign popcount36_2ba4_core_205 = input_a[35] ^ input_a[18];
  assign popcount36_2ba4_core_207 = popcount36_2ba4_core_198 ^ popcount36_2ba4_core_203;
  assign popcount36_2ba4_core_208 = popcount36_2ba4_core_198 & popcount36_2ba4_core_203;
  assign popcount36_2ba4_core_209 = input_a[33] ^ input_a[29];
  assign popcount36_2ba4_core_212 = popcount36_2ba4_core_204 ^ popcount36_2ba4_core_208;
  assign popcount36_2ba4_core_213 = popcount36_2ba4_core_204 & input_a[1];
  assign popcount36_2ba4_core_214 = input_a[30] ^ input_a[17];
  assign popcount36_2ba4_core_215 = input_a[2] & popcount36_2ba4_core_205;
  assign popcount36_2ba4_core_216 = ~(popcount36_2ba4_core_194 & popcount36_2ba4_core_209);
  assign popcount36_2ba4_core_217 = popcount36_2ba4_core_194 & popcount36_2ba4_core_209;
  assign popcount36_2ba4_core_218 = popcount36_2ba4_core_216 ^ popcount36_2ba4_core_215;
  assign popcount36_2ba4_core_219 = popcount36_2ba4_core_216 & popcount36_2ba4_core_215;
  assign popcount36_2ba4_core_220 = popcount36_2ba4_core_217 | popcount36_2ba4_core_219;
  assign popcount36_2ba4_core_221 = popcount36_2ba4_core_193 ^ popcount36_2ba4_core_212;
  assign popcount36_2ba4_core_223 = popcount36_2ba4_core_221 ^ popcount36_2ba4_core_220;
  assign popcount36_2ba4_core_224 = popcount36_2ba4_core_221 & popcount36_2ba4_core_220;
  assign popcount36_2ba4_core_226 = popcount36_2ba4_core_213 ^ popcount36_2ba4_core_224;
  assign popcount36_2ba4_core_227 = popcount36_2ba4_core_213 & popcount36_2ba4_core_224;
  assign popcount36_2ba4_core_228 = input_a[22] | popcount36_2ba4_core_214;
  assign popcount36_2ba4_core_229 = input_a[22] & input_a[23];
  assign popcount36_2ba4_core_230 = popcount36_2ba4_core_176 ^ popcount36_2ba4_core_218;
  assign popcount36_2ba4_core_231 = popcount36_2ba4_core_176 & popcount36_2ba4_core_218;
  assign popcount36_2ba4_core_232 = popcount36_2ba4_core_230 ^ popcount36_2ba4_core_229;
  assign popcount36_2ba4_core_233 = input_a[31] & popcount36_2ba4_core_229;
  assign popcount36_2ba4_core_234 = popcount36_2ba4_core_231 | popcount36_2ba4_core_233;
  assign popcount36_2ba4_core_235 = popcount36_2ba4_core_177 ^ popcount36_2ba4_core_223;
  assign popcount36_2ba4_core_236 = popcount36_2ba4_core_177 & popcount36_2ba4_core_223;
  assign popcount36_2ba4_core_237 = popcount36_2ba4_core_235 ^ popcount36_2ba4_core_234;
  assign popcount36_2ba4_core_238 = popcount36_2ba4_core_235 & popcount36_2ba4_core_234;
  assign popcount36_2ba4_core_239 = popcount36_2ba4_core_236 | popcount36_2ba4_core_238;
  assign popcount36_2ba4_core_240 = popcount36_2ba4_core_162 ^ popcount36_2ba4_core_226;
  assign popcount36_2ba4_core_241 = popcount36_2ba4_core_162 & input_a[16];
  assign popcount36_2ba4_core_242 = popcount36_2ba4_core_240 ^ popcount36_2ba4_core_239;
  assign popcount36_2ba4_core_243 = ~(popcount36_2ba4_core_240 & popcount36_2ba4_core_239);
  assign popcount36_2ba4_core_244 = ~popcount36_2ba4_core_241;
  assign popcount36_2ba4_core_247 = popcount36_2ba4_core_227 & input_a[2];
  assign popcount36_2ba4_core_248 = popcount36_2ba4_core_227 & input_a[2];
  assign popcount36_2ba4_core_250 = input_a[34] ^ input_a[32];
  assign popcount36_2ba4_core_257 = popcount36_2ba4_core_131 ^ popcount36_2ba4_core_237;
  assign popcount36_2ba4_core_258 = popcount36_2ba4_core_131 & popcount36_2ba4_core_237;
  assign popcount36_2ba4_core_259 = popcount36_2ba4_core_257 ^ popcount36_2ba4_core_232;
  assign popcount36_2ba4_core_260 = popcount36_2ba4_core_257 & popcount36_2ba4_core_232;
  assign popcount36_2ba4_core_261 = popcount36_2ba4_core_258 | popcount36_2ba4_core_260;
  assign popcount36_2ba4_core_262 = popcount36_2ba4_core_136 ^ popcount36_2ba4_core_242;
  assign popcount36_2ba4_core_263 = popcount36_2ba4_core_136 & popcount36_2ba4_core_242;
  assign popcount36_2ba4_core_264 = popcount36_2ba4_core_262 ^ popcount36_2ba4_core_261;
  assign popcount36_2ba4_core_265 = popcount36_2ba4_core_262 & popcount36_2ba4_core_261;
  assign popcount36_2ba4_core_266 = popcount36_2ba4_core_263 | popcount36_2ba4_core_265;
  assign popcount36_2ba4_core_267 = popcount36_2ba4_core_137 ^ popcount36_2ba4_core_247;
  assign popcount36_2ba4_core_268 = popcount36_2ba4_core_137 & popcount36_2ba4_core_247;
  assign popcount36_2ba4_core_269 = popcount36_2ba4_core_267 ^ popcount36_2ba4_core_266;
  assign popcount36_2ba4_core_270 = popcount36_2ba4_core_267 & popcount36_2ba4_core_266;
  assign popcount36_2ba4_core_271 = popcount36_2ba4_core_268 | popcount36_2ba4_core_270;
  assign popcount36_2ba4_core_274 = popcount36_2ba4_core_248 ^ popcount36_2ba4_core_271;
  assign popcount36_2ba4_core_275 = popcount36_2ba4_core_248 & popcount36_2ba4_core_271;

  assign popcount36_2ba4_out[0] = 1'b1;
  assign popcount36_2ba4_out[1] = 1'b0;
  assign popcount36_2ba4_out[2] = popcount36_2ba4_core_259;
  assign popcount36_2ba4_out[3] = popcount36_2ba4_core_264;
  assign popcount36_2ba4_out[4] = popcount36_2ba4_core_269;
  assign popcount36_2ba4_out[5] = popcount36_2ba4_core_274;
endmodule