// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.37709
// WCE=18.0
// EP=0.867939%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_up9p(input [35:0] input_a, output [5:0] popcount36_up9p_out);
  wire popcount36_up9p_core_038;
  wire popcount36_up9p_core_039;
  wire popcount36_up9p_core_040;
  wire popcount36_up9p_core_041;
  wire popcount36_up9p_core_043;
  wire popcount36_up9p_core_044;
  wire popcount36_up9p_core_045;
  wire popcount36_up9p_core_047;
  wire popcount36_up9p_core_048;
  wire popcount36_up9p_core_049;
  wire popcount36_up9p_core_050;
  wire popcount36_up9p_core_052;
  wire popcount36_up9p_core_054;
  wire popcount36_up9p_core_055;
  wire popcount36_up9p_core_056;
  wire popcount36_up9p_core_057;
  wire popcount36_up9p_core_059;
  wire popcount36_up9p_core_060;
  wire popcount36_up9p_core_061;
  wire popcount36_up9p_core_062;
  wire popcount36_up9p_core_063;
  wire popcount36_up9p_core_064;
  wire popcount36_up9p_core_065_not;
  wire popcount36_up9p_core_068;
  wire popcount36_up9p_core_070;
  wire popcount36_up9p_core_071;
  wire popcount36_up9p_core_072;
  wire popcount36_up9p_core_075;
  wire popcount36_up9p_core_076;
  wire popcount36_up9p_core_077;
  wire popcount36_up9p_core_080;
  wire popcount36_up9p_core_082;
  wire popcount36_up9p_core_083;
  wire popcount36_up9p_core_084;
  wire popcount36_up9p_core_086;
  wire popcount36_up9p_core_091;
  wire popcount36_up9p_core_092;
  wire popcount36_up9p_core_093;
  wire popcount36_up9p_core_096;
  wire popcount36_up9p_core_098;
  wire popcount36_up9p_core_100;
  wire popcount36_up9p_core_101;
  wire popcount36_up9p_core_103;
  wire popcount36_up9p_core_105;
  wire popcount36_up9p_core_106;
  wire popcount36_up9p_core_107;
  wire popcount36_up9p_core_108;
  wire popcount36_up9p_core_109;
  wire popcount36_up9p_core_111_not;
  wire popcount36_up9p_core_112;
  wire popcount36_up9p_core_117;
  wire popcount36_up9p_core_118;
  wire popcount36_up9p_core_120;
  wire popcount36_up9p_core_121;
  wire popcount36_up9p_core_122;
  wire popcount36_up9p_core_124;
  wire popcount36_up9p_core_125;
  wire popcount36_up9p_core_126;
  wire popcount36_up9p_core_128;
  wire popcount36_up9p_core_131;
  wire popcount36_up9p_core_132;
  wire popcount36_up9p_core_133;
  wire popcount36_up9p_core_135;
  wire popcount36_up9p_core_136;
  wire popcount36_up9p_core_137;
  wire popcount36_up9p_core_138;
  wire popcount36_up9p_core_139;
  wire popcount36_up9p_core_142;
  wire popcount36_up9p_core_143;
  wire popcount36_up9p_core_146;
  wire popcount36_up9p_core_149;
  wire popcount36_up9p_core_152;
  wire popcount36_up9p_core_153;
  wire popcount36_up9p_core_154;
  wire popcount36_up9p_core_155;
  wire popcount36_up9p_core_156;
  wire popcount36_up9p_core_157;
  wire popcount36_up9p_core_158;
  wire popcount36_up9p_core_159;
  wire popcount36_up9p_core_161;
  wire popcount36_up9p_core_164;
  wire popcount36_up9p_core_165;
  wire popcount36_up9p_core_166;
  wire popcount36_up9p_core_167;
  wire popcount36_up9p_core_168;
  wire popcount36_up9p_core_169;
  wire popcount36_up9p_core_170;
  wire popcount36_up9p_core_172;
  wire popcount36_up9p_core_173;
  wire popcount36_up9p_core_174;
  wire popcount36_up9p_core_175;
  wire popcount36_up9p_core_180;
  wire popcount36_up9p_core_182;
  wire popcount36_up9p_core_185;
  wire popcount36_up9p_core_186;
  wire popcount36_up9p_core_187;
  wire popcount36_up9p_core_188_not;
  wire popcount36_up9p_core_190;
  wire popcount36_up9p_core_191;
  wire popcount36_up9p_core_192;
  wire popcount36_up9p_core_193;
  wire popcount36_up9p_core_195;
  wire popcount36_up9p_core_197;
  wire popcount36_up9p_core_198;
  wire popcount36_up9p_core_199;
  wire popcount36_up9p_core_202;
  wire popcount36_up9p_core_203;
  wire popcount36_up9p_core_204;
  wire popcount36_up9p_core_205;
  wire popcount36_up9p_core_206;
  wire popcount36_up9p_core_207;
  wire popcount36_up9p_core_208;
  wire popcount36_up9p_core_210;
  wire popcount36_up9p_core_212_not;
  wire popcount36_up9p_core_213;
  wire popcount36_up9p_core_214;
  wire popcount36_up9p_core_216;
  wire popcount36_up9p_core_218;
  wire popcount36_up9p_core_220;
  wire popcount36_up9p_core_221_not;
  wire popcount36_up9p_core_223_not;
  wire popcount36_up9p_core_224;
  wire popcount36_up9p_core_228;
  wire popcount36_up9p_core_229;
  wire popcount36_up9p_core_230;
  wire popcount36_up9p_core_231;
  wire popcount36_up9p_core_237;
  wire popcount36_up9p_core_238;
  wire popcount36_up9p_core_239;
  wire popcount36_up9p_core_240;
  wire popcount36_up9p_core_243;
  wire popcount36_up9p_core_244;
  wire popcount36_up9p_core_245;
  wire popcount36_up9p_core_246;
  wire popcount36_up9p_core_247;
  wire popcount36_up9p_core_251;
  wire popcount36_up9p_core_253;
  wire popcount36_up9p_core_254_not;
  wire popcount36_up9p_core_255;
  wire popcount36_up9p_core_258;
  wire popcount36_up9p_core_259;
  wire popcount36_up9p_core_260;
  wire popcount36_up9p_core_261;
  wire popcount36_up9p_core_263;
  wire popcount36_up9p_core_264;
  wire popcount36_up9p_core_266;
  wire popcount36_up9p_core_267;
  wire popcount36_up9p_core_270;
  wire popcount36_up9p_core_272;
  wire popcount36_up9p_core_276;

  assign popcount36_up9p_core_038 = input_a[26] ^ input_a[27];
  assign popcount36_up9p_core_039 = ~(input_a[29] | input_a[16]);
  assign popcount36_up9p_core_040 = input_a[33] ^ input_a[14];
  assign popcount36_up9p_core_041 = input_a[27] ^ input_a[33];
  assign popcount36_up9p_core_043 = input_a[25] & input_a[9];
  assign popcount36_up9p_core_044 = ~input_a[21];
  assign popcount36_up9p_core_045 = ~input_a[25];
  assign popcount36_up9p_core_047 = ~(input_a[4] & input_a[10]);
  assign popcount36_up9p_core_048 = ~input_a[34];
  assign popcount36_up9p_core_049 = input_a[4] | input_a[31];
  assign popcount36_up9p_core_050 = ~(input_a[2] | input_a[30]);
  assign popcount36_up9p_core_052 = input_a[18] | input_a[16];
  assign popcount36_up9p_core_054 = input_a[30] | input_a[29];
  assign popcount36_up9p_core_055 = ~(input_a[12] ^ input_a[12]);
  assign popcount36_up9p_core_056 = ~(input_a[3] & input_a[22]);
  assign popcount36_up9p_core_057 = ~input_a[5];
  assign popcount36_up9p_core_059 = ~(input_a[6] & input_a[31]);
  assign popcount36_up9p_core_060 = input_a[24] | input_a[18];
  assign popcount36_up9p_core_061 = input_a[34] & input_a[17];
  assign popcount36_up9p_core_062 = input_a[20] ^ input_a[27];
  assign popcount36_up9p_core_063 = input_a[35] | input_a[31];
  assign popcount36_up9p_core_064 = ~input_a[18];
  assign popcount36_up9p_core_065_not = ~input_a[3];
  assign popcount36_up9p_core_068 = ~(input_a[9] ^ input_a[16]);
  assign popcount36_up9p_core_070 = ~(input_a[17] | input_a[34]);
  assign popcount36_up9p_core_071 = ~(input_a[1] | input_a[17]);
  assign popcount36_up9p_core_072 = ~(input_a[14] ^ input_a[6]);
  assign popcount36_up9p_core_075 = ~(input_a[16] | input_a[11]);
  assign popcount36_up9p_core_076 = input_a[31] | input_a[7];
  assign popcount36_up9p_core_077 = ~(input_a[29] ^ input_a[25]);
  assign popcount36_up9p_core_080 = ~(input_a[0] | input_a[26]);
  assign popcount36_up9p_core_082 = ~input_a[3];
  assign popcount36_up9p_core_083 = input_a[2] ^ input_a[26];
  assign popcount36_up9p_core_084 = input_a[32] | input_a[13];
  assign popcount36_up9p_core_086 = input_a[17] ^ input_a[6];
  assign popcount36_up9p_core_091 = ~(input_a[20] ^ input_a[10]);
  assign popcount36_up9p_core_092 = ~(input_a[14] | input_a[27]);
  assign popcount36_up9p_core_093 = input_a[1] | input_a[33];
  assign popcount36_up9p_core_096 = ~(input_a[1] & input_a[10]);
  assign popcount36_up9p_core_098 = ~(input_a[5] ^ input_a[9]);
  assign popcount36_up9p_core_100 = input_a[27] ^ input_a[6];
  assign popcount36_up9p_core_101 = ~(input_a[34] & input_a[15]);
  assign popcount36_up9p_core_103 = input_a[9] & input_a[35];
  assign popcount36_up9p_core_105 = input_a[24] | input_a[11];
  assign popcount36_up9p_core_106 = input_a[34] & input_a[22];
  assign popcount36_up9p_core_107 = input_a[9] & input_a[11];
  assign popcount36_up9p_core_108 = ~(input_a[5] ^ input_a[0]);
  assign popcount36_up9p_core_109 = input_a[20] ^ input_a[22];
  assign popcount36_up9p_core_111_not = ~input_a[19];
  assign popcount36_up9p_core_112 = input_a[21] & input_a[11];
  assign popcount36_up9p_core_117 = ~input_a[35];
  assign popcount36_up9p_core_118 = ~input_a[2];
  assign popcount36_up9p_core_120 = ~(input_a[8] ^ input_a[29]);
  assign popcount36_up9p_core_121 = ~input_a[5];
  assign popcount36_up9p_core_122 = input_a[17] & input_a[21];
  assign popcount36_up9p_core_124 = ~(input_a[1] ^ input_a[25]);
  assign popcount36_up9p_core_125 = input_a[28] | input_a[28];
  assign popcount36_up9p_core_126 = ~(input_a[31] | input_a[14]);
  assign popcount36_up9p_core_128 = ~(input_a[20] ^ input_a[26]);
  assign popcount36_up9p_core_131 = ~(input_a[15] ^ input_a[4]);
  assign popcount36_up9p_core_132 = ~(input_a[17] & input_a[30]);
  assign popcount36_up9p_core_133 = input_a[10] & input_a[30];
  assign popcount36_up9p_core_135 = input_a[35] ^ input_a[34];
  assign popcount36_up9p_core_136 = input_a[6] & input_a[7];
  assign popcount36_up9p_core_137 = ~(input_a[24] ^ input_a[29]);
  assign popcount36_up9p_core_138 = ~input_a[30];
  assign popcount36_up9p_core_139 = ~(input_a[1] ^ input_a[7]);
  assign popcount36_up9p_core_142 = ~(input_a[12] | input_a[23]);
  assign popcount36_up9p_core_143 = ~input_a[28];
  assign popcount36_up9p_core_146 = input_a[32] | input_a[9];
  assign popcount36_up9p_core_149 = input_a[25] | input_a[14];
  assign popcount36_up9p_core_152 = ~(input_a[11] ^ input_a[21]);
  assign popcount36_up9p_core_153 = input_a[11] | input_a[16];
  assign popcount36_up9p_core_154 = ~(input_a[27] ^ input_a[8]);
  assign popcount36_up9p_core_155 = ~input_a[28];
  assign popcount36_up9p_core_156 = input_a[17] & input_a[7];
  assign popcount36_up9p_core_157 = input_a[1] | input_a[18];
  assign popcount36_up9p_core_158 = ~(input_a[9] & input_a[5]);
  assign popcount36_up9p_core_159 = ~(input_a[30] & input_a[12]);
  assign popcount36_up9p_core_161 = input_a[8] ^ input_a[15];
  assign popcount36_up9p_core_164 = input_a[4] | input_a[6];
  assign popcount36_up9p_core_165 = ~(input_a[11] & input_a[4]);
  assign popcount36_up9p_core_166 = input_a[35] ^ input_a[23];
  assign popcount36_up9p_core_167 = ~(input_a[0] ^ input_a[13]);
  assign popcount36_up9p_core_168 = ~input_a[25];
  assign popcount36_up9p_core_169 = input_a[6] ^ input_a[23];
  assign popcount36_up9p_core_170 = ~input_a[17];
  assign popcount36_up9p_core_172 = input_a[23] & input_a[27];
  assign popcount36_up9p_core_173 = ~(input_a[25] ^ input_a[27]);
  assign popcount36_up9p_core_174 = input_a[19] & input_a[16];
  assign popcount36_up9p_core_175 = ~(input_a[9] ^ input_a[27]);
  assign popcount36_up9p_core_180 = ~(input_a[0] & input_a[9]);
  assign popcount36_up9p_core_182 = ~(input_a[18] & input_a[31]);
  assign popcount36_up9p_core_185 = input_a[16] & input_a[14];
  assign popcount36_up9p_core_186 = ~input_a[11];
  assign popcount36_up9p_core_187 = ~(input_a[22] ^ input_a[5]);
  assign popcount36_up9p_core_188_not = ~input_a[23];
  assign popcount36_up9p_core_190 = ~(input_a[25] | input_a[22]);
  assign popcount36_up9p_core_191 = ~input_a[20];
  assign popcount36_up9p_core_192 = ~input_a[30];
  assign popcount36_up9p_core_193 = ~(input_a[2] & input_a[35]);
  assign popcount36_up9p_core_195 = ~(input_a[4] | input_a[17]);
  assign popcount36_up9p_core_197 = ~(input_a[13] | input_a[14]);
  assign popcount36_up9p_core_198 = ~(input_a[28] | input_a[11]);
  assign popcount36_up9p_core_199 = ~(input_a[21] | input_a[16]);
  assign popcount36_up9p_core_202 = input_a[16] ^ input_a[19];
  assign popcount36_up9p_core_203 = ~input_a[13];
  assign popcount36_up9p_core_204 = input_a[20] & input_a[16];
  assign popcount36_up9p_core_205 = ~input_a[14];
  assign popcount36_up9p_core_206 = ~(input_a[13] | input_a[14]);
  assign popcount36_up9p_core_207 = input_a[22] & input_a[30];
  assign popcount36_up9p_core_208 = input_a[4] | input_a[15];
  assign popcount36_up9p_core_210 = ~(input_a[2] & input_a[22]);
  assign popcount36_up9p_core_212_not = ~input_a[35];
  assign popcount36_up9p_core_213 = ~(input_a[20] | input_a[20]);
  assign popcount36_up9p_core_214 = ~(input_a[19] | input_a[26]);
  assign popcount36_up9p_core_216 = ~(input_a[20] & input_a[30]);
  assign popcount36_up9p_core_218 = input_a[2] | input_a[2];
  assign popcount36_up9p_core_220 = ~(input_a[30] & input_a[4]);
  assign popcount36_up9p_core_221_not = ~input_a[15];
  assign popcount36_up9p_core_223_not = ~input_a[12];
  assign popcount36_up9p_core_224 = input_a[11] ^ input_a[15];
  assign popcount36_up9p_core_228 = input_a[22] | input_a[15];
  assign popcount36_up9p_core_229 = ~input_a[17];
  assign popcount36_up9p_core_230 = input_a[8] | input_a[8];
  assign popcount36_up9p_core_231 = ~(input_a[7] & input_a[16]);
  assign popcount36_up9p_core_237 = ~input_a[21];
  assign popcount36_up9p_core_238 = input_a[31] | input_a[0];
  assign popcount36_up9p_core_239 = ~(input_a[28] & input_a[11]);
  assign popcount36_up9p_core_240 = input_a[19] & input_a[33];
  assign popcount36_up9p_core_243 = input_a[18] | input_a[19];
  assign popcount36_up9p_core_244 = input_a[14] & input_a[35];
  assign popcount36_up9p_core_245 = ~input_a[5];
  assign popcount36_up9p_core_246 = ~(input_a[23] | input_a[0]);
  assign popcount36_up9p_core_247 = ~input_a[25];
  assign popcount36_up9p_core_251 = ~(input_a[15] ^ input_a[14]);
  assign popcount36_up9p_core_253 = input_a[3] & input_a[35];
  assign popcount36_up9p_core_254_not = ~input_a[20];
  assign popcount36_up9p_core_255 = ~input_a[32];
  assign popcount36_up9p_core_258 = ~(input_a[23] & input_a[29]);
  assign popcount36_up9p_core_259 = input_a[15] ^ input_a[35];
  assign popcount36_up9p_core_260 = ~input_a[20];
  assign popcount36_up9p_core_261 = input_a[8] & input_a[14];
  assign popcount36_up9p_core_263 = input_a[32] & input_a[9];
  assign popcount36_up9p_core_264 = ~(input_a[30] | input_a[0]);
  assign popcount36_up9p_core_266 = input_a[25] & input_a[34];
  assign popcount36_up9p_core_267 = ~(input_a[7] & input_a[30]);
  assign popcount36_up9p_core_270 = input_a[24] | input_a[6];
  assign popcount36_up9p_core_272 = ~input_a[22];
  assign popcount36_up9p_core_276 = ~(input_a[22] ^ input_a[10]);

  assign popcount36_up9p_out[0] = input_a[7];
  assign popcount36_up9p_out[1] = input_a[3];
  assign popcount36_up9p_out[2] = 1'b0;
  assign popcount36_up9p_out[3] = 1'b0;
  assign popcount36_up9p_out[4] = 1'b1;
  assign popcount36_up9p_out[5] = 1'b0;
endmodule