// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.65018
// WCE=16.0
// EP=0.882934%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_qkp5(input [26:0] input_a, output [4:0] popcount27_qkp5_out);
  wire popcount27_qkp5_core_029;
  wire popcount27_qkp5_core_030;
  wire popcount27_qkp5_core_032;
  wire popcount27_qkp5_core_033;
  wire popcount27_qkp5_core_034;
  wire popcount27_qkp5_core_035;
  wire popcount27_qkp5_core_036;
  wire popcount27_qkp5_core_038;
  wire popcount27_qkp5_core_039;
  wire popcount27_qkp5_core_040;
  wire popcount27_qkp5_core_043;
  wire popcount27_qkp5_core_044;
  wire popcount27_qkp5_core_045;
  wire popcount27_qkp5_core_048;
  wire popcount27_qkp5_core_049;
  wire popcount27_qkp5_core_050;
  wire popcount27_qkp5_core_051;
  wire popcount27_qkp5_core_052;
  wire popcount27_qkp5_core_053;
  wire popcount27_qkp5_core_054;
  wire popcount27_qkp5_core_055;
  wire popcount27_qkp5_core_057;
  wire popcount27_qkp5_core_059;
  wire popcount27_qkp5_core_060;
  wire popcount27_qkp5_core_061;
  wire popcount27_qkp5_core_062;
  wire popcount27_qkp5_core_064;
  wire popcount27_qkp5_core_065;
  wire popcount27_qkp5_core_067;
  wire popcount27_qkp5_core_069;
  wire popcount27_qkp5_core_070;
  wire popcount27_qkp5_core_071;
  wire popcount27_qkp5_core_072;
  wire popcount27_qkp5_core_074;
  wire popcount27_qkp5_core_075;
  wire popcount27_qkp5_core_076;
  wire popcount27_qkp5_core_078;
  wire popcount27_qkp5_core_081;
  wire popcount27_qkp5_core_082;
  wire popcount27_qkp5_core_086;
  wire popcount27_qkp5_core_089;
  wire popcount27_qkp5_core_091;
  wire popcount27_qkp5_core_092;
  wire popcount27_qkp5_core_093;
  wire popcount27_qkp5_core_096;
  wire popcount27_qkp5_core_097;
  wire popcount27_qkp5_core_098;
  wire popcount27_qkp5_core_099;
  wire popcount27_qkp5_core_100;
  wire popcount27_qkp5_core_102;
  wire popcount27_qkp5_core_104;
  wire popcount27_qkp5_core_105;
  wire popcount27_qkp5_core_108;
  wire popcount27_qkp5_core_110;
  wire popcount27_qkp5_core_111;
  wire popcount27_qkp5_core_112;
  wire popcount27_qkp5_core_113;
  wire popcount27_qkp5_core_117;
  wire popcount27_qkp5_core_120;
  wire popcount27_qkp5_core_121;
  wire popcount27_qkp5_core_122;
  wire popcount27_qkp5_core_123;
  wire popcount27_qkp5_core_124;
  wire popcount27_qkp5_core_127;
  wire popcount27_qkp5_core_129;
  wire popcount27_qkp5_core_131_not;
  wire popcount27_qkp5_core_132;
  wire popcount27_qkp5_core_134;
  wire popcount27_qkp5_core_138;
  wire popcount27_qkp5_core_139;
  wire popcount27_qkp5_core_142;
  wire popcount27_qkp5_core_143;
  wire popcount27_qkp5_core_144;
  wire popcount27_qkp5_core_145;
  wire popcount27_qkp5_core_148;
  wire popcount27_qkp5_core_149;
  wire popcount27_qkp5_core_150;
  wire popcount27_qkp5_core_152_not;
  wire popcount27_qkp5_core_153;
  wire popcount27_qkp5_core_154;
  wire popcount27_qkp5_core_157;
  wire popcount27_qkp5_core_158;
  wire popcount27_qkp5_core_159;
  wire popcount27_qkp5_core_160;
  wire popcount27_qkp5_core_162;
  wire popcount27_qkp5_core_163;
  wire popcount27_qkp5_core_166;
  wire popcount27_qkp5_core_167;
  wire popcount27_qkp5_core_168;
  wire popcount27_qkp5_core_169;
  wire popcount27_qkp5_core_171;
  wire popcount27_qkp5_core_172;
  wire popcount27_qkp5_core_173;
  wire popcount27_qkp5_core_174_not;
  wire popcount27_qkp5_core_176;
  wire popcount27_qkp5_core_179;
  wire popcount27_qkp5_core_182;
  wire popcount27_qkp5_core_183;
  wire popcount27_qkp5_core_185;
  wire popcount27_qkp5_core_187;
  wire popcount27_qkp5_core_190;
  wire popcount27_qkp5_core_191;
  wire popcount27_qkp5_core_192;
  wire popcount27_qkp5_core_193;
  wire popcount27_qkp5_core_194;
  wire popcount27_qkp5_core_195;

  assign popcount27_qkp5_core_029 = ~input_a[20];
  assign popcount27_qkp5_core_030 = input_a[2] & input_a[7];
  assign popcount27_qkp5_core_032 = ~input_a[10];
  assign popcount27_qkp5_core_033 = input_a[11] & input_a[6];
  assign popcount27_qkp5_core_034 = ~input_a[21];
  assign popcount27_qkp5_core_035 = input_a[7] ^ input_a[14];
  assign popcount27_qkp5_core_036 = ~input_a[20];
  assign popcount27_qkp5_core_038 = input_a[18] ^ input_a[4];
  assign popcount27_qkp5_core_039 = ~(input_a[18] ^ input_a[25]);
  assign popcount27_qkp5_core_040 = ~(input_a[26] | input_a[19]);
  assign popcount27_qkp5_core_043 = input_a[9] ^ input_a[12];
  assign popcount27_qkp5_core_044 = ~input_a[2];
  assign popcount27_qkp5_core_045 = ~(input_a[20] | input_a[25]);
  assign popcount27_qkp5_core_048 = ~(input_a[15] | input_a[3]);
  assign popcount27_qkp5_core_049 = input_a[7] ^ input_a[21];
  assign popcount27_qkp5_core_050 = ~input_a[11];
  assign popcount27_qkp5_core_051 = ~input_a[14];
  assign popcount27_qkp5_core_052 = input_a[18] | input_a[9];
  assign popcount27_qkp5_core_053 = input_a[4] & input_a[3];
  assign popcount27_qkp5_core_054 = ~(input_a[0] | input_a[21]);
  assign popcount27_qkp5_core_055 = ~(input_a[23] & input_a[4]);
  assign popcount27_qkp5_core_057 = ~(input_a[22] ^ input_a[7]);
  assign popcount27_qkp5_core_059 = ~input_a[4];
  assign popcount27_qkp5_core_060 = ~(input_a[23] | input_a[9]);
  assign popcount27_qkp5_core_061 = ~(input_a[17] & input_a[8]);
  assign popcount27_qkp5_core_062 = ~(input_a[17] ^ input_a[21]);
  assign popcount27_qkp5_core_064 = ~(input_a[5] ^ input_a[21]);
  assign popcount27_qkp5_core_065 = ~(input_a[10] & input_a[7]);
  assign popcount27_qkp5_core_067 = ~(input_a[23] | input_a[20]);
  assign popcount27_qkp5_core_069 = input_a[26] | input_a[2];
  assign popcount27_qkp5_core_070 = input_a[14] & input_a[22];
  assign popcount27_qkp5_core_071 = input_a[6] & input_a[16];
  assign popcount27_qkp5_core_072 = input_a[24] | input_a[13];
  assign popcount27_qkp5_core_074 = input_a[16] & input_a[18];
  assign popcount27_qkp5_core_075 = input_a[25] | input_a[19];
  assign popcount27_qkp5_core_076 = ~(input_a[6] ^ input_a[4]);
  assign popcount27_qkp5_core_078 = input_a[4] & input_a[15];
  assign popcount27_qkp5_core_081 = input_a[7] ^ input_a[15];
  assign popcount27_qkp5_core_082 = input_a[19] ^ input_a[10];
  assign popcount27_qkp5_core_086 = ~(input_a[25] ^ input_a[24]);
  assign popcount27_qkp5_core_089 = input_a[15] ^ input_a[8];
  assign popcount27_qkp5_core_091 = input_a[9] & input_a[25];
  assign popcount27_qkp5_core_092 = ~input_a[23];
  assign popcount27_qkp5_core_093 = ~(input_a[26] | input_a[5]);
  assign popcount27_qkp5_core_096 = ~(input_a[15] & input_a[1]);
  assign popcount27_qkp5_core_097 = ~(input_a[21] & input_a[26]);
  assign popcount27_qkp5_core_098 = ~input_a[11];
  assign popcount27_qkp5_core_099 = ~(input_a[6] & input_a[12]);
  assign popcount27_qkp5_core_100 = ~input_a[24];
  assign popcount27_qkp5_core_102 = input_a[12] & input_a[18];
  assign popcount27_qkp5_core_104 = input_a[9] & input_a[2];
  assign popcount27_qkp5_core_105 = ~(input_a[13] ^ input_a[24]);
  assign popcount27_qkp5_core_108 = ~(input_a[19] & input_a[16]);
  assign popcount27_qkp5_core_110 = ~input_a[17];
  assign popcount27_qkp5_core_111 = input_a[14] | input_a[1];
  assign popcount27_qkp5_core_112 = input_a[1] ^ input_a[7];
  assign popcount27_qkp5_core_113 = ~(input_a[22] | input_a[16]);
  assign popcount27_qkp5_core_117 = ~(input_a[18] & input_a[3]);
  assign popcount27_qkp5_core_120 = ~(input_a[0] & input_a[21]);
  assign popcount27_qkp5_core_121 = ~(input_a[25] ^ input_a[23]);
  assign popcount27_qkp5_core_122 = ~(input_a[2] | input_a[1]);
  assign popcount27_qkp5_core_123 = input_a[0] | input_a[23];
  assign popcount27_qkp5_core_124 = ~input_a[16];
  assign popcount27_qkp5_core_127 = ~(input_a[14] ^ input_a[9]);
  assign popcount27_qkp5_core_129 = input_a[9] | input_a[5];
  assign popcount27_qkp5_core_131_not = ~input_a[16];
  assign popcount27_qkp5_core_132 = ~(input_a[22] ^ input_a[21]);
  assign popcount27_qkp5_core_134 = ~(input_a[7] | input_a[18]);
  assign popcount27_qkp5_core_138 = input_a[19] ^ input_a[25];
  assign popcount27_qkp5_core_139 = ~(input_a[9] & input_a[18]);
  assign popcount27_qkp5_core_142 = ~(input_a[7] ^ input_a[16]);
  assign popcount27_qkp5_core_143 = ~input_a[24];
  assign popcount27_qkp5_core_144 = ~input_a[20];
  assign popcount27_qkp5_core_145 = input_a[3] ^ input_a[24];
  assign popcount27_qkp5_core_148 = ~(input_a[16] | input_a[12]);
  assign popcount27_qkp5_core_149 = ~input_a[21];
  assign popcount27_qkp5_core_150 = ~input_a[5];
  assign popcount27_qkp5_core_152_not = ~input_a[20];
  assign popcount27_qkp5_core_153 = ~input_a[2];
  assign popcount27_qkp5_core_154 = input_a[15] | input_a[15];
  assign popcount27_qkp5_core_157 = input_a[9] ^ input_a[18];
  assign popcount27_qkp5_core_158 = ~(input_a[18] ^ input_a[11]);
  assign popcount27_qkp5_core_159 = input_a[22] ^ input_a[7];
  assign popcount27_qkp5_core_160 = input_a[11] | input_a[15];
  assign popcount27_qkp5_core_162 = ~input_a[22];
  assign popcount27_qkp5_core_163 = input_a[10] ^ input_a[21];
  assign popcount27_qkp5_core_166 = input_a[7] ^ input_a[24];
  assign popcount27_qkp5_core_167 = input_a[22] & input_a[26];
  assign popcount27_qkp5_core_168 = input_a[6] | input_a[26];
  assign popcount27_qkp5_core_169 = input_a[8] | input_a[6];
  assign popcount27_qkp5_core_171 = ~(input_a[21] & input_a[7]);
  assign popcount27_qkp5_core_172 = ~(input_a[1] | input_a[1]);
  assign popcount27_qkp5_core_173 = input_a[17] | input_a[4];
  assign popcount27_qkp5_core_174_not = ~input_a[9];
  assign popcount27_qkp5_core_176 = input_a[6] | input_a[7];
  assign popcount27_qkp5_core_179 = ~input_a[20];
  assign popcount27_qkp5_core_182 = ~(input_a[22] & input_a[12]);
  assign popcount27_qkp5_core_183 = ~(input_a[25] & input_a[20]);
  assign popcount27_qkp5_core_185 = input_a[11] | input_a[10];
  assign popcount27_qkp5_core_187 = input_a[8] & input_a[2];
  assign popcount27_qkp5_core_190 = ~input_a[25];
  assign popcount27_qkp5_core_191 = input_a[13] ^ input_a[3];
  assign popcount27_qkp5_core_192 = ~(input_a[3] | input_a[13]);
  assign popcount27_qkp5_core_193 = ~(input_a[1] ^ input_a[21]);
  assign popcount27_qkp5_core_194 = input_a[9] | input_a[16];
  assign popcount27_qkp5_core_195 = ~input_a[6];

  assign popcount27_qkp5_out[0] = 1'b1;
  assign popcount27_qkp5_out[1] = input_a[8];
  assign popcount27_qkp5_out[2] = input_a[14];
  assign popcount27_qkp5_out[3] = 1'b1;
  assign popcount27_qkp5_out[4] = 1'b0;
endmodule