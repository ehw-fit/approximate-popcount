// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.09504
// WCE=16.0
// EP=0.956163%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_avee(input [23:0] input_a, output [4:0] popcount24_avee_out);
  wire popcount24_avee_core_026;
  wire popcount24_avee_core_027;
  wire popcount24_avee_core_028;
  wire popcount24_avee_core_029;
  wire popcount24_avee_core_030;
  wire popcount24_avee_core_032;
  wire popcount24_avee_core_033;
  wire popcount24_avee_core_034;
  wire popcount24_avee_core_036;
  wire popcount24_avee_core_037;
  wire popcount24_avee_core_038;
  wire popcount24_avee_core_039;
  wire popcount24_avee_core_041_not;
  wire popcount24_avee_core_042_not;
  wire popcount24_avee_core_045;
  wire popcount24_avee_core_046;
  wire popcount24_avee_core_050;
  wire popcount24_avee_core_052;
  wire popcount24_avee_core_055;
  wire popcount24_avee_core_057;
  wire popcount24_avee_core_058;
  wire popcount24_avee_core_059;
  wire popcount24_avee_core_060;
  wire popcount24_avee_core_061;
  wire popcount24_avee_core_062;
  wire popcount24_avee_core_063;
  wire popcount24_avee_core_064;
  wire popcount24_avee_core_066;
  wire popcount24_avee_core_068;
  wire popcount24_avee_core_069;
  wire popcount24_avee_core_070;
  wire popcount24_avee_core_072;
  wire popcount24_avee_core_073;
  wire popcount24_avee_core_074;
  wire popcount24_avee_core_075_not;
  wire popcount24_avee_core_076;
  wire popcount24_avee_core_078;
  wire popcount24_avee_core_079;
  wire popcount24_avee_core_080;
  wire popcount24_avee_core_081;
  wire popcount24_avee_core_082;
  wire popcount24_avee_core_084;
  wire popcount24_avee_core_085;
  wire popcount24_avee_core_087;
  wire popcount24_avee_core_088;
  wire popcount24_avee_core_092;
  wire popcount24_avee_core_093;
  wire popcount24_avee_core_094;
  wire popcount24_avee_core_095;
  wire popcount24_avee_core_096;
  wire popcount24_avee_core_098;
  wire popcount24_avee_core_100;
  wire popcount24_avee_core_101;
  wire popcount24_avee_core_104;
  wire popcount24_avee_core_106;
  wire popcount24_avee_core_107;
  wire popcount24_avee_core_108;
  wire popcount24_avee_core_111;
  wire popcount24_avee_core_112;
  wire popcount24_avee_core_113;
  wire popcount24_avee_core_114;
  wire popcount24_avee_core_116;
  wire popcount24_avee_core_117;
  wire popcount24_avee_core_118;
  wire popcount24_avee_core_119;
  wire popcount24_avee_core_120;
  wire popcount24_avee_core_122;
  wire popcount24_avee_core_123;
  wire popcount24_avee_core_124;
  wire popcount24_avee_core_126;
  wire popcount24_avee_core_127;
  wire popcount24_avee_core_128;
  wire popcount24_avee_core_129;
  wire popcount24_avee_core_130;
  wire popcount24_avee_core_131_not;
  wire popcount24_avee_core_132;
  wire popcount24_avee_core_133;
  wire popcount24_avee_core_135;
  wire popcount24_avee_core_137;
  wire popcount24_avee_core_139;
  wire popcount24_avee_core_140;
  wire popcount24_avee_core_141;
  wire popcount24_avee_core_143;
  wire popcount24_avee_core_145;
  wire popcount24_avee_core_146;
  wire popcount24_avee_core_148;
  wire popcount24_avee_core_150;
  wire popcount24_avee_core_152;
  wire popcount24_avee_core_153;
  wire popcount24_avee_core_154;
  wire popcount24_avee_core_157;
  wire popcount24_avee_core_158;
  wire popcount24_avee_core_159;
  wire popcount24_avee_core_161;
  wire popcount24_avee_core_162;
  wire popcount24_avee_core_164;
  wire popcount24_avee_core_165;
  wire popcount24_avee_core_166;
  wire popcount24_avee_core_167;
  wire popcount24_avee_core_168;
  wire popcount24_avee_core_169;
  wire popcount24_avee_core_173;
  wire popcount24_avee_core_174;
  wire popcount24_avee_core_175;
  wire popcount24_avee_core_176;

  assign popcount24_avee_core_026 = ~(input_a[5] & input_a[23]);
  assign popcount24_avee_core_027 = ~input_a[1];
  assign popcount24_avee_core_028 = input_a[17] ^ input_a[1];
  assign popcount24_avee_core_029 = input_a[8] | input_a[8];
  assign popcount24_avee_core_030 = ~(input_a[1] ^ input_a[16]);
  assign popcount24_avee_core_032 = input_a[12] | input_a[11];
  assign popcount24_avee_core_033 = input_a[12] | input_a[8];
  assign popcount24_avee_core_034 = ~input_a[23];
  assign popcount24_avee_core_036 = input_a[13] ^ input_a[1];
  assign popcount24_avee_core_037 = ~(input_a[9] | input_a[12]);
  assign popcount24_avee_core_038 = ~(input_a[5] ^ input_a[20]);
  assign popcount24_avee_core_039 = input_a[11] & input_a[15];
  assign popcount24_avee_core_041_not = ~input_a[2];
  assign popcount24_avee_core_042_not = ~input_a[5];
  assign popcount24_avee_core_045 = ~(input_a[9] | input_a[8]);
  assign popcount24_avee_core_046 = input_a[11] ^ input_a[1];
  assign popcount24_avee_core_050 = ~(input_a[4] | input_a[3]);
  assign popcount24_avee_core_052 = input_a[9] ^ input_a[8];
  assign popcount24_avee_core_055 = input_a[18] | input_a[5];
  assign popcount24_avee_core_057 = ~(input_a[16] ^ input_a[7]);
  assign popcount24_avee_core_058 = ~(input_a[6] & input_a[23]);
  assign popcount24_avee_core_059 = input_a[16] ^ input_a[2];
  assign popcount24_avee_core_060 = input_a[19] ^ input_a[21];
  assign popcount24_avee_core_061 = ~input_a[14];
  assign popcount24_avee_core_062 = input_a[9] & input_a[4];
  assign popcount24_avee_core_063 = ~(input_a[2] | input_a[0]);
  assign popcount24_avee_core_064 = ~(input_a[13] | input_a[22]);
  assign popcount24_avee_core_066 = ~(input_a[14] & input_a[15]);
  assign popcount24_avee_core_068 = input_a[2] | input_a[15];
  assign popcount24_avee_core_069 = input_a[11] & input_a[15];
  assign popcount24_avee_core_070 = input_a[2] ^ input_a[11];
  assign popcount24_avee_core_072 = ~input_a[23];
  assign popcount24_avee_core_073 = input_a[13] ^ input_a[2];
  assign popcount24_avee_core_074 = ~(input_a[7] ^ input_a[9]);
  assign popcount24_avee_core_075_not = ~input_a[3];
  assign popcount24_avee_core_076 = ~(input_a[9] | input_a[14]);
  assign popcount24_avee_core_078 = input_a[9] | input_a[14];
  assign popcount24_avee_core_079 = input_a[23] ^ input_a[14];
  assign popcount24_avee_core_080 = ~(input_a[20] | input_a[19]);
  assign popcount24_avee_core_081 = ~input_a[2];
  assign popcount24_avee_core_082 = ~(input_a[4] ^ input_a[1]);
  assign popcount24_avee_core_084 = ~(input_a[9] | input_a[12]);
  assign popcount24_avee_core_085 = input_a[13] | input_a[1];
  assign popcount24_avee_core_087 = input_a[23] & input_a[3];
  assign popcount24_avee_core_088 = ~input_a[18];
  assign popcount24_avee_core_092 = ~(input_a[21] & input_a[6]);
  assign popcount24_avee_core_093 = ~(input_a[1] ^ input_a[12]);
  assign popcount24_avee_core_094 = ~(input_a[7] & input_a[23]);
  assign popcount24_avee_core_095 = input_a[17] | input_a[19];
  assign popcount24_avee_core_096 = ~(input_a[17] | input_a[0]);
  assign popcount24_avee_core_098 = ~(input_a[1] & input_a[18]);
  assign popcount24_avee_core_100 = ~(input_a[1] ^ input_a[4]);
  assign popcount24_avee_core_101 = ~(input_a[12] ^ input_a[9]);
  assign popcount24_avee_core_104 = input_a[22] | input_a[16];
  assign popcount24_avee_core_106 = input_a[14] ^ input_a[13];
  assign popcount24_avee_core_107 = input_a[17] | input_a[5];
  assign popcount24_avee_core_108 = input_a[14] & input_a[9];
  assign popcount24_avee_core_111 = ~(input_a[13] ^ input_a[21]);
  assign popcount24_avee_core_112 = input_a[14] ^ input_a[19];
  assign popcount24_avee_core_113 = input_a[0] & input_a[20];
  assign popcount24_avee_core_114 = ~(input_a[8] ^ input_a[12]);
  assign popcount24_avee_core_116 = ~(input_a[13] ^ input_a[2]);
  assign popcount24_avee_core_117 = input_a[16] ^ input_a[21];
  assign popcount24_avee_core_118 = input_a[2] ^ input_a[7];
  assign popcount24_avee_core_119 = input_a[4] & input_a[10];
  assign popcount24_avee_core_120 = input_a[8] ^ input_a[15];
  assign popcount24_avee_core_122 = ~(input_a[15] | input_a[22]);
  assign popcount24_avee_core_123 = ~(input_a[8] | input_a[16]);
  assign popcount24_avee_core_124 = input_a[19] ^ input_a[9];
  assign popcount24_avee_core_126 = ~(input_a[19] | input_a[15]);
  assign popcount24_avee_core_127 = ~(input_a[8] | input_a[7]);
  assign popcount24_avee_core_128 = input_a[8] & input_a[6];
  assign popcount24_avee_core_129 = ~input_a[14];
  assign popcount24_avee_core_130 = input_a[7] | input_a[16];
  assign popcount24_avee_core_131_not = ~input_a[20];
  assign popcount24_avee_core_132 = ~(input_a[12] ^ input_a[16]);
  assign popcount24_avee_core_133 = ~(input_a[23] ^ input_a[19]);
  assign popcount24_avee_core_135 = ~(input_a[13] & input_a[22]);
  assign popcount24_avee_core_137 = ~(input_a[16] & input_a[13]);
  assign popcount24_avee_core_139 = input_a[20] | input_a[11];
  assign popcount24_avee_core_140 = ~(input_a[21] | input_a[9]);
  assign popcount24_avee_core_141 = input_a[9] ^ input_a[15];
  assign popcount24_avee_core_143 = input_a[17] & input_a[2];
  assign popcount24_avee_core_145 = input_a[23] ^ input_a[21];
  assign popcount24_avee_core_146 = ~(input_a[14] ^ input_a[9]);
  assign popcount24_avee_core_148 = ~(input_a[6] & input_a[22]);
  assign popcount24_avee_core_150 = input_a[14] & input_a[2];
  assign popcount24_avee_core_152 = ~(input_a[7] & input_a[15]);
  assign popcount24_avee_core_153 = ~(input_a[16] ^ input_a[18]);
  assign popcount24_avee_core_154 = ~(input_a[22] & input_a[19]);
  assign popcount24_avee_core_157 = input_a[17] | input_a[13];
  assign popcount24_avee_core_158 = ~(input_a[2] | input_a[14]);
  assign popcount24_avee_core_159 = input_a[7] ^ input_a[11];
  assign popcount24_avee_core_161 = ~input_a[23];
  assign popcount24_avee_core_162 = ~(input_a[5] & input_a[0]);
  assign popcount24_avee_core_164 = ~(input_a[6] | input_a[23]);
  assign popcount24_avee_core_165 = input_a[15] | input_a[12];
  assign popcount24_avee_core_166 = ~input_a[4];
  assign popcount24_avee_core_167 = ~input_a[13];
  assign popcount24_avee_core_168 = ~input_a[21];
  assign popcount24_avee_core_169 = ~(input_a[4] | input_a[3]);
  assign popcount24_avee_core_173 = ~(input_a[12] ^ input_a[16]);
  assign popcount24_avee_core_174 = input_a[20] & input_a[15];
  assign popcount24_avee_core_175 = ~(input_a[7] & input_a[5]);
  assign popcount24_avee_core_176 = ~input_a[13];

  assign popcount24_avee_out[0] = 1'b0;
  assign popcount24_avee_out[1] = 1'b0;
  assign popcount24_avee_out[2] = 1'b0;
  assign popcount24_avee_out[3] = 1'b1;
  assign popcount24_avee_out[4] = 1'b0;
endmodule