// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.55958
// WCE=10.0
// EP=0.894341%
// Printed PDK parameters:
//  Area=5993720.0
//  Delay=14305946.0
//  Power=261280.0

module popcount19_w96b(input [18:0] input_a, output [4:0] popcount19_w96b_out);
  wire popcount19_w96b_core_021;
  wire popcount19_w96b_core_022;
  wire popcount19_w96b_core_023;
  wire popcount19_w96b_core_025;
  wire popcount19_w96b_core_028;
  wire popcount19_w96b_core_029_not;
  wire popcount19_w96b_core_033;
  wire popcount19_w96b_core_035;
  wire popcount19_w96b_core_036;
  wire popcount19_w96b_core_037;
  wire popcount19_w96b_core_041;
  wire popcount19_w96b_core_044;
  wire popcount19_w96b_core_046;
  wire popcount19_w96b_core_047;
  wire popcount19_w96b_core_048;
  wire popcount19_w96b_core_049;
  wire popcount19_w96b_core_051;
  wire popcount19_w96b_core_052;
  wire popcount19_w96b_core_053;
  wire popcount19_w96b_core_055;
  wire popcount19_w96b_core_057;
  wire popcount19_w96b_core_058;
  wire popcount19_w96b_core_059;
  wire popcount19_w96b_core_061;
  wire popcount19_w96b_core_062;
  wire popcount19_w96b_core_063;
  wire popcount19_w96b_core_067;
  wire popcount19_w96b_core_069;
  wire popcount19_w96b_core_070;
  wire popcount19_w96b_core_071;
  wire popcount19_w96b_core_073;
  wire popcount19_w96b_core_074;
  wire popcount19_w96b_core_075;
  wire popcount19_w96b_core_076;
  wire popcount19_w96b_core_078;
  wire popcount19_w96b_core_079;
  wire popcount19_w96b_core_081;
  wire popcount19_w96b_core_082;
  wire popcount19_w96b_core_083;
  wire popcount19_w96b_core_084;
  wire popcount19_w96b_core_085;
  wire popcount19_w96b_core_086;
  wire popcount19_w96b_core_087;
  wire popcount19_w96b_core_089;
  wire popcount19_w96b_core_090;
  wire popcount19_w96b_core_091;
  wire popcount19_w96b_core_092;
  wire popcount19_w96b_core_093;
  wire popcount19_w96b_core_095;
  wire popcount19_w96b_core_096;
  wire popcount19_w96b_core_097;
  wire popcount19_w96b_core_099;
  wire popcount19_w96b_core_100;
  wire popcount19_w96b_core_102;
  wire popcount19_w96b_core_106;
  wire popcount19_w96b_core_107;
  wire popcount19_w96b_core_108;
  wire popcount19_w96b_core_110;
  wire popcount19_w96b_core_111;
  wire popcount19_w96b_core_113;
  wire popcount19_w96b_core_114;
  wire popcount19_w96b_core_116;
  wire popcount19_w96b_core_117;
  wire popcount19_w96b_core_118;
  wire popcount19_w96b_core_121;
  wire popcount19_w96b_core_122;
  wire popcount19_w96b_core_123;
  wire popcount19_w96b_core_126;
  wire popcount19_w96b_core_128;
  wire popcount19_w96b_core_131;
  wire popcount19_w96b_core_132;
  wire popcount19_w96b_core_133;

  assign popcount19_w96b_core_021 = input_a[4] | input_a[11];
  assign popcount19_w96b_core_022 = input_a[15] & input_a[18];
  assign popcount19_w96b_core_023 = input_a[17] ^ input_a[8];
  assign popcount19_w96b_core_025 = ~(input_a[10] | input_a[1]);
  assign popcount19_w96b_core_028 = input_a[9] | input_a[11];
  assign popcount19_w96b_core_029_not = ~input_a[18];
  assign popcount19_w96b_core_033 = ~input_a[10];
  assign popcount19_w96b_core_035 = ~(input_a[10] & input_a[12]);
  assign popcount19_w96b_core_036 = input_a[4] & input_a[9];
  assign popcount19_w96b_core_037 = input_a[4] ^ input_a[2];
  assign popcount19_w96b_core_041 = ~(input_a[11] ^ input_a[15]);
  assign popcount19_w96b_core_044 = ~(input_a[13] & input_a[16]);
  assign popcount19_w96b_core_046 = ~(input_a[9] | input_a[14]);
  assign popcount19_w96b_core_047 = ~(input_a[8] & input_a[7]);
  assign popcount19_w96b_core_048 = ~(input_a[17] & input_a[13]);
  assign popcount19_w96b_core_049 = ~input_a[18];
  assign popcount19_w96b_core_051 = ~input_a[9];
  assign popcount19_w96b_core_052 = ~(input_a[18] | input_a[8]);
  assign popcount19_w96b_core_053 = input_a[10] | input_a[11];
  assign popcount19_w96b_core_055 = input_a[7] | input_a[0];
  assign popcount19_w96b_core_057 = input_a[9] | input_a[7];
  assign popcount19_w96b_core_058 = input_a[1] | popcount19_w96b_core_055;
  assign popcount19_w96b_core_059 = input_a[2] | input_a[15];
  assign popcount19_w96b_core_061 = input_a[16] ^ input_a[7];
  assign popcount19_w96b_core_062 = input_a[15] ^ input_a[10];
  assign popcount19_w96b_core_063 = input_a[16] & input_a[17];
  assign popcount19_w96b_core_067 = input_a[9] | input_a[17];
  assign popcount19_w96b_core_069 = ~input_a[8];
  assign popcount19_w96b_core_070 = input_a[17] ^ input_a[2];
  assign popcount19_w96b_core_071 = ~input_a[0];
  assign popcount19_w96b_core_073 = input_a[9] & input_a[14];
  assign popcount19_w96b_core_074 = ~(input_a[5] ^ input_a[15]);
  assign popcount19_w96b_core_075 = ~(input_a[12] & input_a[13]);
  assign popcount19_w96b_core_076 = input_a[0] & input_a[5];
  assign popcount19_w96b_core_078 = ~(input_a[11] | input_a[15]);
  assign popcount19_w96b_core_079 = input_a[2] | input_a[17];
  assign popcount19_w96b_core_081 = ~input_a[17];
  assign popcount19_w96b_core_082 = input_a[12] ^ input_a[4];
  assign popcount19_w96b_core_083 = ~(input_a[7] & input_a[17]);
  assign popcount19_w96b_core_084 = ~input_a[17];
  assign popcount19_w96b_core_085 = input_a[5] | input_a[16];
  assign popcount19_w96b_core_086 = ~input_a[18];
  assign popcount19_w96b_core_087 = ~(input_a[16] ^ input_a[18]);
  assign popcount19_w96b_core_089 = input_a[10] ^ input_a[18];
  assign popcount19_w96b_core_090 = ~input_a[18];
  assign popcount19_w96b_core_091 = input_a[13] & input_a[18];
  assign popcount19_w96b_core_092 = input_a[17] | input_a[11];
  assign popcount19_w96b_core_093 = input_a[1] ^ input_a[7];
  assign popcount19_w96b_core_095 = input_a[12] | input_a[14];
  assign popcount19_w96b_core_096 = ~(input_a[9] | input_a[7]);
  assign popcount19_w96b_core_097 = input_a[1] & input_a[3];
  assign popcount19_w96b_core_099 = ~(input_a[6] & popcount19_w96b_core_092);
  assign popcount19_w96b_core_100 = input_a[6] & popcount19_w96b_core_092;
  assign popcount19_w96b_core_102 = ~(input_a[10] & input_a[11]);
  assign popcount19_w96b_core_106 = ~input_a[6];
  assign popcount19_w96b_core_107 = input_a[6] & popcount19_w96b_core_100;
  assign popcount19_w96b_core_108 = input_a[2] | popcount19_w96b_core_107;
  assign popcount19_w96b_core_110 = ~input_a[4];
  assign popcount19_w96b_core_111 = input_a[2] | popcount19_w96b_core_108;
  assign popcount19_w96b_core_113 = input_a[14] | input_a[13];
  assign popcount19_w96b_core_114 = input_a[7] | input_a[12];
  assign popcount19_w96b_core_116 = input_a[2] ^ popcount19_w96b_core_099;
  assign popcount19_w96b_core_117 = input_a[2] & popcount19_w96b_core_099;
  assign popcount19_w96b_core_118 = ~(input_a[3] ^ input_a[14]);
  assign popcount19_w96b_core_121 = popcount19_w96b_core_058 ^ popcount19_w96b_core_106;
  assign popcount19_w96b_core_122 = popcount19_w96b_core_058 & popcount19_w96b_core_106;
  assign popcount19_w96b_core_123 = popcount19_w96b_core_121 ^ popcount19_w96b_core_117;
  assign popcount19_w96b_core_126 = input_a[2] | popcount19_w96b_core_111;
  assign popcount19_w96b_core_128 = popcount19_w96b_core_126 | popcount19_w96b_core_122;
  assign popcount19_w96b_core_131 = ~(input_a[14] | input_a[7]);
  assign popcount19_w96b_core_132 = ~(input_a[11] ^ input_a[4]);
  assign popcount19_w96b_core_133 = input_a[5] ^ input_a[14];

  assign popcount19_w96b_out[0] = input_a[8];
  assign popcount19_w96b_out[1] = popcount19_w96b_core_116;
  assign popcount19_w96b_out[2] = popcount19_w96b_core_123;
  assign popcount19_w96b_out[3] = popcount19_w96b_core_128;
  assign popcount19_w96b_out[4] = 1'b0;
endmodule