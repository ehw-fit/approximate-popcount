// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.37915
// WCE=17.0
// EP=0.868282%
// Printed PDK parameters:
//  Area=1123640.0
//  Delay=4181376.75
//  Power=39342.0

module popcount34_28tv(input [33:0] input_a, output [5:0] popcount34_28tv_out);
  wire popcount34_28tv_core_036;
  wire popcount34_28tv_core_040_not;
  wire popcount34_28tv_core_041;
  wire popcount34_28tv_core_042;
  wire popcount34_28tv_core_044;
  wire popcount34_28tv_core_052;
  wire popcount34_28tv_core_053;
  wire popcount34_28tv_core_054;
  wire popcount34_28tv_core_055;
  wire popcount34_28tv_core_056;
  wire popcount34_28tv_core_058;
  wire popcount34_28tv_core_059;
  wire popcount34_28tv_core_062;
  wire popcount34_28tv_core_063;
  wire popcount34_28tv_core_065;
  wire popcount34_28tv_core_067;
  wire popcount34_28tv_core_068;
  wire popcount34_28tv_core_069;
  wire popcount34_28tv_core_070;
  wire popcount34_28tv_core_071;
  wire popcount34_28tv_core_073;
  wire popcount34_28tv_core_075;
  wire popcount34_28tv_core_076;
  wire popcount34_28tv_core_077;
  wire popcount34_28tv_core_078;
  wire popcount34_28tv_core_080;
  wire popcount34_28tv_core_083_not;
  wire popcount34_28tv_core_085;
  wire popcount34_28tv_core_086;
  wire popcount34_28tv_core_087;
  wire popcount34_28tv_core_088;
  wire popcount34_28tv_core_089;
  wire popcount34_28tv_core_092;
  wire popcount34_28tv_core_093;
  wire popcount34_28tv_core_094;
  wire popcount34_28tv_core_099;
  wire popcount34_28tv_core_101;
  wire popcount34_28tv_core_103;
  wire popcount34_28tv_core_104;
  wire popcount34_28tv_core_105;
  wire popcount34_28tv_core_107;
  wire popcount34_28tv_core_108;
  wire popcount34_28tv_core_115;
  wire popcount34_28tv_core_116;
  wire popcount34_28tv_core_118;
  wire popcount34_28tv_core_119;
  wire popcount34_28tv_core_120_not;
  wire popcount34_28tv_core_121;
  wire popcount34_28tv_core_122;
  wire popcount34_28tv_core_124;
  wire popcount34_28tv_core_126;
  wire popcount34_28tv_core_128;
  wire popcount34_28tv_core_129;
  wire popcount34_28tv_core_131;
  wire popcount34_28tv_core_132;
  wire popcount34_28tv_core_133;
  wire popcount34_28tv_core_134;
  wire popcount34_28tv_core_135;
  wire popcount34_28tv_core_137;
  wire popcount34_28tv_core_138;
  wire popcount34_28tv_core_139;
  wire popcount34_28tv_core_142;
  wire popcount34_28tv_core_143;
  wire popcount34_28tv_core_144;
  wire popcount34_28tv_core_145;
  wire popcount34_28tv_core_146;
  wire popcount34_28tv_core_147;
  wire popcount34_28tv_core_148;
  wire popcount34_28tv_core_149;
  wire popcount34_28tv_core_150;
  wire popcount34_28tv_core_151;
  wire popcount34_28tv_core_154;
  wire popcount34_28tv_core_156;
  wire popcount34_28tv_core_157;
  wire popcount34_28tv_core_159;
  wire popcount34_28tv_core_162;
  wire popcount34_28tv_core_164;
  wire popcount34_28tv_core_166;
  wire popcount34_28tv_core_168;
  wire popcount34_28tv_core_169;
  wire popcount34_28tv_core_170;
  wire popcount34_28tv_core_172;
  wire popcount34_28tv_core_175;
  wire popcount34_28tv_core_176;
  wire popcount34_28tv_core_177;
  wire popcount34_28tv_core_178;
  wire popcount34_28tv_core_179;
  wire popcount34_28tv_core_181;
  wire popcount34_28tv_core_183;
  wire popcount34_28tv_core_185;
  wire popcount34_28tv_core_186;
  wire popcount34_28tv_core_187;
  wire popcount34_28tv_core_188;
  wire popcount34_28tv_core_189;
  wire popcount34_28tv_core_190;
  wire popcount34_28tv_core_193;
  wire popcount34_28tv_core_195;
  wire popcount34_28tv_core_196;
  wire popcount34_28tv_core_198;
  wire popcount34_28tv_core_199_not;
  wire popcount34_28tv_core_201;
  wire popcount34_28tv_core_204;
  wire popcount34_28tv_core_205;
  wire popcount34_28tv_core_207;
  wire popcount34_28tv_core_208;
  wire popcount34_28tv_core_209;
  wire popcount34_28tv_core_210;
  wire popcount34_28tv_core_211;
  wire popcount34_28tv_core_213;
  wire popcount34_28tv_core_216;
  wire popcount34_28tv_core_220;
  wire popcount34_28tv_core_221;
  wire popcount34_28tv_core_222;
  wire popcount34_28tv_core_223;
  wire popcount34_28tv_core_225;
  wire popcount34_28tv_core_226;
  wire popcount34_28tv_core_227;
  wire popcount34_28tv_core_230;
  wire popcount34_28tv_core_235;
  wire popcount34_28tv_core_236;
  wire popcount34_28tv_core_238;
  wire popcount34_28tv_core_240;
  wire popcount34_28tv_core_241;
  wire popcount34_28tv_core_242;
  wire popcount34_28tv_core_243;
  wire popcount34_28tv_core_244;
  wire popcount34_28tv_core_245;
  wire popcount34_28tv_core_246;
  wire popcount34_28tv_core_249;
  wire popcount34_28tv_core_250;
  wire popcount34_28tv_core_251_not;
  wire popcount34_28tv_core_252;

  assign popcount34_28tv_core_036 = ~(input_a[11] & input_a[11]);
  assign popcount34_28tv_core_040_not = ~input_a[11];
  assign popcount34_28tv_core_041 = ~(input_a[11] | input_a[6]);
  assign popcount34_28tv_core_042 = input_a[18] & input_a[18];
  assign popcount34_28tv_core_044 = input_a[25] | input_a[27];
  assign popcount34_28tv_core_052 = ~(input_a[8] & input_a[19]);
  assign popcount34_28tv_core_053 = input_a[29] | input_a[12];
  assign popcount34_28tv_core_054 = ~(input_a[33] | input_a[20]);
  assign popcount34_28tv_core_055 = input_a[7] ^ input_a[19];
  assign popcount34_28tv_core_056 = ~(input_a[14] & input_a[26]);
  assign popcount34_28tv_core_058 = input_a[13] | input_a[33];
  assign popcount34_28tv_core_059 = input_a[0] | input_a[17];
  assign popcount34_28tv_core_062 = input_a[19] | input_a[16];
  assign popcount34_28tv_core_063 = input_a[26] ^ input_a[18];
  assign popcount34_28tv_core_065 = ~input_a[12];
  assign popcount34_28tv_core_067 = input_a[18] | input_a[26];
  assign popcount34_28tv_core_068 = ~(input_a[22] & input_a[10]);
  assign popcount34_28tv_core_069 = ~input_a[29];
  assign popcount34_28tv_core_070 = input_a[2] | input_a[18];
  assign popcount34_28tv_core_071 = ~(input_a[12] | input_a[15]);
  assign popcount34_28tv_core_073 = ~input_a[15];
  assign popcount34_28tv_core_075 = ~(input_a[10] & input_a[3]);
  assign popcount34_28tv_core_076 = ~(input_a[18] & input_a[18]);
  assign popcount34_28tv_core_077 = input_a[5] ^ input_a[14];
  assign popcount34_28tv_core_078 = ~(input_a[28] | input_a[28]);
  assign popcount34_28tv_core_080 = ~(input_a[6] & input_a[17]);
  assign popcount34_28tv_core_083_not = ~input_a[27];
  assign popcount34_28tv_core_085 = ~(input_a[23] ^ input_a[21]);
  assign popcount34_28tv_core_086 = ~(input_a[22] & input_a[6]);
  assign popcount34_28tv_core_087 = ~(input_a[33] | input_a[4]);
  assign popcount34_28tv_core_088 = ~(input_a[29] | input_a[10]);
  assign popcount34_28tv_core_089 = input_a[33] & input_a[33];
  assign popcount34_28tv_core_092 = ~(input_a[23] | input_a[19]);
  assign popcount34_28tv_core_093 = input_a[10] | input_a[6];
  assign popcount34_28tv_core_094 = ~input_a[20];
  assign popcount34_28tv_core_099 = ~input_a[15];
  assign popcount34_28tv_core_101 = input_a[33] & input_a[15];
  assign popcount34_28tv_core_103 = ~input_a[9];
  assign popcount34_28tv_core_104 = input_a[8] | input_a[4];
  assign popcount34_28tv_core_105 = ~(input_a[7] | input_a[13]);
  assign popcount34_28tv_core_107 = ~(input_a[29] | input_a[23]);
  assign popcount34_28tv_core_108 = input_a[9] | input_a[18];
  assign popcount34_28tv_core_115 = ~(input_a[18] | input_a[2]);
  assign popcount34_28tv_core_116 = input_a[21] & input_a[3];
  assign popcount34_28tv_core_118 = ~(input_a[11] | input_a[13]);
  assign popcount34_28tv_core_119 = input_a[12] | input_a[1];
  assign popcount34_28tv_core_120_not = ~input_a[1];
  assign popcount34_28tv_core_121 = ~popcount34_28tv_core_119;
  assign popcount34_28tv_core_122 = input_a[32] ^ input_a[21];
  assign popcount34_28tv_core_124 = input_a[12] & input_a[27];
  assign popcount34_28tv_core_126 = input_a[12] | input_a[1];
  assign popcount34_28tv_core_128 = input_a[25] & input_a[8];
  assign popcount34_28tv_core_129 = input_a[20] ^ input_a[32];
  assign popcount34_28tv_core_131 = input_a[8] ^ input_a[13];
  assign popcount34_28tv_core_132 = input_a[13] ^ input_a[18];
  assign popcount34_28tv_core_133 = input_a[33] & input_a[22];
  assign popcount34_28tv_core_134 = input_a[33] & input_a[11];
  assign popcount34_28tv_core_135 = input_a[20] & input_a[24];
  assign popcount34_28tv_core_137 = ~(input_a[22] & input_a[25]);
  assign popcount34_28tv_core_138 = input_a[26] | input_a[23];
  assign popcount34_28tv_core_139 = ~(input_a[10] & input_a[8]);
  assign popcount34_28tv_core_142 = input_a[7] | input_a[21];
  assign popcount34_28tv_core_143 = ~(input_a[11] | input_a[9]);
  assign popcount34_28tv_core_144 = ~(input_a[28] & input_a[25]);
  assign popcount34_28tv_core_145 = input_a[29] ^ input_a[23];
  assign popcount34_28tv_core_146 = ~input_a[33];
  assign popcount34_28tv_core_147 = ~(input_a[16] | input_a[4]);
  assign popcount34_28tv_core_148 = ~(input_a[32] | input_a[3]);
  assign popcount34_28tv_core_149 = input_a[17] & input_a[15];
  assign popcount34_28tv_core_150 = ~input_a[13];
  assign popcount34_28tv_core_151 = ~(input_a[2] ^ input_a[11]);
  assign popcount34_28tv_core_154 = input_a[29] ^ input_a[24];
  assign popcount34_28tv_core_156 = input_a[18] ^ input_a[1];
  assign popcount34_28tv_core_157 = input_a[20] | input_a[4];
  assign popcount34_28tv_core_159 = input_a[7] & input_a[13];
  assign popcount34_28tv_core_162 = ~(input_a[1] & input_a[23]);
  assign popcount34_28tv_core_164 = input_a[24] | input_a[17];
  assign popcount34_28tv_core_166 = ~(input_a[18] | input_a[18]);
  assign popcount34_28tv_core_168 = ~(input_a[23] ^ input_a[19]);
  assign popcount34_28tv_core_169 = ~(input_a[8] | input_a[11]);
  assign popcount34_28tv_core_170 = ~input_a[10];
  assign popcount34_28tv_core_172 = input_a[13] | input_a[23];
  assign popcount34_28tv_core_175 = ~(input_a[21] | input_a[10]);
  assign popcount34_28tv_core_176 = ~(input_a[27] & input_a[12]);
  assign popcount34_28tv_core_177 = input_a[1] ^ input_a[14];
  assign popcount34_28tv_core_178 = ~input_a[13];
  assign popcount34_28tv_core_179 = ~(input_a[31] ^ input_a[9]);
  assign popcount34_28tv_core_181 = ~(input_a[6] ^ input_a[32]);
  assign popcount34_28tv_core_183 = ~(input_a[0] | input_a[14]);
  assign popcount34_28tv_core_185 = input_a[7] ^ input_a[32];
  assign popcount34_28tv_core_186 = input_a[29] & input_a[13];
  assign popcount34_28tv_core_187 = input_a[11] | input_a[31];
  assign popcount34_28tv_core_188 = ~(input_a[2] & input_a[7]);
  assign popcount34_28tv_core_189 = ~(input_a[27] ^ input_a[30]);
  assign popcount34_28tv_core_190 = ~(input_a[15] ^ input_a[1]);
  assign popcount34_28tv_core_193 = ~(input_a[10] ^ input_a[19]);
  assign popcount34_28tv_core_195 = ~(input_a[21] & input_a[3]);
  assign popcount34_28tv_core_196 = input_a[4] | input_a[21];
  assign popcount34_28tv_core_198 = ~input_a[5];
  assign popcount34_28tv_core_199_not = ~input_a[2];
  assign popcount34_28tv_core_201 = ~input_a[24];
  assign popcount34_28tv_core_204 = ~(input_a[32] ^ input_a[15]);
  assign popcount34_28tv_core_205 = input_a[6] | input_a[15];
  assign popcount34_28tv_core_207 = ~(input_a[7] & input_a[14]);
  assign popcount34_28tv_core_208 = ~input_a[5];
  assign popcount34_28tv_core_209 = ~input_a[27];
  assign popcount34_28tv_core_210 = ~input_a[6];
  assign popcount34_28tv_core_211 = ~(input_a[12] | input_a[17]);
  assign popcount34_28tv_core_213 = ~input_a[19];
  assign popcount34_28tv_core_216 = ~(input_a[30] & input_a[19]);
  assign popcount34_28tv_core_220 = ~(input_a[11] | input_a[6]);
  assign popcount34_28tv_core_221 = ~input_a[9];
  assign popcount34_28tv_core_222 = input_a[5] | input_a[31];
  assign popcount34_28tv_core_223 = ~input_a[16];
  assign popcount34_28tv_core_225 = ~(input_a[29] & input_a[4]);
  assign popcount34_28tv_core_226 = ~(input_a[17] | input_a[30]);
  assign popcount34_28tv_core_227 = input_a[17] | input_a[1];
  assign popcount34_28tv_core_230 = ~(input_a[19] & input_a[32]);
  assign popcount34_28tv_core_235 = ~input_a[11];
  assign popcount34_28tv_core_236 = popcount34_28tv_core_121 & popcount34_28tv_core_116;
  assign popcount34_28tv_core_238 = ~popcount34_28tv_core_126;
  assign popcount34_28tv_core_240 = popcount34_28tv_core_238 ^ popcount34_28tv_core_236;
  assign popcount34_28tv_core_241 = input_a[21] & input_a[3];
  assign popcount34_28tv_core_242 = popcount34_28tv_core_126 | popcount34_28tv_core_241;
  assign popcount34_28tv_core_243 = input_a[8] | input_a[2];
  assign popcount34_28tv_core_244 = ~(input_a[20] & input_a[19]);
  assign popcount34_28tv_core_245 = ~input_a[6];
  assign popcount34_28tv_core_246 = ~input_a[20];
  assign popcount34_28tv_core_249 = input_a[30] ^ input_a[9];
  assign popcount34_28tv_core_250 = input_a[24] & input_a[8];
  assign popcount34_28tv_core_251_not = ~input_a[25];
  assign popcount34_28tv_core_252 = ~(input_a[31] | input_a[22]);

  assign popcount34_28tv_out[0] = input_a[21];
  assign popcount34_28tv_out[1] = popcount34_28tv_core_238;
  assign popcount34_28tv_out[2] = popcount34_28tv_core_240;
  assign popcount34_28tv_out[3] = popcount34_28tv_core_240;
  assign popcount34_28tv_out[4] = popcount34_28tv_core_242;
  assign popcount34_28tv_out[5] = 1'b0;
endmodule