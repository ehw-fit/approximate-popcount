// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=0.637355
// WCE=15.0
// EP=0.396253%
// Printed PDK parameters:
//  Area=98520798.0
//  Delay=70690992.0
//  Power=5265700.0

module popcount32_9jxh(input [31:0] input_a, output [5:0] popcount32_9jxh_out);
  wire popcount32_9jxh_core_034;
  wire popcount32_9jxh_core_035;
  wire popcount32_9jxh_core_036;
  wire popcount32_9jxh_core_037;
  wire popcount32_9jxh_core_038;
  wire popcount32_9jxh_core_039;
  wire popcount32_9jxh_core_040;
  wire popcount32_9jxh_core_042;
  wire popcount32_9jxh_core_043;
  wire popcount32_9jxh_core_044;
  wire popcount32_9jxh_core_045;
  wire popcount32_9jxh_core_046;
  wire popcount32_9jxh_core_047;
  wire popcount32_9jxh_core_048;
  wire popcount32_9jxh_core_049;
  wire popcount32_9jxh_core_050;
  wire popcount32_9jxh_core_051;
  wire popcount32_9jxh_core_052;
  wire popcount32_9jxh_core_053;
  wire popcount32_9jxh_core_054;
  wire popcount32_9jxh_core_055;
  wire popcount32_9jxh_core_056;
  wire popcount32_9jxh_core_057;
  wire popcount32_9jxh_core_058;
  wire popcount32_9jxh_core_059;
  wire popcount32_9jxh_core_060;
  wire popcount32_9jxh_core_061;
  wire popcount32_9jxh_core_062;
  wire popcount32_9jxh_core_064;
  wire popcount32_9jxh_core_068;
  wire popcount32_9jxh_core_069;
  wire popcount32_9jxh_core_070;
  wire popcount32_9jxh_core_071;
  wire popcount32_9jxh_core_072;
  wire popcount32_9jxh_core_073;
  wire popcount32_9jxh_core_074;
  wire popcount32_9jxh_core_075;
  wire popcount32_9jxh_core_076;
  wire popcount32_9jxh_core_077;
  wire popcount32_9jxh_core_079;
  wire popcount32_9jxh_core_080;
  wire popcount32_9jxh_core_081;
  wire popcount32_9jxh_core_082;
  wire popcount32_9jxh_core_083;
  wire popcount32_9jxh_core_084;
  wire popcount32_9jxh_core_085;
  wire popcount32_9jxh_core_086;
  wire popcount32_9jxh_core_087;
  wire popcount32_9jxh_core_088;
  wire popcount32_9jxh_core_090;
  wire popcount32_9jxh_core_091;
  wire popcount32_9jxh_core_092;
  wire popcount32_9jxh_core_093;
  wire popcount32_9jxh_core_094;
  wire popcount32_9jxh_core_095;
  wire popcount32_9jxh_core_096;
  wire popcount32_9jxh_core_097;
  wire popcount32_9jxh_core_098;
  wire popcount32_9jxh_core_099;
  wire popcount32_9jxh_core_100;
  wire popcount32_9jxh_core_101;
  wire popcount32_9jxh_core_102;
  wire popcount32_9jxh_core_103;
  wire popcount32_9jxh_core_104;
  wire popcount32_9jxh_core_105;
  wire popcount32_9jxh_core_106;
  wire popcount32_9jxh_core_107;
  wire popcount32_9jxh_core_108;
  wire popcount32_9jxh_core_109;
  wire popcount32_9jxh_core_110;
  wire popcount32_9jxh_core_111;
  wire popcount32_9jxh_core_112;
  wire popcount32_9jxh_core_113;
  wire popcount32_9jxh_core_115;
  wire popcount32_9jxh_core_117;
  wire popcount32_9jxh_core_118;
  wire popcount32_9jxh_core_119;
  wire popcount32_9jxh_core_120;
  wire popcount32_9jxh_core_121;
  wire popcount32_9jxh_core_122;
  wire popcount32_9jxh_core_123;
  wire popcount32_9jxh_core_124;
  wire popcount32_9jxh_core_125;
  wire popcount32_9jxh_core_126_not;
  wire popcount32_9jxh_core_127;
  wire popcount32_9jxh_core_128;
  wire popcount32_9jxh_core_129;
  wire popcount32_9jxh_core_130;
  wire popcount32_9jxh_core_131;
  wire popcount32_9jxh_core_132;
  wire popcount32_9jxh_core_133;
  wire popcount32_9jxh_core_134;
  wire popcount32_9jxh_core_135;
  wire popcount32_9jxh_core_136;
  wire popcount32_9jxh_core_138;
  wire popcount32_9jxh_core_139_not;
  wire popcount32_9jxh_core_140;
  wire popcount32_9jxh_core_141;
  wire popcount32_9jxh_core_142;
  wire popcount32_9jxh_core_143;
  wire popcount32_9jxh_core_144;
  wire popcount32_9jxh_core_145;
  wire popcount32_9jxh_core_146;
  wire popcount32_9jxh_core_147;
  wire popcount32_9jxh_core_151;
  wire popcount32_9jxh_core_152;
  wire popcount32_9jxh_core_153;
  wire popcount32_9jxh_core_154;
  wire popcount32_9jxh_core_155;
  wire popcount32_9jxh_core_156;
  wire popcount32_9jxh_core_157;
  wire popcount32_9jxh_core_158;
  wire popcount32_9jxh_core_159;
  wire popcount32_9jxh_core_160;
  wire popcount32_9jxh_core_161;
  wire popcount32_9jxh_core_164;
  wire popcount32_9jxh_core_165;
  wire popcount32_9jxh_core_166;
  wire popcount32_9jxh_core_167;
  wire popcount32_9jxh_core_168;
  wire popcount32_9jxh_core_169;
  wire popcount32_9jxh_core_170;
  wire popcount32_9jxh_core_171;
  wire popcount32_9jxh_core_172;
  wire popcount32_9jxh_core_173;
  wire popcount32_9jxh_core_175;
  wire popcount32_9jxh_core_176;
  wire popcount32_9jxh_core_177;
  wire popcount32_9jxh_core_178;
  wire popcount32_9jxh_core_179;
  wire popcount32_9jxh_core_180;
  wire popcount32_9jxh_core_181;
  wire popcount32_9jxh_core_182;
  wire popcount32_9jxh_core_183;
  wire popcount32_9jxh_core_184;
  wire popcount32_9jxh_core_185;
  wire popcount32_9jxh_core_186;
  wire popcount32_9jxh_core_187;
  wire popcount32_9jxh_core_188;
  wire popcount32_9jxh_core_189;
  wire popcount32_9jxh_core_190;
  wire popcount32_9jxh_core_191;
  wire popcount32_9jxh_core_192;
  wire popcount32_9jxh_core_193;
  wire popcount32_9jxh_core_194;
  wire popcount32_9jxh_core_195;
  wire popcount32_9jxh_core_196;
  wire popcount32_9jxh_core_197;
  wire popcount32_9jxh_core_198;
  wire popcount32_9jxh_core_200;
  wire popcount32_9jxh_core_204;
  wire popcount32_9jxh_core_205;
  wire popcount32_9jxh_core_206;
  wire popcount32_9jxh_core_207;
  wire popcount32_9jxh_core_208;
  wire popcount32_9jxh_core_209;
  wire popcount32_9jxh_core_210;
  wire popcount32_9jxh_core_211;
  wire popcount32_9jxh_core_212;
  wire popcount32_9jxh_core_213;
  wire popcount32_9jxh_core_214;
  wire popcount32_9jxh_core_215;
  wire popcount32_9jxh_core_216;
  wire popcount32_9jxh_core_217;
  wire popcount32_9jxh_core_218;
  wire popcount32_9jxh_core_219;
  wire popcount32_9jxh_core_220;
  wire popcount32_9jxh_core_221;
  wire popcount32_9jxh_core_222;
  wire popcount32_9jxh_core_223;
  wire popcount32_9jxh_core_225;

  assign popcount32_9jxh_core_034 = input_a[0] ^ input_a[1];
  assign popcount32_9jxh_core_035 = input_a[0] & input_a[1];
  assign popcount32_9jxh_core_036 = input_a[2] ^ input_a[3];
  assign popcount32_9jxh_core_037 = input_a[2] & input_a[3];
  assign popcount32_9jxh_core_038 = popcount32_9jxh_core_034 ^ popcount32_9jxh_core_036;
  assign popcount32_9jxh_core_039 = popcount32_9jxh_core_034 & popcount32_9jxh_core_036;
  assign popcount32_9jxh_core_040 = popcount32_9jxh_core_035 | popcount32_9jxh_core_037;
  assign popcount32_9jxh_core_042 = popcount32_9jxh_core_040 | popcount32_9jxh_core_039;
  assign popcount32_9jxh_core_043 = ~input_a[15];
  assign popcount32_9jxh_core_044 = input_a[21] ^ input_a[2];
  assign popcount32_9jxh_core_045 = input_a[4] ^ input_a[5];
  assign popcount32_9jxh_core_046 = input_a[4] & input_a[5];
  assign popcount32_9jxh_core_047 = input_a[6] ^ input_a[7];
  assign popcount32_9jxh_core_048 = input_a[6] & input_a[7];
  assign popcount32_9jxh_core_049 = popcount32_9jxh_core_045 ^ popcount32_9jxh_core_047;
  assign popcount32_9jxh_core_050 = popcount32_9jxh_core_045 & popcount32_9jxh_core_047;
  assign popcount32_9jxh_core_051 = popcount32_9jxh_core_046 | popcount32_9jxh_core_048;
  assign popcount32_9jxh_core_052 = ~input_a[18];
  assign popcount32_9jxh_core_053 = popcount32_9jxh_core_051 | popcount32_9jxh_core_050;
  assign popcount32_9jxh_core_054 = ~input_a[9];
  assign popcount32_9jxh_core_055 = input_a[3] & input_a[8];
  assign popcount32_9jxh_core_056 = popcount32_9jxh_core_038 ^ popcount32_9jxh_core_049;
  assign popcount32_9jxh_core_057 = popcount32_9jxh_core_038 & popcount32_9jxh_core_049;
  assign popcount32_9jxh_core_058 = popcount32_9jxh_core_042 ^ popcount32_9jxh_core_053;
  assign popcount32_9jxh_core_059 = popcount32_9jxh_core_042 & popcount32_9jxh_core_053;
  assign popcount32_9jxh_core_060 = popcount32_9jxh_core_058 ^ popcount32_9jxh_core_057;
  assign popcount32_9jxh_core_061 = popcount32_9jxh_core_058 & popcount32_9jxh_core_057;
  assign popcount32_9jxh_core_062 = popcount32_9jxh_core_059 | popcount32_9jxh_core_061;
  assign popcount32_9jxh_core_064 = ~(input_a[20] & input_a[15]);
  assign popcount32_9jxh_core_068 = input_a[8] ^ input_a[9];
  assign popcount32_9jxh_core_069 = input_a[8] & input_a[9];
  assign popcount32_9jxh_core_070 = input_a[10] ^ input_a[11];
  assign popcount32_9jxh_core_071 = input_a[10] & input_a[11];
  assign popcount32_9jxh_core_072 = popcount32_9jxh_core_068 ^ popcount32_9jxh_core_070;
  assign popcount32_9jxh_core_073 = popcount32_9jxh_core_068 & popcount32_9jxh_core_070;
  assign popcount32_9jxh_core_074 = popcount32_9jxh_core_069 ^ popcount32_9jxh_core_071;
  assign popcount32_9jxh_core_075 = popcount32_9jxh_core_069 & input_a[11];
  assign popcount32_9jxh_core_076 = popcount32_9jxh_core_074 | popcount32_9jxh_core_073;
  assign popcount32_9jxh_core_077 = ~input_a[21];
  assign popcount32_9jxh_core_079 = input_a[12] ^ input_a[13];
  assign popcount32_9jxh_core_080 = input_a[12] & input_a[13];
  assign popcount32_9jxh_core_081 = input_a[14] ^ input_a[15];
  assign popcount32_9jxh_core_082 = input_a[14] & input_a[15];
  assign popcount32_9jxh_core_083 = popcount32_9jxh_core_079 ^ popcount32_9jxh_core_081;
  assign popcount32_9jxh_core_084 = popcount32_9jxh_core_079 & popcount32_9jxh_core_081;
  assign popcount32_9jxh_core_085 = popcount32_9jxh_core_080 ^ popcount32_9jxh_core_082;
  assign popcount32_9jxh_core_086 = popcount32_9jxh_core_080 & input_a[15];
  assign popcount32_9jxh_core_087 = popcount32_9jxh_core_085 | popcount32_9jxh_core_084;
  assign popcount32_9jxh_core_088 = ~input_a[6];
  assign popcount32_9jxh_core_090 = popcount32_9jxh_core_072 ^ popcount32_9jxh_core_083;
  assign popcount32_9jxh_core_091 = popcount32_9jxh_core_072 & popcount32_9jxh_core_083;
  assign popcount32_9jxh_core_092 = popcount32_9jxh_core_076 ^ popcount32_9jxh_core_087;
  assign popcount32_9jxh_core_093 = popcount32_9jxh_core_076 & popcount32_9jxh_core_087;
  assign popcount32_9jxh_core_094 = popcount32_9jxh_core_092 ^ popcount32_9jxh_core_091;
  assign popcount32_9jxh_core_095 = popcount32_9jxh_core_092 & popcount32_9jxh_core_091;
  assign popcount32_9jxh_core_096 = popcount32_9jxh_core_093 | popcount32_9jxh_core_095;
  assign popcount32_9jxh_core_097 = popcount32_9jxh_core_075 | popcount32_9jxh_core_086;
  assign popcount32_9jxh_core_098 = ~(input_a[9] | input_a[26]);
  assign popcount32_9jxh_core_099 = popcount32_9jxh_core_097 | popcount32_9jxh_core_096;
  assign popcount32_9jxh_core_100 = ~input_a[10];
  assign popcount32_9jxh_core_101 = ~(input_a[7] | input_a[1]);
  assign popcount32_9jxh_core_102 = popcount32_9jxh_core_056 ^ popcount32_9jxh_core_090;
  assign popcount32_9jxh_core_103 = popcount32_9jxh_core_056 & popcount32_9jxh_core_090;
  assign popcount32_9jxh_core_104 = popcount32_9jxh_core_060 ^ popcount32_9jxh_core_094;
  assign popcount32_9jxh_core_105 = popcount32_9jxh_core_060 & popcount32_9jxh_core_094;
  assign popcount32_9jxh_core_106 = popcount32_9jxh_core_104 ^ popcount32_9jxh_core_103;
  assign popcount32_9jxh_core_107 = popcount32_9jxh_core_104 & popcount32_9jxh_core_103;
  assign popcount32_9jxh_core_108 = popcount32_9jxh_core_105 | popcount32_9jxh_core_107;
  assign popcount32_9jxh_core_109 = popcount32_9jxh_core_062 ^ popcount32_9jxh_core_099;
  assign popcount32_9jxh_core_110 = popcount32_9jxh_core_062 & popcount32_9jxh_core_099;
  assign popcount32_9jxh_core_111 = popcount32_9jxh_core_109 ^ popcount32_9jxh_core_108;
  assign popcount32_9jxh_core_112 = popcount32_9jxh_core_109 & popcount32_9jxh_core_108;
  assign popcount32_9jxh_core_113 = popcount32_9jxh_core_110 | popcount32_9jxh_core_112;
  assign popcount32_9jxh_core_115 = ~(input_a[26] ^ input_a[13]);
  assign popcount32_9jxh_core_117 = ~input_a[6];
  assign popcount32_9jxh_core_118 = ~input_a[7];
  assign popcount32_9jxh_core_119 = input_a[16] ^ input_a[17];
  assign popcount32_9jxh_core_120 = input_a[16] & input_a[17];
  assign popcount32_9jxh_core_121 = input_a[18] ^ input_a[19];
  assign popcount32_9jxh_core_122 = input_a[18] & input_a[19];
  assign popcount32_9jxh_core_123 = popcount32_9jxh_core_119 ^ popcount32_9jxh_core_121;
  assign popcount32_9jxh_core_124 = popcount32_9jxh_core_119 & popcount32_9jxh_core_121;
  assign popcount32_9jxh_core_125 = popcount32_9jxh_core_120 | popcount32_9jxh_core_122;
  assign popcount32_9jxh_core_126_not = ~input_a[6];
  assign popcount32_9jxh_core_127 = popcount32_9jxh_core_125 | popcount32_9jxh_core_124;
  assign popcount32_9jxh_core_128 = ~(input_a[12] ^ input_a[0]);
  assign popcount32_9jxh_core_129 = ~(input_a[17] ^ input_a[31]);
  assign popcount32_9jxh_core_130 = input_a[20] ^ input_a[21];
  assign popcount32_9jxh_core_131 = input_a[20] & input_a[21];
  assign popcount32_9jxh_core_132 = input_a[22] ^ input_a[23];
  assign popcount32_9jxh_core_133 = input_a[22] & input_a[23];
  assign popcount32_9jxh_core_134 = ~(popcount32_9jxh_core_130 & popcount32_9jxh_core_132);
  assign popcount32_9jxh_core_135 = popcount32_9jxh_core_130 & popcount32_9jxh_core_132;
  assign popcount32_9jxh_core_136 = popcount32_9jxh_core_131 | popcount32_9jxh_core_133;
  assign popcount32_9jxh_core_138 = popcount32_9jxh_core_136 | popcount32_9jxh_core_135;
  assign popcount32_9jxh_core_139_not = ~input_a[30];
  assign popcount32_9jxh_core_140 = input_a[30] & input_a[28];
  assign popcount32_9jxh_core_141 = popcount32_9jxh_core_123 ^ popcount32_9jxh_core_134;
  assign popcount32_9jxh_core_142 = popcount32_9jxh_core_123 & popcount32_9jxh_core_134;
  assign popcount32_9jxh_core_143 = popcount32_9jxh_core_127 ^ popcount32_9jxh_core_138;
  assign popcount32_9jxh_core_144 = popcount32_9jxh_core_127 & popcount32_9jxh_core_138;
  assign popcount32_9jxh_core_145 = popcount32_9jxh_core_143 ^ popcount32_9jxh_core_142;
  assign popcount32_9jxh_core_146 = popcount32_9jxh_core_143 & popcount32_9jxh_core_142;
  assign popcount32_9jxh_core_147 = popcount32_9jxh_core_144 | popcount32_9jxh_core_146;
  assign popcount32_9jxh_core_151 = input_a[6] | input_a[7];
  assign popcount32_9jxh_core_152 = input_a[2] ^ input_a[15];
  assign popcount32_9jxh_core_153 = input_a[24] ^ input_a[25];
  assign popcount32_9jxh_core_154 = input_a[24] & input_a[25];
  assign popcount32_9jxh_core_155 = input_a[26] ^ input_a[27];
  assign popcount32_9jxh_core_156 = input_a[26] & input_a[27];
  assign popcount32_9jxh_core_157 = popcount32_9jxh_core_153 ^ popcount32_9jxh_core_155;
  assign popcount32_9jxh_core_158 = popcount32_9jxh_core_153 & popcount32_9jxh_core_155;
  assign popcount32_9jxh_core_159 = popcount32_9jxh_core_154 ^ popcount32_9jxh_core_156;
  assign popcount32_9jxh_core_160 = input_a[24] & popcount32_9jxh_core_156;
  assign popcount32_9jxh_core_161 = popcount32_9jxh_core_159 | popcount32_9jxh_core_158;
  assign popcount32_9jxh_core_164 = input_a[28] ^ input_a[29];
  assign popcount32_9jxh_core_165 = input_a[28] & input_a[29];
  assign popcount32_9jxh_core_166 = input_a[30] ^ input_a[31];
  assign popcount32_9jxh_core_167 = input_a[30] & input_a[31];
  assign popcount32_9jxh_core_168 = popcount32_9jxh_core_164 ^ popcount32_9jxh_core_166;
  assign popcount32_9jxh_core_169 = popcount32_9jxh_core_164 & popcount32_9jxh_core_166;
  assign popcount32_9jxh_core_170 = popcount32_9jxh_core_165 ^ popcount32_9jxh_core_167;
  assign popcount32_9jxh_core_171 = popcount32_9jxh_core_165 & input_a[30];
  assign popcount32_9jxh_core_172 = popcount32_9jxh_core_170 | popcount32_9jxh_core_169;
  assign popcount32_9jxh_core_173 = ~input_a[20];
  assign popcount32_9jxh_core_175 = popcount32_9jxh_core_157 ^ popcount32_9jxh_core_168;
  assign popcount32_9jxh_core_176 = popcount32_9jxh_core_157 & popcount32_9jxh_core_168;
  assign popcount32_9jxh_core_177 = popcount32_9jxh_core_161 ^ popcount32_9jxh_core_172;
  assign popcount32_9jxh_core_178 = popcount32_9jxh_core_161 & popcount32_9jxh_core_172;
  assign popcount32_9jxh_core_179 = popcount32_9jxh_core_177 ^ popcount32_9jxh_core_176;
  assign popcount32_9jxh_core_180 = popcount32_9jxh_core_177 & popcount32_9jxh_core_176;
  assign popcount32_9jxh_core_181 = popcount32_9jxh_core_178 | popcount32_9jxh_core_180;
  assign popcount32_9jxh_core_182 = popcount32_9jxh_core_160 | popcount32_9jxh_core_171;
  assign popcount32_9jxh_core_183 = input_a[9] & input_a[3];
  assign popcount32_9jxh_core_184 = popcount32_9jxh_core_182 | popcount32_9jxh_core_181;
  assign popcount32_9jxh_core_185 = ~input_a[22];
  assign popcount32_9jxh_core_186 = input_a[3] ^ input_a[24];
  assign popcount32_9jxh_core_187 = popcount32_9jxh_core_141 ^ popcount32_9jxh_core_175;
  assign popcount32_9jxh_core_188 = popcount32_9jxh_core_141 & popcount32_9jxh_core_175;
  assign popcount32_9jxh_core_189 = popcount32_9jxh_core_145 ^ popcount32_9jxh_core_179;
  assign popcount32_9jxh_core_190 = popcount32_9jxh_core_145 & popcount32_9jxh_core_179;
  assign popcount32_9jxh_core_191 = popcount32_9jxh_core_189 ^ popcount32_9jxh_core_188;
  assign popcount32_9jxh_core_192 = popcount32_9jxh_core_189 & popcount32_9jxh_core_188;
  assign popcount32_9jxh_core_193 = popcount32_9jxh_core_190 | popcount32_9jxh_core_192;
  assign popcount32_9jxh_core_194 = popcount32_9jxh_core_147 ^ popcount32_9jxh_core_184;
  assign popcount32_9jxh_core_195 = popcount32_9jxh_core_147 & popcount32_9jxh_core_184;
  assign popcount32_9jxh_core_196 = popcount32_9jxh_core_194 ^ popcount32_9jxh_core_193;
  assign popcount32_9jxh_core_197 = popcount32_9jxh_core_194 & popcount32_9jxh_core_193;
  assign popcount32_9jxh_core_198 = popcount32_9jxh_core_195 | popcount32_9jxh_core_197;
  assign popcount32_9jxh_core_200 = ~(input_a[3] ^ input_a[29]);
  assign popcount32_9jxh_core_204 = popcount32_9jxh_core_102 ^ popcount32_9jxh_core_187;
  assign popcount32_9jxh_core_205 = popcount32_9jxh_core_102 & popcount32_9jxh_core_187;
  assign popcount32_9jxh_core_206 = popcount32_9jxh_core_106 ^ popcount32_9jxh_core_191;
  assign popcount32_9jxh_core_207 = popcount32_9jxh_core_106 & popcount32_9jxh_core_191;
  assign popcount32_9jxh_core_208 = popcount32_9jxh_core_206 ^ popcount32_9jxh_core_205;
  assign popcount32_9jxh_core_209 = popcount32_9jxh_core_206 & popcount32_9jxh_core_205;
  assign popcount32_9jxh_core_210 = popcount32_9jxh_core_207 | popcount32_9jxh_core_209;
  assign popcount32_9jxh_core_211 = popcount32_9jxh_core_111 ^ popcount32_9jxh_core_196;
  assign popcount32_9jxh_core_212 = popcount32_9jxh_core_111 & popcount32_9jxh_core_196;
  assign popcount32_9jxh_core_213 = popcount32_9jxh_core_211 ^ popcount32_9jxh_core_210;
  assign popcount32_9jxh_core_214 = popcount32_9jxh_core_211 & popcount32_9jxh_core_210;
  assign popcount32_9jxh_core_215 = popcount32_9jxh_core_212 | popcount32_9jxh_core_214;
  assign popcount32_9jxh_core_216 = popcount32_9jxh_core_113 ^ popcount32_9jxh_core_198;
  assign popcount32_9jxh_core_217 = popcount32_9jxh_core_113 & popcount32_9jxh_core_198;
  assign popcount32_9jxh_core_218 = popcount32_9jxh_core_216 ^ popcount32_9jxh_core_215;
  assign popcount32_9jxh_core_219 = popcount32_9jxh_core_216 & popcount32_9jxh_core_215;
  assign popcount32_9jxh_core_220 = popcount32_9jxh_core_217 | popcount32_9jxh_core_219;
  assign popcount32_9jxh_core_221 = ~(input_a[6] | input_a[24]);
  assign popcount32_9jxh_core_222 = input_a[5] | input_a[31];
  assign popcount32_9jxh_core_223 = ~(input_a[0] ^ input_a[21]);
  assign popcount32_9jxh_core_225 = input_a[19] & input_a[7];

  assign popcount32_9jxh_out[0] = popcount32_9jxh_core_204;
  assign popcount32_9jxh_out[1] = popcount32_9jxh_core_208;
  assign popcount32_9jxh_out[2] = popcount32_9jxh_core_213;
  assign popcount32_9jxh_out[3] = popcount32_9jxh_core_218;
  assign popcount32_9jxh_out[4] = popcount32_9jxh_core_220;
  assign popcount32_9jxh_out[5] = 1'b0;
endmodule