// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.99916
// WCE=18.0
// EP=0.899124%
// Printed PDK parameters:
//  Area=4962060.0
//  Delay=10105700.0
//  Power=190790.0

module popcount36_0bei(input [35:0] input_a, output [5:0] popcount36_0bei_out);
  wire popcount36_0bei_core_038;
  wire popcount36_0bei_core_039;
  wire popcount36_0bei_core_040;
  wire popcount36_0bei_core_041;
  wire popcount36_0bei_core_042;
  wire popcount36_0bei_core_043_not;
  wire popcount36_0bei_core_044;
  wire popcount36_0bei_core_045;
  wire popcount36_0bei_core_047;
  wire popcount36_0bei_core_049;
  wire popcount36_0bei_core_050;
  wire popcount36_0bei_core_051;
  wire popcount36_0bei_core_052;
  wire popcount36_0bei_core_053;
  wire popcount36_0bei_core_055;
  wire popcount36_0bei_core_056;
  wire popcount36_0bei_core_057;
  wire popcount36_0bei_core_059;
  wire popcount36_0bei_core_062;
  wire popcount36_0bei_core_064;
  wire popcount36_0bei_core_065_not;
  wire popcount36_0bei_core_066;
  wire popcount36_0bei_core_070;
  wire popcount36_0bei_core_071;
  wire popcount36_0bei_core_072;
  wire popcount36_0bei_core_074;
  wire popcount36_0bei_core_077;
  wire popcount36_0bei_core_080;
  wire popcount36_0bei_core_081;
  wire popcount36_0bei_core_082;
  wire popcount36_0bei_core_086;
  wire popcount36_0bei_core_088;
  wire popcount36_0bei_core_090;
  wire popcount36_0bei_core_091_not;
  wire popcount36_0bei_core_092;
  wire popcount36_0bei_core_093;
  wire popcount36_0bei_core_095;
  wire popcount36_0bei_core_096;
  wire popcount36_0bei_core_097_not;
  wire popcount36_0bei_core_098;
  wire popcount36_0bei_core_099;
  wire popcount36_0bei_core_101;
  wire popcount36_0bei_core_103;
  wire popcount36_0bei_core_104;
  wire popcount36_0bei_core_105;
  wire popcount36_0bei_core_106;
  wire popcount36_0bei_core_107;
  wire popcount36_0bei_core_109;
  wire popcount36_0bei_core_110;
  wire popcount36_0bei_core_111;
  wire popcount36_0bei_core_112;
  wire popcount36_0bei_core_114;
  wire popcount36_0bei_core_115;
  wire popcount36_0bei_core_117;
  wire popcount36_0bei_core_118;
  wire popcount36_0bei_core_119;
  wire popcount36_0bei_core_120;
  wire popcount36_0bei_core_121;
  wire popcount36_0bei_core_122;
  wire popcount36_0bei_core_124;
  wire popcount36_0bei_core_126;
  wire popcount36_0bei_core_127;
  wire popcount36_0bei_core_131;
  wire popcount36_0bei_core_132;
  wire popcount36_0bei_core_135;
  wire popcount36_0bei_core_137;
  wire popcount36_0bei_core_138;
  wire popcount36_0bei_core_139;
  wire popcount36_0bei_core_140;
  wire popcount36_0bei_core_146;
  wire popcount36_0bei_core_150;
  wire popcount36_0bei_core_151;
  wire popcount36_0bei_core_153;
  wire popcount36_0bei_core_154;
  wire popcount36_0bei_core_158;
  wire popcount36_0bei_core_160;
  wire popcount36_0bei_core_162;
  wire popcount36_0bei_core_163;
  wire popcount36_0bei_core_164;
  wire popcount36_0bei_core_165;
  wire popcount36_0bei_core_166;
  wire popcount36_0bei_core_167;
  wire popcount36_0bei_core_168;
  wire popcount36_0bei_core_169;
  wire popcount36_0bei_core_171;
  wire popcount36_0bei_core_172;
  wire popcount36_0bei_core_173;
  wire popcount36_0bei_core_174;
  wire popcount36_0bei_core_177;
  wire popcount36_0bei_core_179;
  wire popcount36_0bei_core_180;
  wire popcount36_0bei_core_181;
  wire popcount36_0bei_core_183;
  wire popcount36_0bei_core_186;
  wire popcount36_0bei_core_188;
  wire popcount36_0bei_core_190;
  wire popcount36_0bei_core_192;
  wire popcount36_0bei_core_194;
  wire popcount36_0bei_core_196;
  wire popcount36_0bei_core_197;
  wire popcount36_0bei_core_199;
  wire popcount36_0bei_core_200;
  wire popcount36_0bei_core_201;
  wire popcount36_0bei_core_202;
  wire popcount36_0bei_core_203;
  wire popcount36_0bei_core_206;
  wire popcount36_0bei_core_207;
  wire popcount36_0bei_core_208;
  wire popcount36_0bei_core_211;
  wire popcount36_0bei_core_212;
  wire popcount36_0bei_core_213;
  wire popcount36_0bei_core_214;
  wire popcount36_0bei_core_215;
  wire popcount36_0bei_core_216;
  wire popcount36_0bei_core_218;
  wire popcount36_0bei_core_219;
  wire popcount36_0bei_core_223;
  wire popcount36_0bei_core_224;
  wire popcount36_0bei_core_225;
  wire popcount36_0bei_core_226;
  wire popcount36_0bei_core_228;
  wire popcount36_0bei_core_229;
  wire popcount36_0bei_core_233;
  wire popcount36_0bei_core_234;
  wire popcount36_0bei_core_235;
  wire popcount36_0bei_core_236;
  wire popcount36_0bei_core_238;
  wire popcount36_0bei_core_242;
  wire popcount36_0bei_core_248;
  wire popcount36_0bei_core_249;
  wire popcount36_0bei_core_250;
  wire popcount36_0bei_core_252;
  wire popcount36_0bei_core_254;
  wire popcount36_0bei_core_255;
  wire popcount36_0bei_core_259;
  wire popcount36_0bei_core_262;
  wire popcount36_0bei_core_264;
  wire popcount36_0bei_core_265;
  wire popcount36_0bei_core_266;
  wire popcount36_0bei_core_268;
  wire popcount36_0bei_core_269;
  wire popcount36_0bei_core_270;
  wire popcount36_0bei_core_272;
  wire popcount36_0bei_core_274;
  wire popcount36_0bei_core_275;
  wire popcount36_0bei_core_276;

  assign popcount36_0bei_core_038 = input_a[15] & input_a[35];
  assign popcount36_0bei_core_039 = input_a[22] & input_a[26];
  assign popcount36_0bei_core_040 = ~input_a[10];
  assign popcount36_0bei_core_041 = input_a[8] & input_a[10];
  assign popcount36_0bei_core_042 = ~(input_a[24] ^ input_a[10]);
  assign popcount36_0bei_core_043_not = ~input_a[14];
  assign popcount36_0bei_core_044 = ~(input_a[10] ^ input_a[2]);
  assign popcount36_0bei_core_045 = popcount36_0bei_core_039 & popcount36_0bei_core_041;
  assign popcount36_0bei_core_047 = input_a[35] & input_a[31];
  assign popcount36_0bei_core_049 = ~input_a[33];
  assign popcount36_0bei_core_050 = ~(input_a[3] ^ input_a[16]);
  assign popcount36_0bei_core_051 = ~(input_a[28] | input_a[35]);
  assign popcount36_0bei_core_052 = ~(input_a[20] ^ input_a[26]);
  assign popcount36_0bei_core_053 = ~input_a[20];
  assign popcount36_0bei_core_055 = input_a[26] & input_a[10];
  assign popcount36_0bei_core_056 = ~(input_a[22] & input_a[9]);
  assign popcount36_0bei_core_057 = ~(input_a[20] | input_a[7]);
  assign popcount36_0bei_core_059 = input_a[24] ^ input_a[13];
  assign popcount36_0bei_core_062 = ~(input_a[32] & input_a[7]);
  assign popcount36_0bei_core_064 = ~input_a[11];
  assign popcount36_0bei_core_065_not = ~input_a[17];
  assign popcount36_0bei_core_066 = ~(input_a[35] ^ input_a[4]);
  assign popcount36_0bei_core_070 = input_a[24] ^ input_a[15];
  assign popcount36_0bei_core_071 = ~(input_a[0] & input_a[26]);
  assign popcount36_0bei_core_072 = ~(input_a[20] & input_a[28]);
  assign popcount36_0bei_core_074 = input_a[4] & input_a[10];
  assign popcount36_0bei_core_077 = input_a[14] | input_a[4];
  assign popcount36_0bei_core_080 = ~(input_a[31] ^ input_a[6]);
  assign popcount36_0bei_core_081 = ~input_a[3];
  assign popcount36_0bei_core_082 = input_a[16] & input_a[25];
  assign popcount36_0bei_core_086 = ~input_a[9];
  assign popcount36_0bei_core_088 = ~(input_a[19] | input_a[4]);
  assign popcount36_0bei_core_090 = ~(input_a[33] & input_a[11]);
  assign popcount36_0bei_core_091_not = ~input_a[32];
  assign popcount36_0bei_core_092 = ~(input_a[17] & input_a[21]);
  assign popcount36_0bei_core_093 = ~(input_a[24] | input_a[15]);
  assign popcount36_0bei_core_095 = input_a[20] ^ input_a[8];
  assign popcount36_0bei_core_096 = input_a[30] ^ input_a[11];
  assign popcount36_0bei_core_097_not = ~input_a[6];
  assign popcount36_0bei_core_098 = ~input_a[30];
  assign popcount36_0bei_core_099 = ~(input_a[20] ^ input_a[3]);
  assign popcount36_0bei_core_101 = ~(input_a[29] | input_a[28]);
  assign popcount36_0bei_core_103 = input_a[2] ^ input_a[10];
  assign popcount36_0bei_core_104 = input_a[22] & input_a[7];
  assign popcount36_0bei_core_105 = input_a[10] & input_a[31];
  assign popcount36_0bei_core_106 = input_a[17] & input_a[12];
  assign popcount36_0bei_core_107 = ~(input_a[7] | input_a[23]);
  assign popcount36_0bei_core_109 = ~(input_a[7] | input_a[32]);
  assign popcount36_0bei_core_110 = input_a[11] ^ input_a[9];
  assign popcount36_0bei_core_111 = input_a[29] ^ input_a[18];
  assign popcount36_0bei_core_112 = input_a[20] & input_a[6];
  assign popcount36_0bei_core_114 = ~(input_a[29] ^ input_a[14]);
  assign popcount36_0bei_core_115 = input_a[32] & input_a[27];
  assign popcount36_0bei_core_117 = input_a[7] & input_a[32];
  assign popcount36_0bei_core_118 = ~(input_a[3] | input_a[11]);
  assign popcount36_0bei_core_119 = ~input_a[20];
  assign popcount36_0bei_core_120 = input_a[30] ^ input_a[6];
  assign popcount36_0bei_core_121 = input_a[20] ^ input_a[35];
  assign popcount36_0bei_core_122 = input_a[18] ^ input_a[4];
  assign popcount36_0bei_core_124 = ~(input_a[15] & input_a[24]);
  assign popcount36_0bei_core_126 = ~(input_a[10] | input_a[2]);
  assign popcount36_0bei_core_127 = input_a[15] & input_a[25];
  assign popcount36_0bei_core_131 = popcount36_0bei_core_045 ^ popcount36_0bei_core_127;
  assign popcount36_0bei_core_132 = popcount36_0bei_core_045 & popcount36_0bei_core_127;
  assign popcount36_0bei_core_135 = input_a[26] ^ input_a[33];
  assign popcount36_0bei_core_137 = ~input_a[23];
  assign popcount36_0bei_core_138 = input_a[26] & input_a[20];
  assign popcount36_0bei_core_139 = ~(input_a[20] ^ input_a[6]);
  assign popcount36_0bei_core_140 = ~(input_a[19] | input_a[20]);
  assign popcount36_0bei_core_146 = ~(input_a[23] ^ input_a[4]);
  assign popcount36_0bei_core_150 = input_a[20] & input_a[21];
  assign popcount36_0bei_core_151 = ~(input_a[11] & input_a[5]);
  assign popcount36_0bei_core_153 = input_a[15] | input_a[2];
  assign popcount36_0bei_core_154 = ~(input_a[35] ^ input_a[12]);
  assign popcount36_0bei_core_158 = input_a[4] & input_a[0];
  assign popcount36_0bei_core_160 = input_a[17] | input_a[29];
  assign popcount36_0bei_core_162 = popcount36_0bei_core_158 & input_a[27];
  assign popcount36_0bei_core_163 = ~(input_a[11] & input_a[15]);
  assign popcount36_0bei_core_164 = input_a[33] & input_a[1];
  assign popcount36_0bei_core_165 = input_a[16] | input_a[13];
  assign popcount36_0bei_core_166 = input_a[8] ^ input_a[12];
  assign popcount36_0bei_core_167 = input_a[24] | input_a[29];
  assign popcount36_0bei_core_168 = input_a[17] | input_a[29];
  assign popcount36_0bei_core_169 = input_a[25] & input_a[6];
  assign popcount36_0bei_core_171 = popcount36_0bei_core_162 & input_a[11];
  assign popcount36_0bei_core_172 = ~input_a[15];
  assign popcount36_0bei_core_173 = ~(input_a[19] ^ input_a[3]);
  assign popcount36_0bei_core_174 = ~(input_a[35] & input_a[26]);
  assign popcount36_0bei_core_177 = ~input_a[14];
  assign popcount36_0bei_core_179 = ~(input_a[11] & input_a[1]);
  assign popcount36_0bei_core_180 = ~(input_a[9] & input_a[32]);
  assign popcount36_0bei_core_181 = ~(input_a[19] ^ input_a[17]);
  assign popcount36_0bei_core_183 = ~(input_a[33] | input_a[3]);
  assign popcount36_0bei_core_186 = input_a[29] | input_a[15];
  assign popcount36_0bei_core_188 = input_a[34] ^ input_a[3];
  assign popcount36_0bei_core_190 = input_a[29] ^ input_a[28];
  assign popcount36_0bei_core_192 = input_a[21] | input_a[19];
  assign popcount36_0bei_core_194 = input_a[5] & input_a[8];
  assign popcount36_0bei_core_196 = ~(input_a[12] ^ input_a[9]);
  assign popcount36_0bei_core_197 = input_a[12] | input_a[32];
  assign popcount36_0bei_core_199 = ~input_a[30];
  assign popcount36_0bei_core_200 = ~input_a[12];
  assign popcount36_0bei_core_201 = ~input_a[11];
  assign popcount36_0bei_core_202 = input_a[24] ^ input_a[13];
  assign popcount36_0bei_core_203 = ~input_a[30];
  assign popcount36_0bei_core_206 = ~input_a[26];
  assign popcount36_0bei_core_207 = input_a[15] | input_a[20];
  assign popcount36_0bei_core_208 = ~(input_a[22] | input_a[26]);
  assign popcount36_0bei_core_211 = input_a[32] ^ input_a[4];
  assign popcount36_0bei_core_212 = ~(input_a[27] & input_a[6]);
  assign popcount36_0bei_core_213 = ~(input_a[23] ^ input_a[23]);
  assign popcount36_0bei_core_214 = ~input_a[10];
  assign popcount36_0bei_core_215 = ~input_a[10];
  assign popcount36_0bei_core_216 = ~(input_a[9] ^ input_a[17]);
  assign popcount36_0bei_core_218 = input_a[19] | input_a[28];
  assign popcount36_0bei_core_219 = input_a[11] ^ input_a[2];
  assign popcount36_0bei_core_223 = ~(input_a[23] ^ input_a[33]);
  assign popcount36_0bei_core_224 = ~(input_a[31] & input_a[10]);
  assign popcount36_0bei_core_225 = ~(input_a[0] ^ input_a[11]);
  assign popcount36_0bei_core_226 = ~input_a[32];
  assign popcount36_0bei_core_228 = input_a[5] & input_a[8];
  assign popcount36_0bei_core_229 = input_a[35] ^ input_a[16];
  assign popcount36_0bei_core_233 = input_a[12] | input_a[35];
  assign popcount36_0bei_core_234 = input_a[21] | input_a[27];
  assign popcount36_0bei_core_235 = input_a[33] | input_a[32];
  assign popcount36_0bei_core_236 = ~input_a[1];
  assign popcount36_0bei_core_238 = ~input_a[23];
  assign popcount36_0bei_core_242 = ~popcount36_0bei_core_171;
  assign popcount36_0bei_core_248 = input_a[5] & input_a[15];
  assign popcount36_0bei_core_249 = input_a[9] & input_a[9];
  assign popcount36_0bei_core_250 = input_a[7] | input_a[15];
  assign popcount36_0bei_core_252 = input_a[22] & input_a[30];
  assign popcount36_0bei_core_254 = ~(input_a[33] | input_a[22]);
  assign popcount36_0bei_core_255 = ~(input_a[5] | input_a[29]);
  assign popcount36_0bei_core_259 = ~popcount36_0bei_core_131;
  assign popcount36_0bei_core_262 = popcount36_0bei_core_132 ^ popcount36_0bei_core_242;
  assign popcount36_0bei_core_264 = popcount36_0bei_core_262 ^ popcount36_0bei_core_131;
  assign popcount36_0bei_core_265 = popcount36_0bei_core_262 & popcount36_0bei_core_131;
  assign popcount36_0bei_core_266 = popcount36_0bei_core_132 | popcount36_0bei_core_265;
  assign popcount36_0bei_core_268 = input_a[22] & input_a[24];
  assign popcount36_0bei_core_269 = popcount36_0bei_core_171 | popcount36_0bei_core_266;
  assign popcount36_0bei_core_270 = ~(input_a[18] | input_a[22]);
  assign popcount36_0bei_core_272 = ~(input_a[2] ^ input_a[1]);
  assign popcount36_0bei_core_274 = input_a[26] & input_a[15];
  assign popcount36_0bei_core_275 = ~(input_a[20] ^ input_a[5]);
  assign popcount36_0bei_core_276 = ~(input_a[28] & input_a[22]);

  assign popcount36_0bei_out[0] = input_a[12];
  assign popcount36_0bei_out[1] = popcount36_0bei_core_242;
  assign popcount36_0bei_out[2] = popcount36_0bei_core_259;
  assign popcount36_0bei_out[3] = popcount36_0bei_core_264;
  assign popcount36_0bei_out[4] = popcount36_0bei_core_269;
  assign popcount36_0bei_out[5] = 1'b0;
endmodule