// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.99764
// WCE=17.0
// EP=0.903336%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_q08w(input [29:0] input_a, output [4:0] popcount30_q08w_out);
  wire popcount30_q08w_core_033_not;
  wire popcount30_q08w_core_034;
  wire popcount30_q08w_core_036;
  wire popcount30_q08w_core_037;
  wire popcount30_q08w_core_039;
  wire popcount30_q08w_core_040;
  wire popcount30_q08w_core_041;
  wire popcount30_q08w_core_043;
  wire popcount30_q08w_core_044;
  wire popcount30_q08w_core_046;
  wire popcount30_q08w_core_049;
  wire popcount30_q08w_core_050;
  wire popcount30_q08w_core_051;
  wire popcount30_q08w_core_054;
  wire popcount30_q08w_core_057;
  wire popcount30_q08w_core_060;
  wire popcount30_q08w_core_062;
  wire popcount30_q08w_core_063;
  wire popcount30_q08w_core_066_not;
  wire popcount30_q08w_core_069_not;
  wire popcount30_q08w_core_070;
  wire popcount30_q08w_core_072;
  wire popcount30_q08w_core_073;
  wire popcount30_q08w_core_074;
  wire popcount30_q08w_core_076;
  wire popcount30_q08w_core_077;
  wire popcount30_q08w_core_078;
  wire popcount30_q08w_core_079;
  wire popcount30_q08w_core_080;
  wire popcount30_q08w_core_081_not;
  wire popcount30_q08w_core_082;
  wire popcount30_q08w_core_086;
  wire popcount30_q08w_core_087;
  wire popcount30_q08w_core_089;
  wire popcount30_q08w_core_090;
  wire popcount30_q08w_core_091;
  wire popcount30_q08w_core_092;
  wire popcount30_q08w_core_093;
  wire popcount30_q08w_core_094;
  wire popcount30_q08w_core_095;
  wire popcount30_q08w_core_096;
  wire popcount30_q08w_core_098;
  wire popcount30_q08w_core_099;
  wire popcount30_q08w_core_100;
  wire popcount30_q08w_core_101;
  wire popcount30_q08w_core_103;
  wire popcount30_q08w_core_106;
  wire popcount30_q08w_core_107;
  wire popcount30_q08w_core_110;
  wire popcount30_q08w_core_111;
  wire popcount30_q08w_core_112;
  wire popcount30_q08w_core_113;
  wire popcount30_q08w_core_114;
  wire popcount30_q08w_core_116;
  wire popcount30_q08w_core_119;
  wire popcount30_q08w_core_120;
  wire popcount30_q08w_core_121;
  wire popcount30_q08w_core_122;
  wire popcount30_q08w_core_123;
  wire popcount30_q08w_core_127_not;
  wire popcount30_q08w_core_128;
  wire popcount30_q08w_core_130;
  wire popcount30_q08w_core_133;
  wire popcount30_q08w_core_134;
  wire popcount30_q08w_core_136;
  wire popcount30_q08w_core_137;
  wire popcount30_q08w_core_139;
  wire popcount30_q08w_core_143;
  wire popcount30_q08w_core_145;
  wire popcount30_q08w_core_146;
  wire popcount30_q08w_core_148_not;
  wire popcount30_q08w_core_149;
  wire popcount30_q08w_core_150;
  wire popcount30_q08w_core_151;
  wire popcount30_q08w_core_152;
  wire popcount30_q08w_core_154;
  wire popcount30_q08w_core_156;
  wire popcount30_q08w_core_157;
  wire popcount30_q08w_core_158;
  wire popcount30_q08w_core_159;
  wire popcount30_q08w_core_164;
  wire popcount30_q08w_core_166;
  wire popcount30_q08w_core_167;
  wire popcount30_q08w_core_168;
  wire popcount30_q08w_core_169;
  wire popcount30_q08w_core_170;
  wire popcount30_q08w_core_171;
  wire popcount30_q08w_core_172;
  wire popcount30_q08w_core_174;
  wire popcount30_q08w_core_175;
  wire popcount30_q08w_core_176;
  wire popcount30_q08w_core_177_not;
  wire popcount30_q08w_core_178;
  wire popcount30_q08w_core_179;
  wire popcount30_q08w_core_180;
  wire popcount30_q08w_core_182;
  wire popcount30_q08w_core_183;
  wire popcount30_q08w_core_184;
  wire popcount30_q08w_core_185;
  wire popcount30_q08w_core_186;
  wire popcount30_q08w_core_189;
  wire popcount30_q08w_core_190;
  wire popcount30_q08w_core_193;
  wire popcount30_q08w_core_194;
  wire popcount30_q08w_core_195;
  wire popcount30_q08w_core_197;
  wire popcount30_q08w_core_199;
  wire popcount30_q08w_core_201;
  wire popcount30_q08w_core_202;
  wire popcount30_q08w_core_206;
  wire popcount30_q08w_core_207;
  wire popcount30_q08w_core_208;
  wire popcount30_q08w_core_209;
  wire popcount30_q08w_core_210;
  wire popcount30_q08w_core_211;
  wire popcount30_q08w_core_213;

  assign popcount30_q08w_core_033_not = ~input_a[7];
  assign popcount30_q08w_core_034 = ~input_a[14];
  assign popcount30_q08w_core_036 = ~(input_a[25] | input_a[5]);
  assign popcount30_q08w_core_037 = ~input_a[6];
  assign popcount30_q08w_core_039 = input_a[19] & input_a[26];
  assign popcount30_q08w_core_040 = ~(input_a[25] | input_a[5]);
  assign popcount30_q08w_core_041 = ~(input_a[29] | input_a[13]);
  assign popcount30_q08w_core_043 = ~input_a[5];
  assign popcount30_q08w_core_044 = input_a[23] & input_a[17];
  assign popcount30_q08w_core_046 = ~(input_a[17] ^ input_a[21]);
  assign popcount30_q08w_core_049 = input_a[17] & input_a[29];
  assign popcount30_q08w_core_050 = ~input_a[26];
  assign popcount30_q08w_core_051 = ~(input_a[11] & input_a[19]);
  assign popcount30_q08w_core_054 = input_a[5] & input_a[29];
  assign popcount30_q08w_core_057 = input_a[21] & input_a[12];
  assign popcount30_q08w_core_060 = input_a[10] & input_a[14];
  assign popcount30_q08w_core_062 = input_a[21] ^ input_a[13];
  assign popcount30_q08w_core_063 = input_a[19] | input_a[19];
  assign popcount30_q08w_core_066_not = ~input_a[12];
  assign popcount30_q08w_core_069_not = ~input_a[21];
  assign popcount30_q08w_core_070 = input_a[11] ^ input_a[3];
  assign popcount30_q08w_core_072 = ~(input_a[5] | input_a[23]);
  assign popcount30_q08w_core_073 = ~(input_a[14] | input_a[14]);
  assign popcount30_q08w_core_074 = ~input_a[18];
  assign popcount30_q08w_core_076 = ~(input_a[27] & input_a[21]);
  assign popcount30_q08w_core_077 = input_a[25] ^ input_a[11];
  assign popcount30_q08w_core_078 = ~(input_a[23] ^ input_a[4]);
  assign popcount30_q08w_core_079 = input_a[14] ^ input_a[3];
  assign popcount30_q08w_core_080 = ~(input_a[0] & input_a[2]);
  assign popcount30_q08w_core_081_not = ~input_a[15];
  assign popcount30_q08w_core_082 = ~input_a[19];
  assign popcount30_q08w_core_086 = ~(input_a[0] & input_a[17]);
  assign popcount30_q08w_core_087 = input_a[5] ^ input_a[22];
  assign popcount30_q08w_core_089 = input_a[22] ^ input_a[14];
  assign popcount30_q08w_core_090 = ~input_a[29];
  assign popcount30_q08w_core_091 = ~(input_a[7] ^ input_a[29]);
  assign popcount30_q08w_core_092 = ~(input_a[8] & input_a[13]);
  assign popcount30_q08w_core_093 = ~(input_a[6] | input_a[2]);
  assign popcount30_q08w_core_094 = ~(input_a[20] | input_a[15]);
  assign popcount30_q08w_core_095 = input_a[10] & input_a[29];
  assign popcount30_q08w_core_096 = ~(input_a[3] ^ input_a[20]);
  assign popcount30_q08w_core_098 = input_a[26] | input_a[7];
  assign popcount30_q08w_core_099 = ~(input_a[27] & input_a[26]);
  assign popcount30_q08w_core_100 = input_a[23] | input_a[3];
  assign popcount30_q08w_core_101 = input_a[3] | input_a[29];
  assign popcount30_q08w_core_103 = ~(input_a[8] & input_a[4]);
  assign popcount30_q08w_core_106 = input_a[1] & input_a[21];
  assign popcount30_q08w_core_107 = ~input_a[1];
  assign popcount30_q08w_core_110 = input_a[28] | input_a[15];
  assign popcount30_q08w_core_111 = input_a[24] ^ input_a[2];
  assign popcount30_q08w_core_112 = ~input_a[8];
  assign popcount30_q08w_core_113 = ~(input_a[7] & input_a[16]);
  assign popcount30_q08w_core_114 = ~(input_a[14] ^ input_a[22]);
  assign popcount30_q08w_core_116 = ~(input_a[11] ^ input_a[26]);
  assign popcount30_q08w_core_119 = input_a[3] | input_a[6];
  assign popcount30_q08w_core_120 = input_a[26] | input_a[14];
  assign popcount30_q08w_core_121 = input_a[2] ^ input_a[11];
  assign popcount30_q08w_core_122 = ~input_a[21];
  assign popcount30_q08w_core_123 = ~(input_a[12] | input_a[12]);
  assign popcount30_q08w_core_127_not = ~input_a[22];
  assign popcount30_q08w_core_128 = ~input_a[17];
  assign popcount30_q08w_core_130 = ~(input_a[11] ^ input_a[8]);
  assign popcount30_q08w_core_133 = ~(input_a[22] & input_a[23]);
  assign popcount30_q08w_core_134 = ~(input_a[15] ^ input_a[19]);
  assign popcount30_q08w_core_136 = ~(input_a[24] & input_a[28]);
  assign popcount30_q08w_core_137 = input_a[9] & input_a[26];
  assign popcount30_q08w_core_139 = ~(input_a[0] | input_a[29]);
  assign popcount30_q08w_core_143 = ~(input_a[15] & input_a[2]);
  assign popcount30_q08w_core_145 = ~(input_a[1] | input_a[16]);
  assign popcount30_q08w_core_146 = ~(input_a[23] ^ input_a[23]);
  assign popcount30_q08w_core_148_not = ~input_a[15];
  assign popcount30_q08w_core_149 = ~input_a[4];
  assign popcount30_q08w_core_150 = input_a[8] & input_a[10];
  assign popcount30_q08w_core_151 = ~(input_a[0] ^ input_a[8]);
  assign popcount30_q08w_core_152 = input_a[15] & input_a[20];
  assign popcount30_q08w_core_154 = ~(input_a[29] | input_a[17]);
  assign popcount30_q08w_core_156 = ~(input_a[13] | input_a[5]);
  assign popcount30_q08w_core_157 = ~(input_a[17] ^ input_a[27]);
  assign popcount30_q08w_core_158 = ~(input_a[0] | input_a[23]);
  assign popcount30_q08w_core_159 = ~(input_a[18] ^ input_a[22]);
  assign popcount30_q08w_core_164 = ~(input_a[27] & input_a[4]);
  assign popcount30_q08w_core_166 = ~(input_a[18] | input_a[22]);
  assign popcount30_q08w_core_167 = input_a[5] ^ input_a[0];
  assign popcount30_q08w_core_168 = ~input_a[4];
  assign popcount30_q08w_core_169 = ~(input_a[8] | input_a[19]);
  assign popcount30_q08w_core_170 = ~(input_a[24] & input_a[29]);
  assign popcount30_q08w_core_171 = ~input_a[26];
  assign popcount30_q08w_core_172 = ~(input_a[7] ^ input_a[14]);
  assign popcount30_q08w_core_174 = ~(input_a[1] ^ input_a[0]);
  assign popcount30_q08w_core_175 = ~(input_a[10] | input_a[26]);
  assign popcount30_q08w_core_176 = ~(input_a[17] & input_a[11]);
  assign popcount30_q08w_core_177_not = ~input_a[24];
  assign popcount30_q08w_core_178 = ~(input_a[4] | input_a[11]);
  assign popcount30_q08w_core_179 = ~input_a[12];
  assign popcount30_q08w_core_180 = ~(input_a[6] & input_a[29]);
  assign popcount30_q08w_core_182 = input_a[28] ^ input_a[7];
  assign popcount30_q08w_core_183 = ~(input_a[16] & input_a[24]);
  assign popcount30_q08w_core_184 = ~(input_a[11] & input_a[17]);
  assign popcount30_q08w_core_185 = input_a[24] | input_a[6];
  assign popcount30_q08w_core_186 = ~(input_a[22] ^ input_a[2]);
  assign popcount30_q08w_core_189 = input_a[9] & input_a[13];
  assign popcount30_q08w_core_190 = input_a[3] | input_a[25];
  assign popcount30_q08w_core_193 = ~input_a[16];
  assign popcount30_q08w_core_194 = ~input_a[27];
  assign popcount30_q08w_core_195 = input_a[29] | input_a[0];
  assign popcount30_q08w_core_197 = ~(input_a[21] & input_a[21]);
  assign popcount30_q08w_core_199 = input_a[17] ^ input_a[11];
  assign popcount30_q08w_core_201 = ~(input_a[7] & input_a[1]);
  assign popcount30_q08w_core_202 = ~(input_a[13] | input_a[12]);
  assign popcount30_q08w_core_206 = ~input_a[28];
  assign popcount30_q08w_core_207 = ~input_a[2];
  assign popcount30_q08w_core_208 = ~(input_a[17] | input_a[6]);
  assign popcount30_q08w_core_209 = input_a[0] & input_a[23];
  assign popcount30_q08w_core_210 = input_a[23] ^ input_a[6];
  assign popcount30_q08w_core_211 = input_a[27] ^ input_a[15];
  assign popcount30_q08w_core_213 = input_a[23] | input_a[1];

  assign popcount30_q08w_out[0] = input_a[26];
  assign popcount30_q08w_out[1] = input_a[23];
  assign popcount30_q08w_out[2] = 1'b0;
  assign popcount30_q08w_out[3] = 1'b0;
  assign popcount30_q08w_out[4] = 1'b1;
endmodule