// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=9.04401
// WCE=27.0
// EP=0.974125%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_ltw2(input [20:0] input_a, output [4:0] popcount21_ltw2_out);
  wire popcount21_ltw2_core_023;
  wire popcount21_ltw2_core_024_not;
  wire popcount21_ltw2_core_025;
  wire popcount21_ltw2_core_026;
  wire popcount21_ltw2_core_027;
  wire popcount21_ltw2_core_028_not;
  wire popcount21_ltw2_core_029;
  wire popcount21_ltw2_core_030;
  wire popcount21_ltw2_core_031;
  wire popcount21_ltw2_core_032;
  wire popcount21_ltw2_core_034;
  wire popcount21_ltw2_core_035;
  wire popcount21_ltw2_core_036;
  wire popcount21_ltw2_core_037;
  wire popcount21_ltw2_core_039_not;
  wire popcount21_ltw2_core_040;
  wire popcount21_ltw2_core_042;
  wire popcount21_ltw2_core_044;
  wire popcount21_ltw2_core_046;
  wire popcount21_ltw2_core_048;
  wire popcount21_ltw2_core_049;
  wire popcount21_ltw2_core_051;
  wire popcount21_ltw2_core_055;
  wire popcount21_ltw2_core_061;
  wire popcount21_ltw2_core_063;
  wire popcount21_ltw2_core_064;
  wire popcount21_ltw2_core_065;
  wire popcount21_ltw2_core_066;
  wire popcount21_ltw2_core_067;
  wire popcount21_ltw2_core_068;
  wire popcount21_ltw2_core_069;
  wire popcount21_ltw2_core_070;
  wire popcount21_ltw2_core_076;
  wire popcount21_ltw2_core_082;
  wire popcount21_ltw2_core_084;
  wire popcount21_ltw2_core_085;
  wire popcount21_ltw2_core_086;
  wire popcount21_ltw2_core_087;
  wire popcount21_ltw2_core_088_not;
  wire popcount21_ltw2_core_090;
  wire popcount21_ltw2_core_092;
  wire popcount21_ltw2_core_094;
  wire popcount21_ltw2_core_096;
  wire popcount21_ltw2_core_099_not;
  wire popcount21_ltw2_core_101;
  wire popcount21_ltw2_core_103;
  wire popcount21_ltw2_core_104;
  wire popcount21_ltw2_core_105;
  wire popcount21_ltw2_core_107;
  wire popcount21_ltw2_core_108;
  wire popcount21_ltw2_core_110;
  wire popcount21_ltw2_core_111;
  wire popcount21_ltw2_core_112;
  wire popcount21_ltw2_core_113;
  wire popcount21_ltw2_core_116;
  wire popcount21_ltw2_core_117;
  wire popcount21_ltw2_core_118;
  wire popcount21_ltw2_core_122;
  wire popcount21_ltw2_core_123_not;
  wire popcount21_ltw2_core_125;
  wire popcount21_ltw2_core_126;
  wire popcount21_ltw2_core_128;
  wire popcount21_ltw2_core_129;
  wire popcount21_ltw2_core_130;
  wire popcount21_ltw2_core_133;
  wire popcount21_ltw2_core_134;
  wire popcount21_ltw2_core_135;
  wire popcount21_ltw2_core_137;
  wire popcount21_ltw2_core_139;
  wire popcount21_ltw2_core_140;
  wire popcount21_ltw2_core_141_not;
  wire popcount21_ltw2_core_144;
  wire popcount21_ltw2_core_145;
  wire popcount21_ltw2_core_149;

  assign popcount21_ltw2_core_023 = input_a[1] & input_a[9];
  assign popcount21_ltw2_core_024_not = ~input_a[14];
  assign popcount21_ltw2_core_025 = ~(input_a[5] & input_a[5]);
  assign popcount21_ltw2_core_026 = ~(input_a[15] & input_a[10]);
  assign popcount21_ltw2_core_027 = ~(input_a[10] | input_a[3]);
  assign popcount21_ltw2_core_028_not = ~input_a[8];
  assign popcount21_ltw2_core_029 = input_a[14] | input_a[13];
  assign popcount21_ltw2_core_030 = ~(input_a[19] | input_a[20]);
  assign popcount21_ltw2_core_031 = ~(input_a[20] ^ input_a[20]);
  assign popcount21_ltw2_core_032 = ~(input_a[6] ^ input_a[14]);
  assign popcount21_ltw2_core_034 = ~(input_a[13] ^ input_a[11]);
  assign popcount21_ltw2_core_035 = input_a[14] ^ input_a[3];
  assign popcount21_ltw2_core_036 = input_a[8] ^ input_a[2];
  assign popcount21_ltw2_core_037 = input_a[14] | input_a[4];
  assign popcount21_ltw2_core_039_not = ~input_a[3];
  assign popcount21_ltw2_core_040 = input_a[7] | input_a[20];
  assign popcount21_ltw2_core_042 = input_a[4] & input_a[16];
  assign popcount21_ltw2_core_044 = input_a[15] & input_a[5];
  assign popcount21_ltw2_core_046 = input_a[0] | input_a[1];
  assign popcount21_ltw2_core_048 = ~(input_a[14] ^ input_a[15]);
  assign popcount21_ltw2_core_049 = ~(input_a[19] ^ input_a[8]);
  assign popcount21_ltw2_core_051 = ~(input_a[2] ^ input_a[17]);
  assign popcount21_ltw2_core_055 = input_a[12] & input_a[3];
  assign popcount21_ltw2_core_061 = input_a[1] | input_a[0];
  assign popcount21_ltw2_core_063 = ~(input_a[19] & input_a[17]);
  assign popcount21_ltw2_core_064 = input_a[12] & input_a[7];
  assign popcount21_ltw2_core_065 = input_a[1] ^ input_a[6];
  assign popcount21_ltw2_core_066 = ~(input_a[7] ^ input_a[14]);
  assign popcount21_ltw2_core_067 = ~(input_a[3] ^ input_a[17]);
  assign popcount21_ltw2_core_068 = input_a[5] | input_a[17];
  assign popcount21_ltw2_core_069 = ~(input_a[11] ^ input_a[9]);
  assign popcount21_ltw2_core_070 = ~(input_a[12] ^ input_a[1]);
  assign popcount21_ltw2_core_076 = input_a[15] | input_a[4];
  assign popcount21_ltw2_core_082 = ~(input_a[18] & input_a[17]);
  assign popcount21_ltw2_core_084 = input_a[3] | input_a[18];
  assign popcount21_ltw2_core_085 = ~(input_a[1] & input_a[20]);
  assign popcount21_ltw2_core_086 = input_a[3] ^ input_a[19];
  assign popcount21_ltw2_core_087 = ~(input_a[6] ^ input_a[18]);
  assign popcount21_ltw2_core_088_not = ~input_a[8];
  assign popcount21_ltw2_core_090 = ~(input_a[4] | input_a[0]);
  assign popcount21_ltw2_core_092 = input_a[4] ^ input_a[12];
  assign popcount21_ltw2_core_094 = ~(input_a[1] | input_a[11]);
  assign popcount21_ltw2_core_096 = input_a[2] & input_a[8];
  assign popcount21_ltw2_core_099_not = ~input_a[8];
  assign popcount21_ltw2_core_101 = ~(input_a[4] & input_a[14]);
  assign popcount21_ltw2_core_103 = input_a[17] & input_a[10];
  assign popcount21_ltw2_core_104 = ~(input_a[12] ^ input_a[20]);
  assign popcount21_ltw2_core_105 = ~(input_a[14] | input_a[17]);
  assign popcount21_ltw2_core_107 = ~input_a[13];
  assign popcount21_ltw2_core_108 = ~(input_a[18] ^ input_a[14]);
  assign popcount21_ltw2_core_110 = ~(input_a[10] ^ input_a[16]);
  assign popcount21_ltw2_core_111 = input_a[6] & input_a[19];
  assign popcount21_ltw2_core_112 = ~input_a[9];
  assign popcount21_ltw2_core_113 = ~(input_a[9] & input_a[12]);
  assign popcount21_ltw2_core_116 = ~input_a[1];
  assign popcount21_ltw2_core_117 = ~(input_a[11] & input_a[16]);
  assign popcount21_ltw2_core_118 = input_a[18] | input_a[11];
  assign popcount21_ltw2_core_122 = input_a[18] | input_a[20];
  assign popcount21_ltw2_core_123_not = ~input_a[2];
  assign popcount21_ltw2_core_125 = ~(input_a[11] | input_a[13]);
  assign popcount21_ltw2_core_126 = ~input_a[16];
  assign popcount21_ltw2_core_128 = input_a[17] ^ input_a[15];
  assign popcount21_ltw2_core_129 = input_a[14] ^ input_a[0];
  assign popcount21_ltw2_core_130 = ~(input_a[11] | input_a[1]);
  assign popcount21_ltw2_core_133 = input_a[18] ^ input_a[19];
  assign popcount21_ltw2_core_134 = input_a[12] ^ input_a[12];
  assign popcount21_ltw2_core_135 = input_a[17] ^ input_a[18];
  assign popcount21_ltw2_core_137 = input_a[20] | input_a[6];
  assign popcount21_ltw2_core_139 = ~(input_a[12] ^ input_a[19]);
  assign popcount21_ltw2_core_140 = input_a[9] ^ input_a[16];
  assign popcount21_ltw2_core_141_not = ~input_a[5];
  assign popcount21_ltw2_core_144 = ~input_a[19];
  assign popcount21_ltw2_core_145 = input_a[12] | input_a[12];
  assign popcount21_ltw2_core_149 = input_a[6] | input_a[14];

  assign popcount21_ltw2_out[0] = input_a[6];
  assign popcount21_ltw2_out[1] = input_a[16];
  assign popcount21_ltw2_out[2] = 1'b1;
  assign popcount21_ltw2_out[3] = input_a[19];
  assign popcount21_ltw2_out[4] = input_a[1];
endmodule