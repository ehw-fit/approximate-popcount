// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.52929
// WCE=14.0
// EP=0.877786%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_qgj4(input [23:0] input_a, output [4:0] popcount24_qgj4_out);
  wire popcount24_qgj4_core_028;
  wire popcount24_qgj4_core_029;
  wire popcount24_qgj4_core_030;
  wire popcount24_qgj4_core_032;
  wire popcount24_qgj4_core_034;
  wire popcount24_qgj4_core_035;
  wire popcount24_qgj4_core_036;
  wire popcount24_qgj4_core_038;
  wire popcount24_qgj4_core_040;
  wire popcount24_qgj4_core_041;
  wire popcount24_qgj4_core_045;
  wire popcount24_qgj4_core_046;
  wire popcount24_qgj4_core_047;
  wire popcount24_qgj4_core_049;
  wire popcount24_qgj4_core_051;
  wire popcount24_qgj4_core_052;
  wire popcount24_qgj4_core_053_not;
  wire popcount24_qgj4_core_054;
  wire popcount24_qgj4_core_055;
  wire popcount24_qgj4_core_056;
  wire popcount24_qgj4_core_058;
  wire popcount24_qgj4_core_059;
  wire popcount24_qgj4_core_060;
  wire popcount24_qgj4_core_062;
  wire popcount24_qgj4_core_063;
  wire popcount24_qgj4_core_066;
  wire popcount24_qgj4_core_067;
  wire popcount24_qgj4_core_068;
  wire popcount24_qgj4_core_071;
  wire popcount24_qgj4_core_072;
  wire popcount24_qgj4_core_073;
  wire popcount24_qgj4_core_074;
  wire popcount24_qgj4_core_076;
  wire popcount24_qgj4_core_077;
  wire popcount24_qgj4_core_078;
  wire popcount24_qgj4_core_081;
  wire popcount24_qgj4_core_083;
  wire popcount24_qgj4_core_084;
  wire popcount24_qgj4_core_086;
  wire popcount24_qgj4_core_088;
  wire popcount24_qgj4_core_090;
  wire popcount24_qgj4_core_092;
  wire popcount24_qgj4_core_093;
  wire popcount24_qgj4_core_095;
  wire popcount24_qgj4_core_096;
  wire popcount24_qgj4_core_097;
  wire popcount24_qgj4_core_098;
  wire popcount24_qgj4_core_100;
  wire popcount24_qgj4_core_101;
  wire popcount24_qgj4_core_102;
  wire popcount24_qgj4_core_103;
  wire popcount24_qgj4_core_105;
  wire popcount24_qgj4_core_106;
  wire popcount24_qgj4_core_107;
  wire popcount24_qgj4_core_108;
  wire popcount24_qgj4_core_112;
  wire popcount24_qgj4_core_113;
  wire popcount24_qgj4_core_114;
  wire popcount24_qgj4_core_116;
  wire popcount24_qgj4_core_117;
  wire popcount24_qgj4_core_118;
  wire popcount24_qgj4_core_120;
  wire popcount24_qgj4_core_122;
  wire popcount24_qgj4_core_123;
  wire popcount24_qgj4_core_125;
  wire popcount24_qgj4_core_126;
  wire popcount24_qgj4_core_128;
  wire popcount24_qgj4_core_129_not;
  wire popcount24_qgj4_core_131;
  wire popcount24_qgj4_core_133;
  wire popcount24_qgj4_core_134;
  wire popcount24_qgj4_core_135;
  wire popcount24_qgj4_core_136;
  wire popcount24_qgj4_core_138;
  wire popcount24_qgj4_core_139;
  wire popcount24_qgj4_core_140;
  wire popcount24_qgj4_core_142;
  wire popcount24_qgj4_core_143;
  wire popcount24_qgj4_core_144;
  wire popcount24_qgj4_core_146;
  wire popcount24_qgj4_core_147;
  wire popcount24_qgj4_core_148;
  wire popcount24_qgj4_core_149;
  wire popcount24_qgj4_core_150;
  wire popcount24_qgj4_core_151_not;
  wire popcount24_qgj4_core_153;
  wire popcount24_qgj4_core_155;
  wire popcount24_qgj4_core_158;
  wire popcount24_qgj4_core_159;
  wire popcount24_qgj4_core_162;
  wire popcount24_qgj4_core_163;
  wire popcount24_qgj4_core_164;
  wire popcount24_qgj4_core_166;
  wire popcount24_qgj4_core_167;
  wire popcount24_qgj4_core_171;
  wire popcount24_qgj4_core_172;
  wire popcount24_qgj4_core_173;
  wire popcount24_qgj4_core_174;
  wire popcount24_qgj4_core_175;

  assign popcount24_qgj4_core_028 = ~input_a[16];
  assign popcount24_qgj4_core_029 = ~(input_a[9] | input_a[8]);
  assign popcount24_qgj4_core_030 = input_a[11] ^ input_a[18];
  assign popcount24_qgj4_core_032 = ~(input_a[1] & input_a[6]);
  assign popcount24_qgj4_core_034 = ~(input_a[5] ^ input_a[20]);
  assign popcount24_qgj4_core_035 = ~input_a[6];
  assign popcount24_qgj4_core_036 = input_a[21] & input_a[16];
  assign popcount24_qgj4_core_038 = ~(input_a[8] ^ input_a[8]);
  assign popcount24_qgj4_core_040 = ~(input_a[1] & input_a[11]);
  assign popcount24_qgj4_core_041 = ~(input_a[14] | input_a[19]);
  assign popcount24_qgj4_core_045 = ~input_a[3];
  assign popcount24_qgj4_core_046 = input_a[0] & input_a[12];
  assign popcount24_qgj4_core_047 = input_a[22] & input_a[23];
  assign popcount24_qgj4_core_049 = input_a[23] ^ input_a[6];
  assign popcount24_qgj4_core_051 = input_a[2] | input_a[7];
  assign popcount24_qgj4_core_052 = input_a[20] | input_a[15];
  assign popcount24_qgj4_core_053_not = ~input_a[12];
  assign popcount24_qgj4_core_054 = input_a[11] ^ input_a[19];
  assign popcount24_qgj4_core_055 = ~(input_a[10] ^ input_a[13]);
  assign popcount24_qgj4_core_056 = input_a[16] ^ input_a[13];
  assign popcount24_qgj4_core_058 = input_a[13] | input_a[19];
  assign popcount24_qgj4_core_059 = input_a[1] ^ input_a[7];
  assign popcount24_qgj4_core_060 = ~input_a[9];
  assign popcount24_qgj4_core_062 = input_a[23] ^ input_a[5];
  assign popcount24_qgj4_core_063 = ~(input_a[15] ^ input_a[19]);
  assign popcount24_qgj4_core_066 = ~(input_a[11] | input_a[1]);
  assign popcount24_qgj4_core_067 = input_a[16] ^ input_a[9];
  assign popcount24_qgj4_core_068 = ~(input_a[1] & input_a[11]);
  assign popcount24_qgj4_core_071 = input_a[4] ^ input_a[20];
  assign popcount24_qgj4_core_072 = ~(input_a[4] & input_a[5]);
  assign popcount24_qgj4_core_073 = input_a[23] ^ input_a[19];
  assign popcount24_qgj4_core_074 = ~(input_a[14] & input_a[8]);
  assign popcount24_qgj4_core_076 = ~(input_a[4] ^ input_a[14]);
  assign popcount24_qgj4_core_077 = input_a[7] ^ input_a[18];
  assign popcount24_qgj4_core_078 = ~(input_a[3] & input_a[13]);
  assign popcount24_qgj4_core_081 = input_a[19] | input_a[20];
  assign popcount24_qgj4_core_083 = input_a[22] ^ input_a[18];
  assign popcount24_qgj4_core_084 = ~(input_a[3] ^ input_a[6]);
  assign popcount24_qgj4_core_086 = input_a[4] & input_a[20];
  assign popcount24_qgj4_core_088 = ~(input_a[11] & input_a[4]);
  assign popcount24_qgj4_core_090 = input_a[16] & input_a[9];
  assign popcount24_qgj4_core_092 = input_a[5] ^ input_a[21];
  assign popcount24_qgj4_core_093 = input_a[13] | input_a[6];
  assign popcount24_qgj4_core_095 = input_a[22] ^ input_a[22];
  assign popcount24_qgj4_core_096 = ~(input_a[18] & input_a[23]);
  assign popcount24_qgj4_core_097 = ~input_a[11];
  assign popcount24_qgj4_core_098 = ~input_a[16];
  assign popcount24_qgj4_core_100 = input_a[23] ^ input_a[8];
  assign popcount24_qgj4_core_101 = input_a[7] | input_a[12];
  assign popcount24_qgj4_core_102 = ~(input_a[22] ^ input_a[2]);
  assign popcount24_qgj4_core_103 = ~(input_a[5] & input_a[19]);
  assign popcount24_qgj4_core_105 = input_a[13] & input_a[7];
  assign popcount24_qgj4_core_106 = ~input_a[16];
  assign popcount24_qgj4_core_107 = input_a[13] | input_a[13];
  assign popcount24_qgj4_core_108 = input_a[21] | input_a[9];
  assign popcount24_qgj4_core_112 = input_a[6] & input_a[17];
  assign popcount24_qgj4_core_113 = input_a[9] & input_a[4];
  assign popcount24_qgj4_core_114 = ~(input_a[10] | input_a[20]);
  assign popcount24_qgj4_core_116 = input_a[21] & input_a[11];
  assign popcount24_qgj4_core_117 = ~input_a[1];
  assign popcount24_qgj4_core_118 = ~(input_a[8] ^ input_a[4]);
  assign popcount24_qgj4_core_120 = input_a[6] & input_a[6];
  assign popcount24_qgj4_core_122 = input_a[6] & input_a[17];
  assign popcount24_qgj4_core_123 = input_a[4] ^ input_a[7];
  assign popcount24_qgj4_core_125 = input_a[13] & input_a[16];
  assign popcount24_qgj4_core_126 = input_a[10] ^ input_a[19];
  assign popcount24_qgj4_core_128 = input_a[12] ^ input_a[12];
  assign popcount24_qgj4_core_129_not = ~input_a[6];
  assign popcount24_qgj4_core_131 = input_a[0] ^ input_a[13];
  assign popcount24_qgj4_core_133 = input_a[16] & input_a[8];
  assign popcount24_qgj4_core_134 = ~(input_a[2] & input_a[16]);
  assign popcount24_qgj4_core_135 = ~input_a[2];
  assign popcount24_qgj4_core_136 = input_a[20] ^ input_a[14];
  assign popcount24_qgj4_core_138 = input_a[16] ^ input_a[3];
  assign popcount24_qgj4_core_139 = input_a[10] & input_a[8];
  assign popcount24_qgj4_core_140 = input_a[12] & input_a[16];
  assign popcount24_qgj4_core_142 = input_a[12] | input_a[2];
  assign popcount24_qgj4_core_143 = input_a[13] & input_a[9];
  assign popcount24_qgj4_core_144 = ~(input_a[16] ^ input_a[5]);
  assign popcount24_qgj4_core_146 = input_a[3] & input_a[10];
  assign popcount24_qgj4_core_147 = input_a[17] | input_a[1];
  assign popcount24_qgj4_core_148 = ~input_a[0];
  assign popcount24_qgj4_core_149 = input_a[20] ^ input_a[7];
  assign popcount24_qgj4_core_150 = input_a[13] ^ input_a[19];
  assign popcount24_qgj4_core_151_not = ~input_a[14];
  assign popcount24_qgj4_core_153 = ~(input_a[0] ^ input_a[3]);
  assign popcount24_qgj4_core_155 = ~(input_a[23] | input_a[17]);
  assign popcount24_qgj4_core_158 = ~input_a[2];
  assign popcount24_qgj4_core_159 = ~input_a[10];
  assign popcount24_qgj4_core_162 = input_a[21] ^ input_a[9];
  assign popcount24_qgj4_core_163 = ~(input_a[20] | input_a[14]);
  assign popcount24_qgj4_core_164 = input_a[2] ^ input_a[19];
  assign popcount24_qgj4_core_166 = ~(input_a[23] ^ input_a[18]);
  assign popcount24_qgj4_core_167 = ~(input_a[15] ^ input_a[1]);
  assign popcount24_qgj4_core_171 = ~(input_a[8] ^ input_a[20]);
  assign popcount24_qgj4_core_172 = ~(input_a[22] | input_a[18]);
  assign popcount24_qgj4_core_173 = ~input_a[19];
  assign popcount24_qgj4_core_174 = ~input_a[6];
  assign popcount24_qgj4_core_175 = ~(input_a[1] | input_a[12]);

  assign popcount24_qgj4_out[0] = input_a[22];
  assign popcount24_qgj4_out[1] = 1'b0;
  assign popcount24_qgj4_out[2] = input_a[18];
  assign popcount24_qgj4_out[3] = 1'b1;
  assign popcount24_qgj4_out[4] = 1'b0;
endmodule