// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.12191
// WCE=21.0
// EP=0.963781%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_wicn(input [29:0] input_a, output [4:0] popcount30_wicn_out);
  wire popcount30_wicn_core_032;
  wire popcount30_wicn_core_034;
  wire popcount30_wicn_core_035;
  wire popcount30_wicn_core_038;
  wire popcount30_wicn_core_039;
  wire popcount30_wicn_core_040;
  wire popcount30_wicn_core_041;
  wire popcount30_wicn_core_042;
  wire popcount30_wicn_core_043;
  wire popcount30_wicn_core_044;
  wire popcount30_wicn_core_045;
  wire popcount30_wicn_core_046;
  wire popcount30_wicn_core_047;
  wire popcount30_wicn_core_048;
  wire popcount30_wicn_core_049;
  wire popcount30_wicn_core_052;
  wire popcount30_wicn_core_053;
  wire popcount30_wicn_core_055;
  wire popcount30_wicn_core_058;
  wire popcount30_wicn_core_061;
  wire popcount30_wicn_core_062;
  wire popcount30_wicn_core_064;
  wire popcount30_wicn_core_065;
  wire popcount30_wicn_core_068;
  wire popcount30_wicn_core_069;
  wire popcount30_wicn_core_071;
  wire popcount30_wicn_core_072;
  wire popcount30_wicn_core_073;
  wire popcount30_wicn_core_074;
  wire popcount30_wicn_core_076;
  wire popcount30_wicn_core_077;
  wire popcount30_wicn_core_078;
  wire popcount30_wicn_core_079;
  wire popcount30_wicn_core_080;
  wire popcount30_wicn_core_081;
  wire popcount30_wicn_core_082;
  wire popcount30_wicn_core_083;
  wire popcount30_wicn_core_084;
  wire popcount30_wicn_core_087;
  wire popcount30_wicn_core_089;
  wire popcount30_wicn_core_090;
  wire popcount30_wicn_core_091;
  wire popcount30_wicn_core_092;
  wire popcount30_wicn_core_093;
  wire popcount30_wicn_core_097;
  wire popcount30_wicn_core_098;
  wire popcount30_wicn_core_099;
  wire popcount30_wicn_core_100;
  wire popcount30_wicn_core_101;
  wire popcount30_wicn_core_102;
  wire popcount30_wicn_core_103;
  wire popcount30_wicn_core_104;
  wire popcount30_wicn_core_105;
  wire popcount30_wicn_core_106;
  wire popcount30_wicn_core_108;
  wire popcount30_wicn_core_111;
  wire popcount30_wicn_core_113;
  wire popcount30_wicn_core_115;
  wire popcount30_wicn_core_117;
  wire popcount30_wicn_core_118;
  wire popcount30_wicn_core_121;
  wire popcount30_wicn_core_122;
  wire popcount30_wicn_core_123;
  wire popcount30_wicn_core_124;
  wire popcount30_wicn_core_125;
  wire popcount30_wicn_core_126_not;
  wire popcount30_wicn_core_127;
  wire popcount30_wicn_core_134;
  wire popcount30_wicn_core_137;
  wire popcount30_wicn_core_139;
  wire popcount30_wicn_core_140;
  wire popcount30_wicn_core_142;
  wire popcount30_wicn_core_143;
  wire popcount30_wicn_core_144;
  wire popcount30_wicn_core_145;
  wire popcount30_wicn_core_146;
  wire popcount30_wicn_core_149;
  wire popcount30_wicn_core_151;
  wire popcount30_wicn_core_152_not;
  wire popcount30_wicn_core_153;
  wire popcount30_wicn_core_154;
  wire popcount30_wicn_core_161;
  wire popcount30_wicn_core_162;
  wire popcount30_wicn_core_164;
  wire popcount30_wicn_core_165;
  wire popcount30_wicn_core_167;
  wire popcount30_wicn_core_168;
  wire popcount30_wicn_core_169;
  wire popcount30_wicn_core_172;
  wire popcount30_wicn_core_173;
  wire popcount30_wicn_core_175;
  wire popcount30_wicn_core_176;
  wire popcount30_wicn_core_177;
  wire popcount30_wicn_core_178;
  wire popcount30_wicn_core_179;
  wire popcount30_wicn_core_182;
  wire popcount30_wicn_core_183;
  wire popcount30_wicn_core_184;
  wire popcount30_wicn_core_185;
  wire popcount30_wicn_core_186;
  wire popcount30_wicn_core_187;
  wire popcount30_wicn_core_188;
  wire popcount30_wicn_core_191;
  wire popcount30_wicn_core_192;
  wire popcount30_wicn_core_194;
  wire popcount30_wicn_core_195;
  wire popcount30_wicn_core_196;
  wire popcount30_wicn_core_197;
  wire popcount30_wicn_core_198;
  wire popcount30_wicn_core_200;
  wire popcount30_wicn_core_201;
  wire popcount30_wicn_core_203;
  wire popcount30_wicn_core_204;
  wire popcount30_wicn_core_208;
  wire popcount30_wicn_core_209;
  wire popcount30_wicn_core_211;
  wire popcount30_wicn_core_212;
  wire popcount30_wicn_core_213;

  assign popcount30_wicn_core_032 = ~(input_a[7] | input_a[0]);
  assign popcount30_wicn_core_034 = input_a[21] & input_a[20];
  assign popcount30_wicn_core_035 = ~(input_a[28] | input_a[1]);
  assign popcount30_wicn_core_038 = ~(input_a[23] & input_a[5]);
  assign popcount30_wicn_core_039 = input_a[14] & input_a[26];
  assign popcount30_wicn_core_040 = input_a[7] | input_a[5];
  assign popcount30_wicn_core_041 = input_a[20] | input_a[20];
  assign popcount30_wicn_core_042 = input_a[25] ^ input_a[7];
  assign popcount30_wicn_core_043 = ~(input_a[15] | input_a[6]);
  assign popcount30_wicn_core_044 = input_a[7] ^ input_a[19];
  assign popcount30_wicn_core_045 = ~(input_a[15] ^ input_a[0]);
  assign popcount30_wicn_core_046 = input_a[0] | input_a[26];
  assign popcount30_wicn_core_047 = ~(input_a[19] ^ input_a[20]);
  assign popcount30_wicn_core_048 = ~input_a[25];
  assign popcount30_wicn_core_049 = ~(input_a[28] & input_a[18]);
  assign popcount30_wicn_core_052 = ~(input_a[1] & input_a[28]);
  assign popcount30_wicn_core_053 = input_a[29] | input_a[5];
  assign popcount30_wicn_core_055 = ~input_a[20];
  assign popcount30_wicn_core_058 = ~(input_a[13] ^ input_a[1]);
  assign popcount30_wicn_core_061 = input_a[14] ^ input_a[15];
  assign popcount30_wicn_core_062 = input_a[27] | input_a[4];
  assign popcount30_wicn_core_064 = ~(input_a[4] | input_a[21]);
  assign popcount30_wicn_core_065 = ~(input_a[28] | input_a[2]);
  assign popcount30_wicn_core_068 = input_a[15] ^ input_a[20];
  assign popcount30_wicn_core_069 = ~(input_a[16] & input_a[14]);
  assign popcount30_wicn_core_071 = input_a[27] ^ input_a[16];
  assign popcount30_wicn_core_072 = ~(input_a[1] & input_a[14]);
  assign popcount30_wicn_core_073 = ~(input_a[13] & input_a[12]);
  assign popcount30_wicn_core_074 = ~input_a[17];
  assign popcount30_wicn_core_076 = ~(input_a[29] ^ input_a[16]);
  assign popcount30_wicn_core_077 = ~(input_a[20] | input_a[6]);
  assign popcount30_wicn_core_078 = ~(input_a[15] ^ input_a[10]);
  assign popcount30_wicn_core_079 = ~input_a[8];
  assign popcount30_wicn_core_080 = input_a[16] | input_a[26];
  assign popcount30_wicn_core_081 = ~(input_a[6] ^ input_a[4]);
  assign popcount30_wicn_core_082 = ~(input_a[12] & input_a[24]);
  assign popcount30_wicn_core_083 = ~input_a[6];
  assign popcount30_wicn_core_084 = input_a[13] | input_a[3];
  assign popcount30_wicn_core_087 = ~(input_a[12] ^ input_a[15]);
  assign popcount30_wicn_core_089 = input_a[27] | input_a[10];
  assign popcount30_wicn_core_090 = ~(input_a[8] ^ input_a[28]);
  assign popcount30_wicn_core_091 = input_a[23] ^ input_a[4];
  assign popcount30_wicn_core_092 = ~input_a[19];
  assign popcount30_wicn_core_093 = input_a[9] & input_a[11];
  assign popcount30_wicn_core_097 = ~(input_a[9] & input_a[22]);
  assign popcount30_wicn_core_098 = ~(input_a[3] ^ input_a[25]);
  assign popcount30_wicn_core_099 = ~(input_a[19] | input_a[27]);
  assign popcount30_wicn_core_100 = input_a[13] & input_a[7];
  assign popcount30_wicn_core_101 = ~input_a[1];
  assign popcount30_wicn_core_102 = input_a[25] & input_a[23];
  assign popcount30_wicn_core_103 = input_a[20] | input_a[9];
  assign popcount30_wicn_core_104 = input_a[29] & input_a[6];
  assign popcount30_wicn_core_105 = ~input_a[21];
  assign popcount30_wicn_core_106 = ~(input_a[0] | input_a[23]);
  assign popcount30_wicn_core_108 = ~(input_a[4] | input_a[17]);
  assign popcount30_wicn_core_111 = input_a[6] ^ input_a[24];
  assign popcount30_wicn_core_113 = ~(input_a[18] & input_a[27]);
  assign popcount30_wicn_core_115 = ~(input_a[15] & input_a[8]);
  assign popcount30_wicn_core_117 = input_a[20] ^ input_a[8];
  assign popcount30_wicn_core_118 = input_a[12] | input_a[11];
  assign popcount30_wicn_core_121 = ~(input_a[21] | input_a[16]);
  assign popcount30_wicn_core_122 = input_a[24] ^ input_a[28];
  assign popcount30_wicn_core_123 = input_a[23] & input_a[22];
  assign popcount30_wicn_core_124 = input_a[20] & input_a[9];
  assign popcount30_wicn_core_125 = input_a[11] & input_a[24];
  assign popcount30_wicn_core_126_not = ~input_a[10];
  assign popcount30_wicn_core_127 = ~input_a[7];
  assign popcount30_wicn_core_134 = ~(input_a[5] & input_a[9]);
  assign popcount30_wicn_core_137 = input_a[14] & input_a[1];
  assign popcount30_wicn_core_139 = ~(input_a[21] ^ input_a[26]);
  assign popcount30_wicn_core_140 = input_a[2] & input_a[16];
  assign popcount30_wicn_core_142 = ~(input_a[4] ^ input_a[6]);
  assign popcount30_wicn_core_143 = input_a[14] ^ input_a[2];
  assign popcount30_wicn_core_144 = input_a[27] ^ input_a[29];
  assign popcount30_wicn_core_145 = ~(input_a[10] ^ input_a[13]);
  assign popcount30_wicn_core_146 = ~(input_a[10] | input_a[11]);
  assign popcount30_wicn_core_149 = ~(input_a[11] | input_a[7]);
  assign popcount30_wicn_core_151 = ~(input_a[16] & input_a[23]);
  assign popcount30_wicn_core_152_not = ~input_a[7];
  assign popcount30_wicn_core_153 = input_a[1] | input_a[21];
  assign popcount30_wicn_core_154 = ~input_a[6];
  assign popcount30_wicn_core_161 = input_a[6] | input_a[29];
  assign popcount30_wicn_core_162 = ~(input_a[23] & input_a[15]);
  assign popcount30_wicn_core_164 = input_a[8] ^ input_a[19];
  assign popcount30_wicn_core_165 = ~(input_a[8] | input_a[2]);
  assign popcount30_wicn_core_167 = input_a[9] ^ input_a[29];
  assign popcount30_wicn_core_168 = ~(input_a[6] ^ input_a[1]);
  assign popcount30_wicn_core_169 = input_a[26] & input_a[19];
  assign popcount30_wicn_core_172 = ~(input_a[15] ^ input_a[10]);
  assign popcount30_wicn_core_173 = ~input_a[17];
  assign popcount30_wicn_core_175 = ~(input_a[1] & input_a[23]);
  assign popcount30_wicn_core_176 = ~(input_a[5] ^ input_a[23]);
  assign popcount30_wicn_core_177 = ~input_a[3];
  assign popcount30_wicn_core_178 = ~(input_a[10] & input_a[20]);
  assign popcount30_wicn_core_179 = ~input_a[6];
  assign popcount30_wicn_core_182 = input_a[20] | input_a[4];
  assign popcount30_wicn_core_183 = input_a[20] & input_a[14];
  assign popcount30_wicn_core_184 = ~input_a[29];
  assign popcount30_wicn_core_185 = ~input_a[29];
  assign popcount30_wicn_core_186 = ~input_a[11];
  assign popcount30_wicn_core_187 = input_a[6] ^ input_a[20];
  assign popcount30_wicn_core_188 = ~(input_a[6] & input_a[13]);
  assign popcount30_wicn_core_191 = ~(input_a[2] & input_a[12]);
  assign popcount30_wicn_core_192 = input_a[4] & input_a[2];
  assign popcount30_wicn_core_194 = ~(input_a[12] ^ input_a[2]);
  assign popcount30_wicn_core_195 = input_a[25] | input_a[9];
  assign popcount30_wicn_core_196 = ~(input_a[7] | input_a[26]);
  assign popcount30_wicn_core_197 = ~(input_a[2] | input_a[27]);
  assign popcount30_wicn_core_198 = input_a[2] & input_a[13];
  assign popcount30_wicn_core_200 = ~(input_a[17] ^ input_a[18]);
  assign popcount30_wicn_core_201 = ~(input_a[0] | input_a[6]);
  assign popcount30_wicn_core_203 = ~(input_a[12] & input_a[29]);
  assign popcount30_wicn_core_204 = ~(input_a[24] ^ input_a[27]);
  assign popcount30_wicn_core_208 = ~input_a[6];
  assign popcount30_wicn_core_209 = ~input_a[26];
  assign popcount30_wicn_core_211 = input_a[8] | input_a[18];
  assign popcount30_wicn_core_212 = input_a[27] & input_a[15];
  assign popcount30_wicn_core_213 = ~(input_a[26] ^ input_a[9]);

  assign popcount30_wicn_out[0] = 1'b0;
  assign popcount30_wicn_out[1] = 1'b0;
  assign popcount30_wicn_out[2] = input_a[4];
  assign popcount30_wicn_out[3] = 1'b1;
  assign popcount30_wicn_out[4] = 1'b0;
endmodule