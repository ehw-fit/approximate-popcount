// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.64769
// WCE=28.0
// EP=0.970739%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_bqn3(input [32:0] input_a, output [5:0] popcount33_bqn3_out);
  wire popcount33_bqn3_core_036;
  wire popcount33_bqn3_core_039;
  wire popcount33_bqn3_core_041;
  wire popcount33_bqn3_core_045;
  wire popcount33_bqn3_core_046;
  wire popcount33_bqn3_core_047;
  wire popcount33_bqn3_core_048;
  wire popcount33_bqn3_core_049;
  wire popcount33_bqn3_core_050;
  wire popcount33_bqn3_core_051;
  wire popcount33_bqn3_core_053;
  wire popcount33_bqn3_core_055;
  wire popcount33_bqn3_core_056;
  wire popcount33_bqn3_core_058;
  wire popcount33_bqn3_core_059;
  wire popcount33_bqn3_core_060;
  wire popcount33_bqn3_core_061;
  wire popcount33_bqn3_core_062;
  wire popcount33_bqn3_core_065;
  wire popcount33_bqn3_core_068;
  wire popcount33_bqn3_core_069;
  wire popcount33_bqn3_core_071;
  wire popcount33_bqn3_core_072;
  wire popcount33_bqn3_core_073;
  wire popcount33_bqn3_core_074;
  wire popcount33_bqn3_core_076;
  wire popcount33_bqn3_core_077;
  wire popcount33_bqn3_core_079;
  wire popcount33_bqn3_core_080;
  wire popcount33_bqn3_core_081;
  wire popcount33_bqn3_core_082;
  wire popcount33_bqn3_core_084;
  wire popcount33_bqn3_core_085;
  wire popcount33_bqn3_core_087;
  wire popcount33_bqn3_core_088;
  wire popcount33_bqn3_core_089;
  wire popcount33_bqn3_core_090;
  wire popcount33_bqn3_core_091;
  wire popcount33_bqn3_core_092;
  wire popcount33_bqn3_core_095;
  wire popcount33_bqn3_core_098;
  wire popcount33_bqn3_core_099;
  wire popcount33_bqn3_core_100;
  wire popcount33_bqn3_core_101;
  wire popcount33_bqn3_core_102;
  wire popcount33_bqn3_core_105;
  wire popcount33_bqn3_core_106;
  wire popcount33_bqn3_core_107;
  wire popcount33_bqn3_core_111;
  wire popcount33_bqn3_core_117;
  wire popcount33_bqn3_core_118;
  wire popcount33_bqn3_core_119;
  wire popcount33_bqn3_core_120;
  wire popcount33_bqn3_core_121;
  wire popcount33_bqn3_core_122;
  wire popcount33_bqn3_core_124_not;
  wire popcount33_bqn3_core_126;
  wire popcount33_bqn3_core_127;
  wire popcount33_bqn3_core_128;
  wire popcount33_bqn3_core_130;
  wire popcount33_bqn3_core_131;
  wire popcount33_bqn3_core_132;
  wire popcount33_bqn3_core_134;
  wire popcount33_bqn3_core_135;
  wire popcount33_bqn3_core_136;
  wire popcount33_bqn3_core_137;
  wire popcount33_bqn3_core_139;
  wire popcount33_bqn3_core_141;
  wire popcount33_bqn3_core_142;
  wire popcount33_bqn3_core_144;
  wire popcount33_bqn3_core_145_not;
  wire popcount33_bqn3_core_146;
  wire popcount33_bqn3_core_147_not;
  wire popcount33_bqn3_core_150;
  wire popcount33_bqn3_core_151;
  wire popcount33_bqn3_core_154;
  wire popcount33_bqn3_core_157;
  wire popcount33_bqn3_core_160;
  wire popcount33_bqn3_core_161;
  wire popcount33_bqn3_core_163;
  wire popcount33_bqn3_core_165;
  wire popcount33_bqn3_core_166;
  wire popcount33_bqn3_core_169;
  wire popcount33_bqn3_core_170;
  wire popcount33_bqn3_core_171;
  wire popcount33_bqn3_core_172;
  wire popcount33_bqn3_core_173;
  wire popcount33_bqn3_core_174;
  wire popcount33_bqn3_core_179;
  wire popcount33_bqn3_core_180;
  wire popcount33_bqn3_core_181;
  wire popcount33_bqn3_core_184;
  wire popcount33_bqn3_core_186;
  wire popcount33_bqn3_core_188;
  wire popcount33_bqn3_core_191;
  wire popcount33_bqn3_core_192;
  wire popcount33_bqn3_core_193;
  wire popcount33_bqn3_core_194;
  wire popcount33_bqn3_core_198;
  wire popcount33_bqn3_core_199_not;
  wire popcount33_bqn3_core_200;
  wire popcount33_bqn3_core_201;
  wire popcount33_bqn3_core_203;
  wire popcount33_bqn3_core_204;
  wire popcount33_bqn3_core_205_not;
  wire popcount33_bqn3_core_206;
  wire popcount33_bqn3_core_207;
  wire popcount33_bqn3_core_208;
  wire popcount33_bqn3_core_209;
  wire popcount33_bqn3_core_211;
  wire popcount33_bqn3_core_212;
  wire popcount33_bqn3_core_213_not;
  wire popcount33_bqn3_core_215;
  wire popcount33_bqn3_core_216;
  wire popcount33_bqn3_core_219;
  wire popcount33_bqn3_core_220;
  wire popcount33_bqn3_core_223;
  wire popcount33_bqn3_core_224;
  wire popcount33_bqn3_core_225;
  wire popcount33_bqn3_core_226;
  wire popcount33_bqn3_core_227;
  wire popcount33_bqn3_core_228;
  wire popcount33_bqn3_core_230;
  wire popcount33_bqn3_core_232;
  wire popcount33_bqn3_core_233;
  wire popcount33_bqn3_core_234;
  wire popcount33_bqn3_core_235;
  wire popcount33_bqn3_core_236;
  wire popcount33_bqn3_core_238;

  assign popcount33_bqn3_core_036 = ~(input_a[20] ^ input_a[15]);
  assign popcount33_bqn3_core_039 = ~(input_a[16] ^ input_a[4]);
  assign popcount33_bqn3_core_041 = input_a[30] & input_a[10];
  assign popcount33_bqn3_core_045 = ~(input_a[16] ^ input_a[13]);
  assign popcount33_bqn3_core_046 = input_a[13] | input_a[8];
  assign popcount33_bqn3_core_047 = input_a[26] ^ input_a[28];
  assign popcount33_bqn3_core_048 = ~input_a[17];
  assign popcount33_bqn3_core_049 = input_a[18] ^ input_a[1];
  assign popcount33_bqn3_core_050 = ~input_a[5];
  assign popcount33_bqn3_core_051 = input_a[18] ^ input_a[1];
  assign popcount33_bqn3_core_053 = input_a[20] & input_a[5];
  assign popcount33_bqn3_core_055 = ~(input_a[30] ^ input_a[30]);
  assign popcount33_bqn3_core_056 = ~(input_a[11] | input_a[1]);
  assign popcount33_bqn3_core_058 = input_a[2] ^ input_a[30];
  assign popcount33_bqn3_core_059 = ~(input_a[19] | input_a[16]);
  assign popcount33_bqn3_core_060 = ~(input_a[26] & input_a[4]);
  assign popcount33_bqn3_core_061 = ~input_a[31];
  assign popcount33_bqn3_core_062 = ~(input_a[12] ^ input_a[28]);
  assign popcount33_bqn3_core_065 = ~input_a[14];
  assign popcount33_bqn3_core_068 = input_a[18] & input_a[4];
  assign popcount33_bqn3_core_069 = input_a[9] ^ input_a[16];
  assign popcount33_bqn3_core_071 = ~(input_a[16] ^ input_a[6]);
  assign popcount33_bqn3_core_072 = ~(input_a[14] ^ input_a[15]);
  assign popcount33_bqn3_core_073 = input_a[28] | input_a[13];
  assign popcount33_bqn3_core_074 = ~(input_a[32] ^ input_a[3]);
  assign popcount33_bqn3_core_076 = input_a[9] & input_a[6];
  assign popcount33_bqn3_core_077 = ~(input_a[11] ^ input_a[2]);
  assign popcount33_bqn3_core_079 = input_a[11] & input_a[11];
  assign popcount33_bqn3_core_080 = ~(input_a[15] | input_a[22]);
  assign popcount33_bqn3_core_081 = ~(input_a[30] & input_a[23]);
  assign popcount33_bqn3_core_082 = ~(input_a[3] & input_a[11]);
  assign popcount33_bqn3_core_084 = ~(input_a[25] | input_a[22]);
  assign popcount33_bqn3_core_085 = ~(input_a[11] | input_a[18]);
  assign popcount33_bqn3_core_087 = ~(input_a[17] ^ input_a[14]);
  assign popcount33_bqn3_core_088 = ~(input_a[32] ^ input_a[14]);
  assign popcount33_bqn3_core_089 = ~(input_a[27] & input_a[30]);
  assign popcount33_bqn3_core_090 = input_a[25] ^ input_a[9];
  assign popcount33_bqn3_core_091 = ~(input_a[13] & input_a[20]);
  assign popcount33_bqn3_core_092 = input_a[15] ^ input_a[20];
  assign popcount33_bqn3_core_095 = input_a[30] & input_a[18];
  assign popcount33_bqn3_core_098 = ~input_a[10];
  assign popcount33_bqn3_core_099 = ~(input_a[28] | input_a[4]);
  assign popcount33_bqn3_core_100 = ~(input_a[22] ^ input_a[3]);
  assign popcount33_bqn3_core_101 = ~(input_a[11] & input_a[27]);
  assign popcount33_bqn3_core_102 = input_a[7] ^ input_a[9];
  assign popcount33_bqn3_core_105 = ~input_a[28];
  assign popcount33_bqn3_core_106 = ~(input_a[8] ^ input_a[11]);
  assign popcount33_bqn3_core_107 = input_a[32] & input_a[27];
  assign popcount33_bqn3_core_111 = input_a[18] ^ input_a[7];
  assign popcount33_bqn3_core_117 = ~(input_a[17] & input_a[23]);
  assign popcount33_bqn3_core_118 = input_a[12] | input_a[8];
  assign popcount33_bqn3_core_119 = ~input_a[23];
  assign popcount33_bqn3_core_120 = ~(input_a[28] | input_a[0]);
  assign popcount33_bqn3_core_121 = input_a[14] ^ input_a[9];
  assign popcount33_bqn3_core_122 = ~(input_a[5] & input_a[30]);
  assign popcount33_bqn3_core_124_not = ~input_a[1];
  assign popcount33_bqn3_core_126 = ~(input_a[27] | input_a[29]);
  assign popcount33_bqn3_core_127 = ~(input_a[13] & input_a[2]);
  assign popcount33_bqn3_core_128 = ~input_a[17];
  assign popcount33_bqn3_core_130 = ~(input_a[11] & input_a[23]);
  assign popcount33_bqn3_core_131 = ~(input_a[1] ^ input_a[16]);
  assign popcount33_bqn3_core_132 = ~(input_a[30] ^ input_a[4]);
  assign popcount33_bqn3_core_134 = ~(input_a[24] ^ input_a[0]);
  assign popcount33_bqn3_core_135 = input_a[21] & input_a[19];
  assign popcount33_bqn3_core_136 = input_a[14] & input_a[25];
  assign popcount33_bqn3_core_137 = input_a[13] | input_a[17];
  assign popcount33_bqn3_core_139 = ~(input_a[2] | input_a[19]);
  assign popcount33_bqn3_core_141 = ~input_a[2];
  assign popcount33_bqn3_core_142 = ~input_a[8];
  assign popcount33_bqn3_core_144 = ~(input_a[31] | input_a[21]);
  assign popcount33_bqn3_core_145_not = ~input_a[5];
  assign popcount33_bqn3_core_146 = ~(input_a[21] | input_a[12]);
  assign popcount33_bqn3_core_147_not = ~input_a[25];
  assign popcount33_bqn3_core_150 = input_a[11] | input_a[26];
  assign popcount33_bqn3_core_151 = input_a[0] | input_a[13];
  assign popcount33_bqn3_core_154 = ~(input_a[19] & input_a[10]);
  assign popcount33_bqn3_core_157 = ~(input_a[4] | input_a[31]);
  assign popcount33_bqn3_core_160 = input_a[1] ^ input_a[10];
  assign popcount33_bqn3_core_161 = input_a[12] | input_a[29];
  assign popcount33_bqn3_core_163 = ~(input_a[19] & input_a[10]);
  assign popcount33_bqn3_core_165 = ~(input_a[5] | input_a[7]);
  assign popcount33_bqn3_core_166 = ~input_a[29];
  assign popcount33_bqn3_core_169 = ~(input_a[20] ^ input_a[29]);
  assign popcount33_bqn3_core_170 = ~input_a[17];
  assign popcount33_bqn3_core_171 = ~(input_a[1] ^ input_a[8]);
  assign popcount33_bqn3_core_172 = ~(input_a[18] & input_a[22]);
  assign popcount33_bqn3_core_173 = input_a[26] | input_a[18];
  assign popcount33_bqn3_core_174 = ~input_a[24];
  assign popcount33_bqn3_core_179 = ~input_a[23];
  assign popcount33_bqn3_core_180 = input_a[4] ^ input_a[28];
  assign popcount33_bqn3_core_181 = ~(input_a[3] & input_a[13]);
  assign popcount33_bqn3_core_184 = ~(input_a[5] ^ input_a[18]);
  assign popcount33_bqn3_core_186 = input_a[19] & input_a[11];
  assign popcount33_bqn3_core_188 = ~(input_a[7] | input_a[6]);
  assign popcount33_bqn3_core_191 = input_a[27] & input_a[13];
  assign popcount33_bqn3_core_192 = ~(input_a[0] ^ input_a[7]);
  assign popcount33_bqn3_core_193 = ~(input_a[24] & input_a[29]);
  assign popcount33_bqn3_core_194 = ~(input_a[27] & input_a[30]);
  assign popcount33_bqn3_core_198 = input_a[5] | input_a[0];
  assign popcount33_bqn3_core_199_not = ~input_a[31];
  assign popcount33_bqn3_core_200 = ~(input_a[8] | input_a[10]);
  assign popcount33_bqn3_core_201 = input_a[8] ^ input_a[32];
  assign popcount33_bqn3_core_203 = ~(input_a[9] | input_a[16]);
  assign popcount33_bqn3_core_204 = input_a[13] | input_a[29];
  assign popcount33_bqn3_core_205_not = ~input_a[11];
  assign popcount33_bqn3_core_206 = ~(input_a[3] ^ input_a[16]);
  assign popcount33_bqn3_core_207 = input_a[28] & input_a[17];
  assign popcount33_bqn3_core_208 = input_a[0] ^ input_a[0];
  assign popcount33_bqn3_core_209 = input_a[21] & input_a[5];
  assign popcount33_bqn3_core_211 = ~(input_a[4] & input_a[2]);
  assign popcount33_bqn3_core_212 = ~(input_a[8] ^ input_a[0]);
  assign popcount33_bqn3_core_213_not = ~input_a[0];
  assign popcount33_bqn3_core_215 = ~input_a[15];
  assign popcount33_bqn3_core_216 = ~input_a[11];
  assign popcount33_bqn3_core_219 = input_a[0] | input_a[12];
  assign popcount33_bqn3_core_220 = input_a[7] & input_a[20];
  assign popcount33_bqn3_core_223 = ~(input_a[5] | input_a[4]);
  assign popcount33_bqn3_core_224 = input_a[21] | input_a[31];
  assign popcount33_bqn3_core_225 = ~(input_a[20] & input_a[1]);
  assign popcount33_bqn3_core_226 = ~(input_a[19] | input_a[32]);
  assign popcount33_bqn3_core_227 = ~input_a[13];
  assign popcount33_bqn3_core_228 = ~input_a[26];
  assign popcount33_bqn3_core_230 = ~(input_a[18] | input_a[17]);
  assign popcount33_bqn3_core_232 = ~(input_a[26] & input_a[2]);
  assign popcount33_bqn3_core_233 = input_a[24] | input_a[26];
  assign popcount33_bqn3_core_234 = input_a[7] | input_a[6];
  assign popcount33_bqn3_core_235 = input_a[30] & input_a[20];
  assign popcount33_bqn3_core_236 = ~input_a[30];
  assign popcount33_bqn3_core_238 = input_a[25] & input_a[16];

  assign popcount33_bqn3_out[0] = 1'b1;
  assign popcount33_bqn3_out[1] = input_a[21];
  assign popcount33_bqn3_out[2] = input_a[24];
  assign popcount33_bqn3_out[3] = input_a[10];
  assign popcount33_bqn3_out[4] = input_a[25];
  assign popcount33_bqn3_out[5] = 1'b0;
endmodule