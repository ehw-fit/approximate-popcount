// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.76197
// WCE=10.0
// EP=0.823803%
// Printed PDK parameters:
//  Area=1104200.0
//  Delay=3380858.25
//  Power=35820.0

module popcount20_429r(input [19:0] input_a, output [4:0] popcount20_429r_out);
  wire popcount20_429r_core_022;
  wire popcount20_429r_core_025_not;
  wire popcount20_429r_core_026;
  wire popcount20_429r_core_032;
  wire popcount20_429r_core_033;
  wire popcount20_429r_core_034;
  wire popcount20_429r_core_035;
  wire popcount20_429r_core_036;
  wire popcount20_429r_core_037;
  wire popcount20_429r_core_038;
  wire popcount20_429r_core_040;
  wire popcount20_429r_core_041;
  wire popcount20_429r_core_042;
  wire popcount20_429r_core_043;
  wire popcount20_429r_core_045;
  wire popcount20_429r_core_046;
  wire popcount20_429r_core_047;
  wire popcount20_429r_core_049;
  wire popcount20_429r_core_050;
  wire popcount20_429r_core_051;
  wire popcount20_429r_core_052_not;
  wire popcount20_429r_core_053;
  wire popcount20_429r_core_056;
  wire popcount20_429r_core_059;
  wire popcount20_429r_core_060;
  wire popcount20_429r_core_061;
  wire popcount20_429r_core_062;
  wire popcount20_429r_core_063;
  wire popcount20_429r_core_065;
  wire popcount20_429r_core_066;
  wire popcount20_429r_core_069;
  wire popcount20_429r_core_070;
  wire popcount20_429r_core_071;
  wire popcount20_429r_core_072;
  wire popcount20_429r_core_073;
  wire popcount20_429r_core_074;
  wire popcount20_429r_core_076;
  wire popcount20_429r_core_077;
  wire popcount20_429r_core_078;
  wire popcount20_429r_core_079;
  wire popcount20_429r_core_082;
  wire popcount20_429r_core_084;
  wire popcount20_429r_core_085;
  wire popcount20_429r_core_086;
  wire popcount20_429r_core_087;
  wire popcount20_429r_core_088;
  wire popcount20_429r_core_089;
  wire popcount20_429r_core_090;
  wire popcount20_429r_core_091;
  wire popcount20_429r_core_096;
  wire popcount20_429r_core_097_not;
  wire popcount20_429r_core_098;
  wire popcount20_429r_core_099_not;
  wire popcount20_429r_core_100;
  wire popcount20_429r_core_102;
  wire popcount20_429r_core_106;
  wire popcount20_429r_core_107;
  wire popcount20_429r_core_109;
  wire popcount20_429r_core_110;
  wire popcount20_429r_core_111;
  wire popcount20_429r_core_112;
  wire popcount20_429r_core_113;
  wire popcount20_429r_core_116_not;
  wire popcount20_429r_core_117;
  wire popcount20_429r_core_120;
  wire popcount20_429r_core_121;
  wire popcount20_429r_core_122;
  wire popcount20_429r_core_123;
  wire popcount20_429r_core_125;
  wire popcount20_429r_core_126;
  wire popcount20_429r_core_127;
  wire popcount20_429r_core_128;
  wire popcount20_429r_core_130;
  wire popcount20_429r_core_131;
  wire popcount20_429r_core_132;
  wire popcount20_429r_core_133;
  wire popcount20_429r_core_135;
  wire popcount20_429r_core_136;
  wire popcount20_429r_core_138;
  wire popcount20_429r_core_140;
  wire popcount20_429r_core_143;
  wire popcount20_429r_core_144;
  wire popcount20_429r_core_145;

  assign popcount20_429r_core_022 = input_a[0] ^ input_a[8];
  assign popcount20_429r_core_025_not = ~input_a[15];
  assign popcount20_429r_core_026 = ~(input_a[14] & input_a[14]);
  assign popcount20_429r_core_032 = ~input_a[1];
  assign popcount20_429r_core_033 = input_a[7] | input_a[9];
  assign popcount20_429r_core_034 = ~(input_a[9] & input_a[16]);
  assign popcount20_429r_core_035 = ~(input_a[8] ^ input_a[13]);
  assign popcount20_429r_core_036 = ~input_a[17];
  assign popcount20_429r_core_037 = ~(input_a[3] ^ input_a[15]);
  assign popcount20_429r_core_038 = input_a[14] | input_a[1];
  assign popcount20_429r_core_040 = ~(input_a[13] ^ input_a[19]);
  assign popcount20_429r_core_041 = ~(input_a[5] & input_a[3]);
  assign popcount20_429r_core_042 = ~(input_a[15] | input_a[3]);
  assign popcount20_429r_core_043 = input_a[0] ^ input_a[17];
  assign popcount20_429r_core_045 = input_a[12] & input_a[3];
  assign popcount20_429r_core_046 = ~(input_a[5] & input_a[4]);
  assign popcount20_429r_core_047 = input_a[12] & input_a[10];
  assign popcount20_429r_core_049 = input_a[14] | input_a[4];
  assign popcount20_429r_core_050 = input_a[11] ^ input_a[1];
  assign popcount20_429r_core_051 = ~(input_a[18] | input_a[8]);
  assign popcount20_429r_core_052_not = ~input_a[9];
  assign popcount20_429r_core_053 = input_a[5] ^ input_a[18];
  assign popcount20_429r_core_056 = ~(input_a[7] & input_a[14]);
  assign popcount20_429r_core_059 = input_a[15] ^ input_a[0];
  assign popcount20_429r_core_060 = input_a[16] ^ input_a[0];
  assign popcount20_429r_core_061 = ~(input_a[7] & input_a[3]);
  assign popcount20_429r_core_062 = input_a[0] & input_a[13];
  assign popcount20_429r_core_063 = ~input_a[8];
  assign popcount20_429r_core_065 = ~(input_a[10] ^ input_a[16]);
  assign popcount20_429r_core_066 = ~(input_a[3] | input_a[1]);
  assign popcount20_429r_core_069 = input_a[7] ^ input_a[3];
  assign popcount20_429r_core_070 = ~(input_a[12] & input_a[17]);
  assign popcount20_429r_core_071 = input_a[3] | input_a[9];
  assign popcount20_429r_core_072 = input_a[10] | input_a[8];
  assign popcount20_429r_core_073 = ~(input_a[8] & input_a[12]);
  assign popcount20_429r_core_074 = ~(input_a[5] & input_a[9]);
  assign popcount20_429r_core_076 = ~(input_a[2] & input_a[1]);
  assign popcount20_429r_core_077 = input_a[10] & input_a[17];
  assign popcount20_429r_core_078 = ~input_a[3];
  assign popcount20_429r_core_079 = ~input_a[10];
  assign popcount20_429r_core_082 = ~(input_a[0] & input_a[9]);
  assign popcount20_429r_core_084 = input_a[7] ^ input_a[16];
  assign popcount20_429r_core_085 = ~(input_a[0] & input_a[0]);
  assign popcount20_429r_core_086 = ~(input_a[12] | input_a[3]);
  assign popcount20_429r_core_087 = input_a[15] ^ input_a[12];
  assign popcount20_429r_core_088 = input_a[18] | input_a[2];
  assign popcount20_429r_core_089 = ~input_a[9];
  assign popcount20_429r_core_090 = ~input_a[15];
  assign popcount20_429r_core_091 = ~(input_a[2] | input_a[19]);
  assign popcount20_429r_core_096 = input_a[9] ^ input_a[2];
  assign popcount20_429r_core_097_not = ~input_a[9];
  assign popcount20_429r_core_098 = input_a[8] ^ input_a[7];
  assign popcount20_429r_core_099_not = ~input_a[12];
  assign popcount20_429r_core_100 = ~(input_a[2] & input_a[4]);
  assign popcount20_429r_core_102 = ~(input_a[18] | input_a[4]);
  assign popcount20_429r_core_106 = ~(input_a[3] | input_a[19]);
  assign popcount20_429r_core_107 = input_a[5] ^ input_a[12];
  assign popcount20_429r_core_109 = ~(input_a[2] | input_a[14]);
  assign popcount20_429r_core_110 = input_a[18] ^ input_a[17];
  assign popcount20_429r_core_111 = ~(input_a[19] | input_a[4]);
  assign popcount20_429r_core_112 = ~input_a[19];
  assign popcount20_429r_core_113 = input_a[4] | input_a[10];
  assign popcount20_429r_core_116_not = ~popcount20_429r_core_113;
  assign popcount20_429r_core_117 = ~(input_a[6] & input_a[11]);
  assign popcount20_429r_core_120 = ~(input_a[16] | input_a[19]);
  assign popcount20_429r_core_121 = ~(input_a[17] & input_a[2]);
  assign popcount20_429r_core_122 = ~(input_a[0] | input_a[8]);
  assign popcount20_429r_core_123 = input_a[11] | input_a[6];
  assign popcount20_429r_core_125 = ~(input_a[1] ^ input_a[7]);
  assign popcount20_429r_core_126 = ~input_a[11];
  assign popcount20_429r_core_127 = ~(input_a[18] ^ input_a[12]);
  assign popcount20_429r_core_128 = ~(input_a[12] | input_a[4]);
  assign popcount20_429r_core_130 = ~(input_a[2] | input_a[3]);
  assign popcount20_429r_core_131 = input_a[19] | popcount20_429r_core_116_not;
  assign popcount20_429r_core_132 = ~(input_a[5] | input_a[18]);
  assign popcount20_429r_core_133 = popcount20_429r_core_131 ^ input_a[19];
  assign popcount20_429r_core_135 = input_a[4] | input_a[19];
  assign popcount20_429r_core_136 = input_a[7] | input_a[11];
  assign popcount20_429r_core_138 = input_a[10] | popcount20_429r_core_135;
  assign popcount20_429r_core_140 = ~(input_a[4] & input_a[0]);
  assign popcount20_429r_core_143 = input_a[2] | input_a[16];
  assign popcount20_429r_core_144 = input_a[19] ^ input_a[6];
  assign popcount20_429r_core_145 = ~(input_a[9] ^ input_a[1]);

  assign popcount20_429r_out[0] = input_a[16];
  assign popcount20_429r_out[1] = 1'b1;
  assign popcount20_429r_out[2] = popcount20_429r_core_133;
  assign popcount20_429r_out[3] = popcount20_429r_core_138;
  assign popcount20_429r_out[4] = 1'b0;
endmodule