// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.14024
// WCE=18.0
// EP=0.951113%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_2a7j(input [27:0] input_a, output [4:0] popcount28_2a7j_out);
  wire popcount28_2a7j_core_032;
  wire popcount28_2a7j_core_033;
  wire popcount28_2a7j_core_034;
  wire popcount28_2a7j_core_036;
  wire popcount28_2a7j_core_037;
  wire popcount28_2a7j_core_038;
  wire popcount28_2a7j_core_039;
  wire popcount28_2a7j_core_040;
  wire popcount28_2a7j_core_042;
  wire popcount28_2a7j_core_043;
  wire popcount28_2a7j_core_046;
  wire popcount28_2a7j_core_047;
  wire popcount28_2a7j_core_049;
  wire popcount28_2a7j_core_050;
  wire popcount28_2a7j_core_051;
  wire popcount28_2a7j_core_053;
  wire popcount28_2a7j_core_054;
  wire popcount28_2a7j_core_055;
  wire popcount28_2a7j_core_056;
  wire popcount28_2a7j_core_058;
  wire popcount28_2a7j_core_060;
  wire popcount28_2a7j_core_062;
  wire popcount28_2a7j_core_063;
  wire popcount28_2a7j_core_064;
  wire popcount28_2a7j_core_065;
  wire popcount28_2a7j_core_066_not;
  wire popcount28_2a7j_core_067;
  wire popcount28_2a7j_core_068;
  wire popcount28_2a7j_core_070;
  wire popcount28_2a7j_core_071_not;
  wire popcount28_2a7j_core_072;
  wire popcount28_2a7j_core_073;
  wire popcount28_2a7j_core_074;
  wire popcount28_2a7j_core_075;
  wire popcount28_2a7j_core_077;
  wire popcount28_2a7j_core_080;
  wire popcount28_2a7j_core_081;
  wire popcount28_2a7j_core_083;
  wire popcount28_2a7j_core_086;
  wire popcount28_2a7j_core_087;
  wire popcount28_2a7j_core_088;
  wire popcount28_2a7j_core_089;
  wire popcount28_2a7j_core_092;
  wire popcount28_2a7j_core_094;
  wire popcount28_2a7j_core_095;
  wire popcount28_2a7j_core_097;
  wire popcount28_2a7j_core_099;
  wire popcount28_2a7j_core_101;
  wire popcount28_2a7j_core_102;
  wire popcount28_2a7j_core_105;
  wire popcount28_2a7j_core_106_not;
  wire popcount28_2a7j_core_108;
  wire popcount28_2a7j_core_109;
  wire popcount28_2a7j_core_110;
  wire popcount28_2a7j_core_112;
  wire popcount28_2a7j_core_113;
  wire popcount28_2a7j_core_115_not;
  wire popcount28_2a7j_core_118;
  wire popcount28_2a7j_core_119;
  wire popcount28_2a7j_core_120;
  wire popcount28_2a7j_core_121;
  wire popcount28_2a7j_core_122;
  wire popcount28_2a7j_core_123;
  wire popcount28_2a7j_core_124;
  wire popcount28_2a7j_core_126;
  wire popcount28_2a7j_core_127;
  wire popcount28_2a7j_core_130;
  wire popcount28_2a7j_core_132;
  wire popcount28_2a7j_core_133_not;
  wire popcount28_2a7j_core_135;
  wire popcount28_2a7j_core_136;
  wire popcount28_2a7j_core_137;
  wire popcount28_2a7j_core_138;
  wire popcount28_2a7j_core_139;
  wire popcount28_2a7j_core_141;
  wire popcount28_2a7j_core_142;
  wire popcount28_2a7j_core_143;
  wire popcount28_2a7j_core_144;
  wire popcount28_2a7j_core_146;
  wire popcount28_2a7j_core_147;
  wire popcount28_2a7j_core_148;
  wire popcount28_2a7j_core_150;
  wire popcount28_2a7j_core_151;
  wire popcount28_2a7j_core_152;
  wire popcount28_2a7j_core_153;
  wire popcount28_2a7j_core_154;
  wire popcount28_2a7j_core_155;
  wire popcount28_2a7j_core_156_not;
  wire popcount28_2a7j_core_157;
  wire popcount28_2a7j_core_161;
  wire popcount28_2a7j_core_162;
  wire popcount28_2a7j_core_163;
  wire popcount28_2a7j_core_164;
  wire popcount28_2a7j_core_165;
  wire popcount28_2a7j_core_166;
  wire popcount28_2a7j_core_167;
  wire popcount28_2a7j_core_168;
  wire popcount28_2a7j_core_169;
  wire popcount28_2a7j_core_170;
  wire popcount28_2a7j_core_172;
  wire popcount28_2a7j_core_173;
  wire popcount28_2a7j_core_174;
  wire popcount28_2a7j_core_175;
  wire popcount28_2a7j_core_176;
  wire popcount28_2a7j_core_177;
  wire popcount28_2a7j_core_178;
  wire popcount28_2a7j_core_179;
  wire popcount28_2a7j_core_182;
  wire popcount28_2a7j_core_184;
  wire popcount28_2a7j_core_185;
  wire popcount28_2a7j_core_186;
  wire popcount28_2a7j_core_187;
  wire popcount28_2a7j_core_188;
  wire popcount28_2a7j_core_189;
  wire popcount28_2a7j_core_191;
  wire popcount28_2a7j_core_195;
  wire popcount28_2a7j_core_196;
  wire popcount28_2a7j_core_198;
  wire popcount28_2a7j_core_200;
  wire popcount28_2a7j_core_201;

  assign popcount28_2a7j_core_032 = input_a[5] | input_a[1];
  assign popcount28_2a7j_core_033 = ~(input_a[24] & input_a[11]);
  assign popcount28_2a7j_core_034 = input_a[11] | input_a[26];
  assign popcount28_2a7j_core_036 = ~(input_a[21] & input_a[7]);
  assign popcount28_2a7j_core_037 = ~(input_a[24] | input_a[9]);
  assign popcount28_2a7j_core_038 = input_a[9] & input_a[15];
  assign popcount28_2a7j_core_039 = ~(input_a[7] ^ input_a[17]);
  assign popcount28_2a7j_core_040 = ~input_a[16];
  assign popcount28_2a7j_core_042 = ~(input_a[2] & input_a[9]);
  assign popcount28_2a7j_core_043 = input_a[7] ^ input_a[24];
  assign popcount28_2a7j_core_046 = ~input_a[23];
  assign popcount28_2a7j_core_047 = input_a[26] | input_a[22];
  assign popcount28_2a7j_core_049 = ~(input_a[17] & input_a[17]);
  assign popcount28_2a7j_core_050 = ~(input_a[3] & input_a[8]);
  assign popcount28_2a7j_core_051 = ~(input_a[19] | input_a[21]);
  assign popcount28_2a7j_core_053 = input_a[11] & input_a[8];
  assign popcount28_2a7j_core_054 = ~input_a[15];
  assign popcount28_2a7j_core_055 = input_a[21] | input_a[24];
  assign popcount28_2a7j_core_056 = ~(input_a[11] ^ input_a[19]);
  assign popcount28_2a7j_core_058 = ~(input_a[12] & input_a[24]);
  assign popcount28_2a7j_core_060 = input_a[7] | input_a[1];
  assign popcount28_2a7j_core_062 = ~(input_a[5] | input_a[2]);
  assign popcount28_2a7j_core_063 = input_a[23] & input_a[22];
  assign popcount28_2a7j_core_064 = ~(input_a[16] & input_a[9]);
  assign popcount28_2a7j_core_065 = input_a[16] ^ input_a[1];
  assign popcount28_2a7j_core_066_not = ~input_a[8];
  assign popcount28_2a7j_core_067 = input_a[1] & input_a[4];
  assign popcount28_2a7j_core_068 = ~input_a[19];
  assign popcount28_2a7j_core_070 = input_a[9] & input_a[3];
  assign popcount28_2a7j_core_071_not = ~input_a[23];
  assign popcount28_2a7j_core_072 = ~input_a[17];
  assign popcount28_2a7j_core_073 = ~(input_a[2] & input_a[3]);
  assign popcount28_2a7j_core_074 = ~(input_a[14] ^ input_a[11]);
  assign popcount28_2a7j_core_075 = ~(input_a[19] | input_a[25]);
  assign popcount28_2a7j_core_077 = ~(input_a[5] & input_a[21]);
  assign popcount28_2a7j_core_080 = ~(input_a[21] ^ input_a[27]);
  assign popcount28_2a7j_core_081 = input_a[20] ^ input_a[10];
  assign popcount28_2a7j_core_083 = ~input_a[12];
  assign popcount28_2a7j_core_086 = input_a[19] | input_a[17];
  assign popcount28_2a7j_core_087 = ~(input_a[2] & input_a[8]);
  assign popcount28_2a7j_core_088 = ~input_a[12];
  assign popcount28_2a7j_core_089 = input_a[27] & input_a[7];
  assign popcount28_2a7j_core_092 = input_a[22] | input_a[14];
  assign popcount28_2a7j_core_094 = ~(input_a[4] & input_a[24]);
  assign popcount28_2a7j_core_095 = ~(input_a[20] | input_a[21]);
  assign popcount28_2a7j_core_097 = input_a[0] | input_a[12];
  assign popcount28_2a7j_core_099 = ~input_a[17];
  assign popcount28_2a7j_core_101 = ~(input_a[14] & input_a[3]);
  assign popcount28_2a7j_core_102 = input_a[26] & input_a[26];
  assign popcount28_2a7j_core_105 = ~input_a[12];
  assign popcount28_2a7j_core_106_not = ~input_a[4];
  assign popcount28_2a7j_core_108 = input_a[10] | input_a[20];
  assign popcount28_2a7j_core_109 = ~(input_a[14] | input_a[20]);
  assign popcount28_2a7j_core_110 = ~(input_a[21] | input_a[5]);
  assign popcount28_2a7j_core_112 = input_a[26] & input_a[0];
  assign popcount28_2a7j_core_113 = input_a[23] ^ input_a[25];
  assign popcount28_2a7j_core_115_not = ~input_a[18];
  assign popcount28_2a7j_core_118 = input_a[9] ^ input_a[22];
  assign popcount28_2a7j_core_119 = ~(input_a[18] | input_a[13]);
  assign popcount28_2a7j_core_120 = input_a[27] & input_a[16];
  assign popcount28_2a7j_core_121 = ~input_a[19];
  assign popcount28_2a7j_core_122 = ~(input_a[18] | input_a[26]);
  assign popcount28_2a7j_core_123 = input_a[24] & input_a[15];
  assign popcount28_2a7j_core_124 = ~(input_a[13] & input_a[15]);
  assign popcount28_2a7j_core_126 = input_a[4] & input_a[15];
  assign popcount28_2a7j_core_127 = ~input_a[7];
  assign popcount28_2a7j_core_130 = input_a[8] ^ input_a[2];
  assign popcount28_2a7j_core_132 = ~(input_a[6] | input_a[26]);
  assign popcount28_2a7j_core_133_not = ~input_a[13];
  assign popcount28_2a7j_core_135 = ~input_a[26];
  assign popcount28_2a7j_core_136 = ~(input_a[1] | input_a[14]);
  assign popcount28_2a7j_core_137 = ~input_a[1];
  assign popcount28_2a7j_core_138 = input_a[18] ^ input_a[13];
  assign popcount28_2a7j_core_139 = input_a[12] ^ input_a[5];
  assign popcount28_2a7j_core_141 = ~input_a[16];
  assign popcount28_2a7j_core_142 = ~input_a[19];
  assign popcount28_2a7j_core_143 = ~input_a[27];
  assign popcount28_2a7j_core_144 = input_a[13] ^ input_a[21];
  assign popcount28_2a7j_core_146 = ~(input_a[16] | input_a[26]);
  assign popcount28_2a7j_core_147 = ~(input_a[5] | input_a[11]);
  assign popcount28_2a7j_core_148 = ~input_a[27];
  assign popcount28_2a7j_core_150 = input_a[3] & input_a[0];
  assign popcount28_2a7j_core_151 = ~(input_a[21] | input_a[2]);
  assign popcount28_2a7j_core_152 = input_a[23] & input_a[14];
  assign popcount28_2a7j_core_153 = ~(input_a[26] & input_a[10]);
  assign popcount28_2a7j_core_154 = input_a[14] | input_a[17];
  assign popcount28_2a7j_core_155 = ~(input_a[15] ^ input_a[21]);
  assign popcount28_2a7j_core_156_not = ~input_a[6];
  assign popcount28_2a7j_core_157 = ~input_a[21];
  assign popcount28_2a7j_core_161 = ~(input_a[24] | input_a[2]);
  assign popcount28_2a7j_core_162 = ~(input_a[11] | input_a[13]);
  assign popcount28_2a7j_core_163 = ~input_a[15];
  assign popcount28_2a7j_core_164 = input_a[22] ^ input_a[9];
  assign popcount28_2a7j_core_165 = ~(input_a[17] | input_a[15]);
  assign popcount28_2a7j_core_166 = ~(input_a[18] ^ input_a[7]);
  assign popcount28_2a7j_core_167 = ~(input_a[4] | input_a[2]);
  assign popcount28_2a7j_core_168 = ~input_a[14];
  assign popcount28_2a7j_core_169 = input_a[12] & input_a[14];
  assign popcount28_2a7j_core_170 = ~input_a[25];
  assign popcount28_2a7j_core_172 = input_a[9] & input_a[21];
  assign popcount28_2a7j_core_173 = ~(input_a[25] | input_a[9]);
  assign popcount28_2a7j_core_174 = input_a[1] & input_a[12];
  assign popcount28_2a7j_core_175 = input_a[6] | input_a[21];
  assign popcount28_2a7j_core_176 = ~(input_a[12] | input_a[19]);
  assign popcount28_2a7j_core_177 = ~(input_a[3] & input_a[7]);
  assign popcount28_2a7j_core_178 = input_a[21] & input_a[26];
  assign popcount28_2a7j_core_179 = ~input_a[22];
  assign popcount28_2a7j_core_182 = input_a[1] | input_a[0];
  assign popcount28_2a7j_core_184 = input_a[17] | input_a[25];
  assign popcount28_2a7j_core_185 = input_a[4] | input_a[17];
  assign popcount28_2a7j_core_186 = input_a[13] ^ input_a[0];
  assign popcount28_2a7j_core_187 = input_a[16] | input_a[16];
  assign popcount28_2a7j_core_188 = ~input_a[2];
  assign popcount28_2a7j_core_189 = input_a[16] | input_a[18];
  assign popcount28_2a7j_core_191 = ~(input_a[24] & input_a[26]);
  assign popcount28_2a7j_core_195 = input_a[21] & input_a[5];
  assign popcount28_2a7j_core_196 = ~(input_a[0] | input_a[19]);
  assign popcount28_2a7j_core_198 = ~(input_a[16] | input_a[15]);
  assign popcount28_2a7j_core_200 = ~input_a[11];
  assign popcount28_2a7j_core_201 = ~(input_a[12] ^ input_a[11]);

  assign popcount28_2a7j_out[0] = 1'b1;
  assign popcount28_2a7j_out[1] = input_a[24];
  assign popcount28_2a7j_out[2] = 1'b0;
  assign popcount28_2a7j_out[3] = 1'b0;
  assign popcount28_2a7j_out[4] = 1'b1;
endmodule