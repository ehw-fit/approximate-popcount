// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.42553
// WCE=18.0
// EP=0.915034%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_5gm3(input [22:0] input_a, output [4:0] popcount23_5gm3_out);
  wire popcount23_5gm3_core_026;
  wire popcount23_5gm3_core_029;
  wire popcount23_5gm3_core_030;
  wire popcount23_5gm3_core_031;
  wire popcount23_5gm3_core_036;
  wire popcount23_5gm3_core_037;
  wire popcount23_5gm3_core_039;
  wire popcount23_5gm3_core_042;
  wire popcount23_5gm3_core_043;
  wire popcount23_5gm3_core_045;
  wire popcount23_5gm3_core_046_not;
  wire popcount23_5gm3_core_048;
  wire popcount23_5gm3_core_049;
  wire popcount23_5gm3_core_050;
  wire popcount23_5gm3_core_052;
  wire popcount23_5gm3_core_055;
  wire popcount23_5gm3_core_058;
  wire popcount23_5gm3_core_059;
  wire popcount23_5gm3_core_062;
  wire popcount23_5gm3_core_065;
  wire popcount23_5gm3_core_066;
  wire popcount23_5gm3_core_067;
  wire popcount23_5gm3_core_069;
  wire popcount23_5gm3_core_071;
  wire popcount23_5gm3_core_072;
  wire popcount23_5gm3_core_073;
  wire popcount23_5gm3_core_074;
  wire popcount23_5gm3_core_076;
  wire popcount23_5gm3_core_077;
  wire popcount23_5gm3_core_080;
  wire popcount23_5gm3_core_081;
  wire popcount23_5gm3_core_082;
  wire popcount23_5gm3_core_086;
  wire popcount23_5gm3_core_090;
  wire popcount23_5gm3_core_093;
  wire popcount23_5gm3_core_096;
  wire popcount23_5gm3_core_097;
  wire popcount23_5gm3_core_098;
  wire popcount23_5gm3_core_099;
  wire popcount23_5gm3_core_102;
  wire popcount23_5gm3_core_103;
  wire popcount23_5gm3_core_106;
  wire popcount23_5gm3_core_107;
  wire popcount23_5gm3_core_108;
  wire popcount23_5gm3_core_109;
  wire popcount23_5gm3_core_110;
  wire popcount23_5gm3_core_112;
  wire popcount23_5gm3_core_113;
  wire popcount23_5gm3_core_114_not;
  wire popcount23_5gm3_core_116;
  wire popcount23_5gm3_core_117;
  wire popcount23_5gm3_core_118;
  wire popcount23_5gm3_core_119;
  wire popcount23_5gm3_core_121;
  wire popcount23_5gm3_core_122;
  wire popcount23_5gm3_core_125;
  wire popcount23_5gm3_core_126;
  wire popcount23_5gm3_core_127;
  wire popcount23_5gm3_core_128;
  wire popcount23_5gm3_core_130;
  wire popcount23_5gm3_core_131;
  wire popcount23_5gm3_core_133;
  wire popcount23_5gm3_core_134;
  wire popcount23_5gm3_core_135;
  wire popcount23_5gm3_core_136;
  wire popcount23_5gm3_core_139;
  wire popcount23_5gm3_core_143;
  wire popcount23_5gm3_core_145;
  wire popcount23_5gm3_core_147;
  wire popcount23_5gm3_core_148;
  wire popcount23_5gm3_core_149;
  wire popcount23_5gm3_core_152;
  wire popcount23_5gm3_core_153;
  wire popcount23_5gm3_core_155;
  wire popcount23_5gm3_core_157_not;
  wire popcount23_5gm3_core_159;
  wire popcount23_5gm3_core_160_not;
  wire popcount23_5gm3_core_161;
  wire popcount23_5gm3_core_162;
  wire popcount23_5gm3_core_163;
  wire popcount23_5gm3_core_166;
  wire popcount23_5gm3_core_169;

  assign popcount23_5gm3_core_026 = ~input_a[20];
  assign popcount23_5gm3_core_029 = input_a[9] ^ input_a[0];
  assign popcount23_5gm3_core_030 = input_a[2] ^ input_a[13];
  assign popcount23_5gm3_core_031 = ~(input_a[20] | input_a[12]);
  assign popcount23_5gm3_core_036 = input_a[12] ^ input_a[6];
  assign popcount23_5gm3_core_037 = ~(input_a[17] ^ input_a[5]);
  assign popcount23_5gm3_core_039 = input_a[7] ^ input_a[9];
  assign popcount23_5gm3_core_042 = ~(input_a[19] ^ input_a[10]);
  assign popcount23_5gm3_core_043 = input_a[6] ^ input_a[17];
  assign popcount23_5gm3_core_045 = ~(input_a[4] & input_a[9]);
  assign popcount23_5gm3_core_046_not = ~input_a[15];
  assign popcount23_5gm3_core_048 = ~(input_a[21] & input_a[21]);
  assign popcount23_5gm3_core_049 = ~(input_a[8] | input_a[1]);
  assign popcount23_5gm3_core_050 = ~(input_a[19] | input_a[6]);
  assign popcount23_5gm3_core_052 = input_a[7] ^ input_a[9];
  assign popcount23_5gm3_core_055 = input_a[9] | input_a[11];
  assign popcount23_5gm3_core_058 = input_a[21] ^ input_a[18];
  assign popcount23_5gm3_core_059 = ~(input_a[18] | input_a[17]);
  assign popcount23_5gm3_core_062 = ~(input_a[11] ^ input_a[10]);
  assign popcount23_5gm3_core_065 = ~input_a[8];
  assign popcount23_5gm3_core_066 = ~(input_a[10] ^ input_a[22]);
  assign popcount23_5gm3_core_067 = input_a[1] & input_a[5];
  assign popcount23_5gm3_core_069 = input_a[10] & input_a[16];
  assign popcount23_5gm3_core_071 = ~(input_a[13] | input_a[2]);
  assign popcount23_5gm3_core_072 = input_a[4] & input_a[7];
  assign popcount23_5gm3_core_073 = ~(input_a[18] & input_a[8]);
  assign popcount23_5gm3_core_074 = ~(input_a[22] | input_a[7]);
  assign popcount23_5gm3_core_076 = ~(input_a[16] & input_a[10]);
  assign popcount23_5gm3_core_077 = input_a[3] | input_a[18];
  assign popcount23_5gm3_core_080 = ~(input_a[3] & input_a[21]);
  assign popcount23_5gm3_core_081 = ~(input_a[19] | input_a[1]);
  assign popcount23_5gm3_core_082 = input_a[2] & input_a[16];
  assign popcount23_5gm3_core_086 = ~(input_a[21] | input_a[4]);
  assign popcount23_5gm3_core_090 = input_a[18] | input_a[11];
  assign popcount23_5gm3_core_093 = ~(input_a[16] ^ input_a[15]);
  assign popcount23_5gm3_core_096 = ~(input_a[15] & input_a[15]);
  assign popcount23_5gm3_core_097 = ~(input_a[9] | input_a[21]);
  assign popcount23_5gm3_core_098 = ~(input_a[18] & input_a[18]);
  assign popcount23_5gm3_core_099 = input_a[7] & input_a[18];
  assign popcount23_5gm3_core_102 = input_a[17] | input_a[7];
  assign popcount23_5gm3_core_103 = ~(input_a[1] ^ input_a[15]);
  assign popcount23_5gm3_core_106 = ~input_a[2];
  assign popcount23_5gm3_core_107 = input_a[1] | input_a[17];
  assign popcount23_5gm3_core_108 = input_a[13] | input_a[4];
  assign popcount23_5gm3_core_109 = ~input_a[3];
  assign popcount23_5gm3_core_110 = input_a[0] | input_a[1];
  assign popcount23_5gm3_core_112 = ~(input_a[4] & input_a[17]);
  assign popcount23_5gm3_core_113 = input_a[16] & input_a[3];
  assign popcount23_5gm3_core_114_not = ~input_a[12];
  assign popcount23_5gm3_core_116 = ~(input_a[6] & input_a[22]);
  assign popcount23_5gm3_core_117 = ~input_a[10];
  assign popcount23_5gm3_core_118 = input_a[8] | input_a[20];
  assign popcount23_5gm3_core_119 = input_a[12] & input_a[7];
  assign popcount23_5gm3_core_121 = ~input_a[7];
  assign popcount23_5gm3_core_122 = ~(input_a[10] & input_a[17]);
  assign popcount23_5gm3_core_125 = ~input_a[15];
  assign popcount23_5gm3_core_126 = input_a[10] | input_a[15];
  assign popcount23_5gm3_core_127 = input_a[12] ^ input_a[3];
  assign popcount23_5gm3_core_128 = input_a[1] ^ input_a[0];
  assign popcount23_5gm3_core_130 = ~input_a[14];
  assign popcount23_5gm3_core_131 = ~(input_a[9] | input_a[7]);
  assign popcount23_5gm3_core_133 = input_a[16] ^ input_a[0];
  assign popcount23_5gm3_core_134 = ~input_a[11];
  assign popcount23_5gm3_core_135 = ~(input_a[19] ^ input_a[3]);
  assign popcount23_5gm3_core_136 = input_a[2] | input_a[19];
  assign popcount23_5gm3_core_139 = ~input_a[9];
  assign popcount23_5gm3_core_143 = ~(input_a[13] & input_a[4]);
  assign popcount23_5gm3_core_145 = ~(input_a[11] ^ input_a[17]);
  assign popcount23_5gm3_core_147 = input_a[4] ^ input_a[11];
  assign popcount23_5gm3_core_148 = input_a[3] & input_a[19];
  assign popcount23_5gm3_core_149 = ~(input_a[10] | input_a[21]);
  assign popcount23_5gm3_core_152 = ~input_a[17];
  assign popcount23_5gm3_core_153 = input_a[4] & input_a[0];
  assign popcount23_5gm3_core_155 = input_a[12] | input_a[15];
  assign popcount23_5gm3_core_157_not = ~input_a[14];
  assign popcount23_5gm3_core_159 = input_a[2] | input_a[14];
  assign popcount23_5gm3_core_160_not = ~input_a[20];
  assign popcount23_5gm3_core_161 = input_a[14] | input_a[12];
  assign popcount23_5gm3_core_162 = ~(input_a[9] & input_a[5]);
  assign popcount23_5gm3_core_163 = ~(input_a[20] | input_a[7]);
  assign popcount23_5gm3_core_166 = input_a[14] | input_a[7];
  assign popcount23_5gm3_core_169 = ~(input_a[12] & input_a[18]);

  assign popcount23_5gm3_out[0] = 1'b0;
  assign popcount23_5gm3_out[1] = 1'b0;
  assign popcount23_5gm3_out[2] = 1'b1;
  assign popcount23_5gm3_out[3] = input_a[11];
  assign popcount23_5gm3_out[4] = 1'b0;
endmodule