// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.541
// WCE=47.0
// EP=0.990451%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount45_vpej(input [44:0] input_a, output [5:0] popcount45_vpej_out);
  wire popcount45_vpej_core_048;
  wire popcount45_vpej_core_049;
  wire popcount45_vpej_core_050_not;
  wire popcount45_vpej_core_052;
  wire popcount45_vpej_core_055;
  wire popcount45_vpej_core_056;
  wire popcount45_vpej_core_062;
  wire popcount45_vpej_core_063;
  wire popcount45_vpej_core_064;
  wire popcount45_vpej_core_065;
  wire popcount45_vpej_core_066;
  wire popcount45_vpej_core_070;
  wire popcount45_vpej_core_072;
  wire popcount45_vpej_core_073;
  wire popcount45_vpej_core_074;
  wire popcount45_vpej_core_075;
  wire popcount45_vpej_core_078;
  wire popcount45_vpej_core_080_not;
  wire popcount45_vpej_core_083;
  wire popcount45_vpej_core_084;
  wire popcount45_vpej_core_087;
  wire popcount45_vpej_core_091;
  wire popcount45_vpej_core_092;
  wire popcount45_vpej_core_093;
  wire popcount45_vpej_core_094;
  wire popcount45_vpej_core_095;
  wire popcount45_vpej_core_098;
  wire popcount45_vpej_core_099;
  wire popcount45_vpej_core_100;
  wire popcount45_vpej_core_101;
  wire popcount45_vpej_core_102;
  wire popcount45_vpej_core_103;
  wire popcount45_vpej_core_104;
  wire popcount45_vpej_core_105;
  wire popcount45_vpej_core_106;
  wire popcount45_vpej_core_107;
  wire popcount45_vpej_core_109;
  wire popcount45_vpej_core_110;
  wire popcount45_vpej_core_111;
  wire popcount45_vpej_core_112;
  wire popcount45_vpej_core_113;
  wire popcount45_vpej_core_114;
  wire popcount45_vpej_core_116;
  wire popcount45_vpej_core_119;
  wire popcount45_vpej_core_120;
  wire popcount45_vpej_core_122;
  wire popcount45_vpej_core_124;
  wire popcount45_vpej_core_126;
  wire popcount45_vpej_core_127;
  wire popcount45_vpej_core_129;
  wire popcount45_vpej_core_130;
  wire popcount45_vpej_core_131_not;
  wire popcount45_vpej_core_132;
  wire popcount45_vpej_core_133;
  wire popcount45_vpej_core_134;
  wire popcount45_vpej_core_137;
  wire popcount45_vpej_core_138;
  wire popcount45_vpej_core_140;
  wire popcount45_vpej_core_142;
  wire popcount45_vpej_core_143;
  wire popcount45_vpej_core_145;
  wire popcount45_vpej_core_146;
  wire popcount45_vpej_core_148;
  wire popcount45_vpej_core_150;
  wire popcount45_vpej_core_151;
  wire popcount45_vpej_core_152;
  wire popcount45_vpej_core_153;
  wire popcount45_vpej_core_155;
  wire popcount45_vpej_core_156;
  wire popcount45_vpej_core_157;
  wire popcount45_vpej_core_158;
  wire popcount45_vpej_core_159;
  wire popcount45_vpej_core_160;
  wire popcount45_vpej_core_161;
  wire popcount45_vpej_core_162;
  wire popcount45_vpej_core_163;
  wire popcount45_vpej_core_164_not;
  wire popcount45_vpej_core_167;
  wire popcount45_vpej_core_169;
  wire popcount45_vpej_core_173;
  wire popcount45_vpej_core_174;
  wire popcount45_vpej_core_175;
  wire popcount45_vpej_core_176;
  wire popcount45_vpej_core_177;
  wire popcount45_vpej_core_178;
  wire popcount45_vpej_core_181;
  wire popcount45_vpej_core_182;
  wire popcount45_vpej_core_183;
  wire popcount45_vpej_core_184;
  wire popcount45_vpej_core_186;
  wire popcount45_vpej_core_187;
  wire popcount45_vpej_core_189;
  wire popcount45_vpej_core_190;
  wire popcount45_vpej_core_191;
  wire popcount45_vpej_core_192;
  wire popcount45_vpej_core_193;
  wire popcount45_vpej_core_195;
  wire popcount45_vpej_core_197;
  wire popcount45_vpej_core_198;
  wire popcount45_vpej_core_203;
  wire popcount45_vpej_core_204_not;
  wire popcount45_vpej_core_206;
  wire popcount45_vpej_core_207;
  wire popcount45_vpej_core_209;
  wire popcount45_vpej_core_210;
  wire popcount45_vpej_core_211;
  wire popcount45_vpej_core_212;
  wire popcount45_vpej_core_213;
  wire popcount45_vpej_core_214;
  wire popcount45_vpej_core_215;
  wire popcount45_vpej_core_216;
  wire popcount45_vpej_core_217;
  wire popcount45_vpej_core_218;
  wire popcount45_vpej_core_221;
  wire popcount45_vpej_core_222;
  wire popcount45_vpej_core_223;
  wire popcount45_vpej_core_224;
  wire popcount45_vpej_core_226;
  wire popcount45_vpej_core_228;
  wire popcount45_vpej_core_232;
  wire popcount45_vpej_core_233;
  wire popcount45_vpej_core_234;
  wire popcount45_vpej_core_235;
  wire popcount45_vpej_core_236;
  wire popcount45_vpej_core_237;
  wire popcount45_vpej_core_239;
  wire popcount45_vpej_core_240;
  wire popcount45_vpej_core_242;
  wire popcount45_vpej_core_243;
  wire popcount45_vpej_core_246;
  wire popcount45_vpej_core_250;
  wire popcount45_vpej_core_251;
  wire popcount45_vpej_core_253;
  wire popcount45_vpej_core_254;
  wire popcount45_vpej_core_255;
  wire popcount45_vpej_core_256;
  wire popcount45_vpej_core_258;
  wire popcount45_vpej_core_259;
  wire popcount45_vpej_core_260;
  wire popcount45_vpej_core_265;
  wire popcount45_vpej_core_266;
  wire popcount45_vpej_core_268;
  wire popcount45_vpej_core_272;
  wire popcount45_vpej_core_274;
  wire popcount45_vpej_core_276;
  wire popcount45_vpej_core_277;
  wire popcount45_vpej_core_278;
  wire popcount45_vpej_core_282;
  wire popcount45_vpej_core_283;
  wire popcount45_vpej_core_285;
  wire popcount45_vpej_core_286;
  wire popcount45_vpej_core_287;
  wire popcount45_vpej_core_288;
  wire popcount45_vpej_core_290;
  wire popcount45_vpej_core_291;
  wire popcount45_vpej_core_292;
  wire popcount45_vpej_core_293;
  wire popcount45_vpej_core_294;
  wire popcount45_vpej_core_295;
  wire popcount45_vpej_core_296;
  wire popcount45_vpej_core_298;
  wire popcount45_vpej_core_299;
  wire popcount45_vpej_core_300;
  wire popcount45_vpej_core_302;
  wire popcount45_vpej_core_304;
  wire popcount45_vpej_core_305;
  wire popcount45_vpej_core_308;
  wire popcount45_vpej_core_314;
  wire popcount45_vpej_core_315;
  wire popcount45_vpej_core_317;
  wire popcount45_vpej_core_318;
  wire popcount45_vpej_core_320;
  wire popcount45_vpej_core_321;
  wire popcount45_vpej_core_323;
  wire popcount45_vpej_core_324;
  wire popcount45_vpej_core_325;
  wire popcount45_vpej_core_326;
  wire popcount45_vpej_core_327;
  wire popcount45_vpej_core_330;
  wire popcount45_vpej_core_332;
  wire popcount45_vpej_core_334;
  wire popcount45_vpej_core_336;
  wire popcount45_vpej_core_338;
  wire popcount45_vpej_core_340;
  wire popcount45_vpej_core_341;
  wire popcount45_vpej_core_343;
  wire popcount45_vpej_core_345;
  wire popcount45_vpej_core_346;
  wire popcount45_vpej_core_348;
  wire popcount45_vpej_core_349;
  wire popcount45_vpej_core_352;
  wire popcount45_vpej_core_353;
  wire popcount45_vpej_core_355;
  wire popcount45_vpej_core_356;

  assign popcount45_vpej_core_048 = input_a[34] | input_a[1];
  assign popcount45_vpej_core_049 = ~input_a[22];
  assign popcount45_vpej_core_050_not = ~input_a[31];
  assign popcount45_vpej_core_052 = ~(input_a[31] & input_a[5]);
  assign popcount45_vpej_core_055 = ~(input_a[13] ^ input_a[26]);
  assign popcount45_vpej_core_056 = input_a[30] & input_a[38];
  assign popcount45_vpej_core_062 = ~(input_a[6] & input_a[27]);
  assign popcount45_vpej_core_063 = input_a[28] | input_a[38];
  assign popcount45_vpej_core_064 = input_a[21] | input_a[34];
  assign popcount45_vpej_core_065 = ~(input_a[41] & input_a[3]);
  assign popcount45_vpej_core_066 = input_a[38] | input_a[31];
  assign popcount45_vpej_core_070 = ~(input_a[35] ^ input_a[37]);
  assign popcount45_vpej_core_072 = ~(input_a[26] & input_a[10]);
  assign popcount45_vpej_core_073 = ~(input_a[35] & input_a[9]);
  assign popcount45_vpej_core_074 = ~input_a[16];
  assign popcount45_vpej_core_075 = ~input_a[0];
  assign popcount45_vpej_core_078 = input_a[7] ^ input_a[12];
  assign popcount45_vpej_core_080_not = ~input_a[36];
  assign popcount45_vpej_core_083 = ~(input_a[28] & input_a[7]);
  assign popcount45_vpej_core_084 = ~input_a[25];
  assign popcount45_vpej_core_087 = ~(input_a[33] & input_a[32]);
  assign popcount45_vpej_core_091 = input_a[29] | input_a[30];
  assign popcount45_vpej_core_092 = ~(input_a[44] ^ input_a[37]);
  assign popcount45_vpej_core_093 = input_a[30] & input_a[29];
  assign popcount45_vpej_core_094 = ~(input_a[11] | input_a[43]);
  assign popcount45_vpej_core_095 = ~(input_a[8] ^ input_a[37]);
  assign popcount45_vpej_core_098 = ~(input_a[35] ^ input_a[38]);
  assign popcount45_vpej_core_099 = input_a[42] | input_a[26];
  assign popcount45_vpej_core_100 = ~input_a[43];
  assign popcount45_vpej_core_101 = input_a[27] | input_a[27];
  assign popcount45_vpej_core_102 = ~(input_a[13] ^ input_a[40]);
  assign popcount45_vpej_core_103 = input_a[20] ^ input_a[44];
  assign popcount45_vpej_core_104 = input_a[29] & input_a[39];
  assign popcount45_vpej_core_105 = ~(input_a[23] | input_a[8]);
  assign popcount45_vpej_core_106 = input_a[7] ^ input_a[13];
  assign popcount45_vpej_core_107 = ~(input_a[3] | input_a[27]);
  assign popcount45_vpej_core_109 = input_a[15] & input_a[5];
  assign popcount45_vpej_core_110 = ~(input_a[44] ^ input_a[24]);
  assign popcount45_vpej_core_111 = input_a[36] | input_a[32];
  assign popcount45_vpej_core_112 = input_a[33] | input_a[13];
  assign popcount45_vpej_core_113 = ~(input_a[34] | input_a[5]);
  assign popcount45_vpej_core_114 = input_a[39] & input_a[40];
  assign popcount45_vpej_core_116 = ~(input_a[29] ^ input_a[29]);
  assign popcount45_vpej_core_119 = ~(input_a[32] | input_a[10]);
  assign popcount45_vpej_core_120 = ~(input_a[35] ^ input_a[13]);
  assign popcount45_vpej_core_122 = input_a[20] & input_a[41];
  assign popcount45_vpej_core_124 = ~(input_a[3] ^ input_a[11]);
  assign popcount45_vpej_core_126 = input_a[13] ^ input_a[23];
  assign popcount45_vpej_core_127 = ~(input_a[37] ^ input_a[32]);
  assign popcount45_vpej_core_129 = ~(input_a[10] | input_a[2]);
  assign popcount45_vpej_core_130 = ~input_a[22];
  assign popcount45_vpej_core_131_not = ~input_a[21];
  assign popcount45_vpej_core_132 = ~(input_a[18] | input_a[35]);
  assign popcount45_vpej_core_133 = input_a[43] ^ input_a[43];
  assign popcount45_vpej_core_134 = ~input_a[12];
  assign popcount45_vpej_core_137 = ~(input_a[40] | input_a[37]);
  assign popcount45_vpej_core_138 = input_a[11] | input_a[43];
  assign popcount45_vpej_core_140 = input_a[8] ^ input_a[33];
  assign popcount45_vpej_core_142 = input_a[18] & input_a[8];
  assign popcount45_vpej_core_143 = ~(input_a[20] | input_a[5]);
  assign popcount45_vpej_core_145 = ~(input_a[24] & input_a[26]);
  assign popcount45_vpej_core_146 = ~(input_a[20] & input_a[23]);
  assign popcount45_vpej_core_148 = input_a[44] & input_a[43];
  assign popcount45_vpej_core_150 = input_a[34] | input_a[21];
  assign popcount45_vpej_core_151 = input_a[13] & input_a[2];
  assign popcount45_vpej_core_152 = input_a[8] & input_a[7];
  assign popcount45_vpej_core_153 = ~(input_a[23] ^ input_a[9]);
  assign popcount45_vpej_core_155 = ~input_a[42];
  assign popcount45_vpej_core_156 = ~(input_a[1] | input_a[10]);
  assign popcount45_vpej_core_157 = ~input_a[8];
  assign popcount45_vpej_core_158 = input_a[21] & input_a[15];
  assign popcount45_vpej_core_159 = input_a[24] | input_a[35];
  assign popcount45_vpej_core_160 = input_a[19] & input_a[29];
  assign popcount45_vpej_core_161 = input_a[32] & input_a[26];
  assign popcount45_vpej_core_162 = ~(input_a[30] ^ input_a[26]);
  assign popcount45_vpej_core_163 = ~input_a[21];
  assign popcount45_vpej_core_164_not = ~input_a[33];
  assign popcount45_vpej_core_167 = input_a[28] & input_a[18];
  assign popcount45_vpej_core_169 = ~(input_a[10] & input_a[34]);
  assign popcount45_vpej_core_173 = ~(input_a[6] & input_a[39]);
  assign popcount45_vpej_core_174 = ~(input_a[21] & input_a[0]);
  assign popcount45_vpej_core_175 = input_a[17] | input_a[9];
  assign popcount45_vpej_core_176 = input_a[34] & input_a[9];
  assign popcount45_vpej_core_177 = ~(input_a[12] | input_a[34]);
  assign popcount45_vpej_core_178 = ~(input_a[22] | input_a[43]);
  assign popcount45_vpej_core_181 = ~(input_a[37] | input_a[35]);
  assign popcount45_vpej_core_182 = ~(input_a[33] ^ input_a[14]);
  assign popcount45_vpej_core_183 = ~(input_a[29] ^ input_a[21]);
  assign popcount45_vpej_core_184 = input_a[42] ^ input_a[13];
  assign popcount45_vpej_core_186 = ~(input_a[5] | input_a[37]);
  assign popcount45_vpej_core_187 = ~(input_a[22] | input_a[6]);
  assign popcount45_vpej_core_189 = ~input_a[25];
  assign popcount45_vpej_core_190 = ~input_a[43];
  assign popcount45_vpej_core_191 = ~(input_a[16] | input_a[20]);
  assign popcount45_vpej_core_192 = input_a[36] & input_a[23];
  assign popcount45_vpej_core_193 = ~input_a[19];
  assign popcount45_vpej_core_195 = input_a[18] | input_a[9];
  assign popcount45_vpej_core_197 = ~(input_a[11] | input_a[42]);
  assign popcount45_vpej_core_198 = ~(input_a[1] | input_a[9]);
  assign popcount45_vpej_core_203 = ~(input_a[14] ^ input_a[22]);
  assign popcount45_vpej_core_204_not = ~input_a[31];
  assign popcount45_vpej_core_206 = input_a[4] ^ input_a[33];
  assign popcount45_vpej_core_207 = input_a[5] ^ input_a[42];
  assign popcount45_vpej_core_209 = input_a[22] ^ input_a[7];
  assign popcount45_vpej_core_210 = input_a[22] ^ input_a[15];
  assign popcount45_vpej_core_211 = input_a[31] & input_a[1];
  assign popcount45_vpej_core_212 = input_a[13] & input_a[24];
  assign popcount45_vpej_core_213 = input_a[14] | input_a[8];
  assign popcount45_vpej_core_214 = ~input_a[10];
  assign popcount45_vpej_core_215 = input_a[12] & input_a[14];
  assign popcount45_vpej_core_216 = ~(input_a[22] & input_a[19]);
  assign popcount45_vpej_core_217 = ~(input_a[26] & input_a[10]);
  assign popcount45_vpej_core_218 = input_a[25] ^ input_a[23];
  assign popcount45_vpej_core_221 = input_a[27] & input_a[24];
  assign popcount45_vpej_core_222 = input_a[7] & input_a[6];
  assign popcount45_vpej_core_223 = ~input_a[9];
  assign popcount45_vpej_core_224 = input_a[42] ^ input_a[44];
  assign popcount45_vpej_core_226 = input_a[16] & input_a[1];
  assign popcount45_vpej_core_228 = input_a[1] | input_a[23];
  assign popcount45_vpej_core_232 = input_a[25] ^ input_a[39];
  assign popcount45_vpej_core_233 = ~(input_a[31] | input_a[42]);
  assign popcount45_vpej_core_234 = ~(input_a[19] | input_a[24]);
  assign popcount45_vpej_core_235 = ~(input_a[13] ^ input_a[7]);
  assign popcount45_vpej_core_236 = ~(input_a[11] | input_a[0]);
  assign popcount45_vpej_core_237 = input_a[19] | input_a[16];
  assign popcount45_vpej_core_239 = ~(input_a[33] | input_a[28]);
  assign popcount45_vpej_core_240 = ~(input_a[3] ^ input_a[7]);
  assign popcount45_vpej_core_242 = ~(input_a[39] ^ input_a[14]);
  assign popcount45_vpej_core_243 = input_a[41] ^ input_a[28];
  assign popcount45_vpej_core_246 = ~(input_a[23] ^ input_a[7]);
  assign popcount45_vpej_core_250 = input_a[14] & input_a[41];
  assign popcount45_vpej_core_251 = ~input_a[29];
  assign popcount45_vpej_core_253 = input_a[32] & input_a[22];
  assign popcount45_vpej_core_254 = ~(input_a[22] & input_a[20]);
  assign popcount45_vpej_core_255 = ~(input_a[1] & input_a[15]);
  assign popcount45_vpej_core_256 = input_a[39] & input_a[12];
  assign popcount45_vpej_core_258 = input_a[5] | input_a[22];
  assign popcount45_vpej_core_259 = ~input_a[44];
  assign popcount45_vpej_core_260 = ~(input_a[25] & input_a[31]);
  assign popcount45_vpej_core_265 = ~input_a[15];
  assign popcount45_vpej_core_266 = ~(input_a[28] | input_a[41]);
  assign popcount45_vpej_core_268 = ~(input_a[11] | input_a[29]);
  assign popcount45_vpej_core_272 = input_a[28] & input_a[26];
  assign popcount45_vpej_core_274 = ~(input_a[33] | input_a[21]);
  assign popcount45_vpej_core_276 = ~input_a[16];
  assign popcount45_vpej_core_277 = ~(input_a[33] ^ input_a[27]);
  assign popcount45_vpej_core_278 = input_a[5] | input_a[4];
  assign popcount45_vpej_core_282 = input_a[37] ^ input_a[38];
  assign popcount45_vpej_core_283 = input_a[13] & input_a[37];
  assign popcount45_vpej_core_285 = ~(input_a[8] | input_a[24]);
  assign popcount45_vpej_core_286 = ~input_a[6];
  assign popcount45_vpej_core_287 = input_a[20] & input_a[24];
  assign popcount45_vpej_core_288 = input_a[29] ^ input_a[38];
  assign popcount45_vpej_core_290 = input_a[22] | input_a[23];
  assign popcount45_vpej_core_291 = ~(input_a[16] ^ input_a[34]);
  assign popcount45_vpej_core_292 = ~(input_a[2] | input_a[2]);
  assign popcount45_vpej_core_293 = ~(input_a[26] ^ input_a[1]);
  assign popcount45_vpej_core_294 = ~(input_a[43] & input_a[43]);
  assign popcount45_vpej_core_295 = input_a[41] ^ input_a[44];
  assign popcount45_vpej_core_296 = input_a[26] ^ input_a[14];
  assign popcount45_vpej_core_298 = ~input_a[42];
  assign popcount45_vpej_core_299 = ~(input_a[18] & input_a[20]);
  assign popcount45_vpej_core_300 = input_a[17] | input_a[21];
  assign popcount45_vpej_core_302 = ~input_a[14];
  assign popcount45_vpej_core_304 = ~input_a[25];
  assign popcount45_vpej_core_305 = ~(input_a[5] | input_a[30]);
  assign popcount45_vpej_core_308 = input_a[4] | input_a[29];
  assign popcount45_vpej_core_314 = ~input_a[20];
  assign popcount45_vpej_core_315 = input_a[21] & input_a[33];
  assign popcount45_vpej_core_317 = input_a[21] & input_a[25];
  assign popcount45_vpej_core_318 = ~input_a[6];
  assign popcount45_vpej_core_320 = ~(input_a[27] ^ input_a[3]);
  assign popcount45_vpej_core_321 = input_a[37] | input_a[30];
  assign popcount45_vpej_core_323 = input_a[41] ^ input_a[17];
  assign popcount45_vpej_core_324 = input_a[40] & input_a[22];
  assign popcount45_vpej_core_325 = ~(input_a[39] ^ input_a[10]);
  assign popcount45_vpej_core_326 = ~input_a[36];
  assign popcount45_vpej_core_327 = input_a[24] & input_a[9];
  assign popcount45_vpej_core_330 = input_a[0] & input_a[8];
  assign popcount45_vpej_core_332 = ~(input_a[21] | input_a[26]);
  assign popcount45_vpej_core_334 = ~(input_a[16] | input_a[37]);
  assign popcount45_vpej_core_336 = ~(input_a[40] & input_a[5]);
  assign popcount45_vpej_core_338 = ~(input_a[25] ^ input_a[41]);
  assign popcount45_vpej_core_340 = ~(input_a[22] & input_a[33]);
  assign popcount45_vpej_core_341 = input_a[0] ^ input_a[4];
  assign popcount45_vpej_core_343 = ~(input_a[7] ^ input_a[7]);
  assign popcount45_vpej_core_345 = input_a[22] & input_a[25];
  assign popcount45_vpej_core_346 = ~(input_a[2] ^ input_a[42]);
  assign popcount45_vpej_core_348 = input_a[26] | input_a[9];
  assign popcount45_vpej_core_349 = input_a[29] & input_a[18];
  assign popcount45_vpej_core_352 = ~input_a[16];
  assign popcount45_vpej_core_353 = input_a[32] ^ input_a[19];
  assign popcount45_vpej_core_355 = ~(input_a[2] | input_a[44]);
  assign popcount45_vpej_core_356 = input_a[24] & input_a[3];

  assign popcount45_vpej_out[0] = input_a[0];
  assign popcount45_vpej_out[1] = input_a[16];
  assign popcount45_vpej_out[2] = 1'b0;
  assign popcount45_vpej_out[3] = 1'b0;
  assign popcount45_vpej_out[4] = input_a[23];
  assign popcount45_vpej_out[5] = input_a[34];
endmodule