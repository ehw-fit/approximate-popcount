// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.56247
// WCE=57.0
// EP=0.95993%
// Printed PDK parameters:
//  Area=70292459.0
//  Delay=87106304.0
//  Power=2869900.0

module popcount45_pvta(input [44:0] input_a, output [5:0] popcount45_pvta_out);
  wire popcount45_pvta_core_047;
  wire popcount45_pvta_core_049;
  wire popcount45_pvta_core_051;
  wire popcount45_pvta_core_052;
  wire popcount45_pvta_core_055;
  wire popcount45_pvta_core_056;
  wire popcount45_pvta_core_057;
  wire popcount45_pvta_core_058;
  wire popcount45_pvta_core_059;
  wire popcount45_pvta_core_060;
  wire popcount45_pvta_core_061;
  wire popcount45_pvta_core_064;
  wire popcount45_pvta_core_065;
  wire popcount45_pvta_core_067;
  wire popcount45_pvta_core_068;
  wire popcount45_pvta_core_069;
  wire popcount45_pvta_core_070;
  wire popcount45_pvta_core_071;
  wire popcount45_pvta_core_072;
  wire popcount45_pvta_core_073;
  wire popcount45_pvta_core_074;
  wire popcount45_pvta_core_075;
  wire popcount45_pvta_core_078;
  wire popcount45_pvta_core_079;
  wire popcount45_pvta_core_083;
  wire popcount45_pvta_core_084;
  wire popcount45_pvta_core_085;
  wire popcount45_pvta_core_086;
  wire popcount45_pvta_core_087;
  wire popcount45_pvta_core_088;
  wire popcount45_pvta_core_089;
  wire popcount45_pvta_core_090;
  wire popcount45_pvta_core_091;
  wire popcount45_pvta_core_092;
  wire popcount45_pvta_core_093;
  wire popcount45_pvta_core_094;
  wire popcount45_pvta_core_095;
  wire popcount45_pvta_core_096;
  wire popcount45_pvta_core_097;
  wire popcount45_pvta_core_098;
  wire popcount45_pvta_core_099;
  wire popcount45_pvta_core_101;
  wire popcount45_pvta_core_102;
  wire popcount45_pvta_core_103;
  wire popcount45_pvta_core_104;
  wire popcount45_pvta_core_105;
  wire popcount45_pvta_core_106;
  wire popcount45_pvta_core_107;
  wire popcount45_pvta_core_108;
  wire popcount45_pvta_core_109;
  wire popcount45_pvta_core_110;
  wire popcount45_pvta_core_111;
  wire popcount45_pvta_core_112;
  wire popcount45_pvta_core_114;
  wire popcount45_pvta_core_115;
  wire popcount45_pvta_core_116;
  wire popcount45_pvta_core_117;
  wire popcount45_pvta_core_118;
  wire popcount45_pvta_core_122;
  wire popcount45_pvta_core_124;
  wire popcount45_pvta_core_125;
  wire popcount45_pvta_core_126;
  wire popcount45_pvta_core_127;
  wire popcount45_pvta_core_128;
  wire popcount45_pvta_core_129;
  wire popcount45_pvta_core_134_not;
  wire popcount45_pvta_core_136;
  wire popcount45_pvta_core_137;
  wire popcount45_pvta_core_138;
  wire popcount45_pvta_core_139;
  wire popcount45_pvta_core_140;
  wire popcount45_pvta_core_143;
  wire popcount45_pvta_core_144;
  wire popcount45_pvta_core_149;
  wire popcount45_pvta_core_152;
  wire popcount45_pvta_core_154;
  wire popcount45_pvta_core_155;
  wire popcount45_pvta_core_156;
  wire popcount45_pvta_core_157;
  wire popcount45_pvta_core_158;
  wire popcount45_pvta_core_159;
  wire popcount45_pvta_core_160;
  wire popcount45_pvta_core_161;
  wire popcount45_pvta_core_164;
  wire popcount45_pvta_core_165;
  wire popcount45_pvta_core_166;
  wire popcount45_pvta_core_167;
  wire popcount45_pvta_core_168;
  wire popcount45_pvta_core_169;
  wire popcount45_pvta_core_170;
  wire popcount45_pvta_core_171;
  wire popcount45_pvta_core_172;
  wire popcount45_pvta_core_173;
  wire popcount45_pvta_core_174;
  wire popcount45_pvta_core_175;
  wire popcount45_pvta_core_176;
  wire popcount45_pvta_core_177;
  wire popcount45_pvta_core_178;
  wire popcount45_pvta_core_179;
  wire popcount45_pvta_core_182;
  wire popcount45_pvta_core_183;
  wire popcount45_pvta_core_185;
  wire popcount45_pvta_core_186;
  wire popcount45_pvta_core_189;
  wire popcount45_pvta_core_193;
  wire popcount45_pvta_core_194;
  wire popcount45_pvta_core_195;
  wire popcount45_pvta_core_196;
  wire popcount45_pvta_core_197;
  wire popcount45_pvta_core_198;
  wire popcount45_pvta_core_199;
  wire popcount45_pvta_core_203;
  wire popcount45_pvta_core_204;
  wire popcount45_pvta_core_206;
  wire popcount45_pvta_core_207;
  wire popcount45_pvta_core_208;
  wire popcount45_pvta_core_209;
  wire popcount45_pvta_core_211;
  wire popcount45_pvta_core_212;
  wire popcount45_pvta_core_213;
  wire popcount45_pvta_core_214_not;
  wire popcount45_pvta_core_216;
  wire popcount45_pvta_core_217;
  wire popcount45_pvta_core_219;
  wire popcount45_pvta_core_220;
  wire popcount45_pvta_core_221;
  wire popcount45_pvta_core_222;
  wire popcount45_pvta_core_223;
  wire popcount45_pvta_core_224;
  wire popcount45_pvta_core_225;
  wire popcount45_pvta_core_226;
  wire popcount45_pvta_core_227;
  wire popcount45_pvta_core_228_not;
  wire popcount45_pvta_core_230;
  wire popcount45_pvta_core_231;
  wire popcount45_pvta_core_232;
  wire popcount45_pvta_core_233_not;
  wire popcount45_pvta_core_234;
  wire popcount45_pvta_core_235;
  wire popcount45_pvta_core_236;
  wire popcount45_pvta_core_237;
  wire popcount45_pvta_core_240;
  wire popcount45_pvta_core_241;
  wire popcount45_pvta_core_243;
  wire popcount45_pvta_core_245;
  wire popcount45_pvta_core_246;
  wire popcount45_pvta_core_249;
  wire popcount45_pvta_core_250;
  wire popcount45_pvta_core_251;
  wire popcount45_pvta_core_252;
  wire popcount45_pvta_core_253;
  wire popcount45_pvta_core_254;
  wire popcount45_pvta_core_255;
  wire popcount45_pvta_core_256;
  wire popcount45_pvta_core_259;
  wire popcount45_pvta_core_260;
  wire popcount45_pvta_core_264;
  wire popcount45_pvta_core_265;
  wire popcount45_pvta_core_267;
  wire popcount45_pvta_core_268;
  wire popcount45_pvta_core_269;
  wire popcount45_pvta_core_270;
  wire popcount45_pvta_core_271;
  wire popcount45_pvta_core_273;
  wire popcount45_pvta_core_274;
  wire popcount45_pvta_core_275;
  wire popcount45_pvta_core_276;
  wire popcount45_pvta_core_277;
  wire popcount45_pvta_core_278;
  wire popcount45_pvta_core_280;
  wire popcount45_pvta_core_281;
  wire popcount45_pvta_core_284;
  wire popcount45_pvta_core_288;
  wire popcount45_pvta_core_292;
  wire popcount45_pvta_core_295;
  wire popcount45_pvta_core_296;
  wire popcount45_pvta_core_298;
  wire popcount45_pvta_core_299;
  wire popcount45_pvta_core_303;
  wire popcount45_pvta_core_304;
  wire popcount45_pvta_core_305;
  wire popcount45_pvta_core_306;
  wire popcount45_pvta_core_308;
  wire popcount45_pvta_core_309;
  wire popcount45_pvta_core_310;
  wire popcount45_pvta_core_311;
  wire popcount45_pvta_core_315;
  wire popcount45_pvta_core_316;
  wire popcount45_pvta_core_317_not;
  wire popcount45_pvta_core_319;
  wire popcount45_pvta_core_320;
  wire popcount45_pvta_core_321;
  wire popcount45_pvta_core_322;
  wire popcount45_pvta_core_323;
  wire popcount45_pvta_core_324;
  wire popcount45_pvta_core_325;
  wire popcount45_pvta_core_326;
  wire popcount45_pvta_core_327;
  wire popcount45_pvta_core_328;
  wire popcount45_pvta_core_329;
  wire popcount45_pvta_core_332;
  wire popcount45_pvta_core_333;
  wire popcount45_pvta_core_336;
  wire popcount45_pvta_core_337;
  wire popcount45_pvta_core_338;
  wire popcount45_pvta_core_339;
  wire popcount45_pvta_core_340;
  wire popcount45_pvta_core_341;
  wire popcount45_pvta_core_342;
  wire popcount45_pvta_core_343;
  wire popcount45_pvta_core_344;
  wire popcount45_pvta_core_345;
  wire popcount45_pvta_core_346;
  wire popcount45_pvta_core_347;
  wire popcount45_pvta_core_348;
  wire popcount45_pvta_core_349;
  wire popcount45_pvta_core_350;
  wire popcount45_pvta_core_351;
  wire popcount45_pvta_core_352;
  wire popcount45_pvta_core_353;
  wire popcount45_pvta_core_354;
  wire popcount45_pvta_core_355;
  wire popcount45_pvta_core_356;

  assign popcount45_pvta_core_047 = input_a[0] ^ input_a[1];
  assign popcount45_pvta_core_049 = input_a[3] ^ input_a[4];
  assign popcount45_pvta_core_051 = input_a[2] ^ input_a[39];
  assign popcount45_pvta_core_052 = input_a[2] & popcount45_pvta_core_049;
  assign popcount45_pvta_core_055 = popcount45_pvta_core_047 | popcount45_pvta_core_051;
  assign popcount45_pvta_core_056 = popcount45_pvta_core_047 & popcount45_pvta_core_051;
  assign popcount45_pvta_core_057 = input_a[0] ^ popcount45_pvta_core_052;
  assign popcount45_pvta_core_058 = input_a[0] & popcount45_pvta_core_052;
  assign popcount45_pvta_core_059 = popcount45_pvta_core_057 ^ popcount45_pvta_core_056;
  assign popcount45_pvta_core_060 = popcount45_pvta_core_057 & popcount45_pvta_core_056;
  assign popcount45_pvta_core_061 = popcount45_pvta_core_058 | popcount45_pvta_core_060;
  assign popcount45_pvta_core_064 = input_a[6] ^ input_a[7];
  assign popcount45_pvta_core_065 = input_a[6] & input_a[7];
  assign popcount45_pvta_core_067 = input_a[5] & input_a[29];
  assign popcount45_pvta_core_068 = popcount45_pvta_core_065 ^ popcount45_pvta_core_067;
  assign popcount45_pvta_core_069 = popcount45_pvta_core_065 & popcount45_pvta_core_067;
  assign popcount45_pvta_core_070 = input_a[9] ^ input_a[10];
  assign popcount45_pvta_core_071 = input_a[9] & input_a[10];
  assign popcount45_pvta_core_072 = input_a[8] ^ popcount45_pvta_core_070;
  assign popcount45_pvta_core_073 = input_a[8] & popcount45_pvta_core_070;
  assign popcount45_pvta_core_074 = ~popcount45_pvta_core_071;
  assign popcount45_pvta_core_075 = popcount45_pvta_core_071 & popcount45_pvta_core_073;
  assign popcount45_pvta_core_078 = popcount45_pvta_core_068 ^ popcount45_pvta_core_074;
  assign popcount45_pvta_core_079 = popcount45_pvta_core_068 & popcount45_pvta_core_074;
  assign popcount45_pvta_core_083 = popcount45_pvta_core_069 ^ popcount45_pvta_core_075;
  assign popcount45_pvta_core_084 = popcount45_pvta_core_069 & popcount45_pvta_core_075;
  assign popcount45_pvta_core_085 = popcount45_pvta_core_083 & popcount45_pvta_core_079;
  assign popcount45_pvta_core_086 = popcount45_pvta_core_083 & popcount45_pvta_core_079;
  assign popcount45_pvta_core_087 = popcount45_pvta_core_084 | popcount45_pvta_core_086;
  assign popcount45_pvta_core_088 = input_a[24] ^ popcount45_pvta_core_072;
  assign popcount45_pvta_core_089 = popcount45_pvta_core_055 & popcount45_pvta_core_072;
  assign popcount45_pvta_core_090 = popcount45_pvta_core_059 ^ popcount45_pvta_core_078;
  assign popcount45_pvta_core_091 = popcount45_pvta_core_059 & popcount45_pvta_core_078;
  assign popcount45_pvta_core_092 = popcount45_pvta_core_090 ^ input_a[29];
  assign popcount45_pvta_core_093 = popcount45_pvta_core_090 & input_a[12];
  assign popcount45_pvta_core_094 = popcount45_pvta_core_091 | popcount45_pvta_core_093;
  assign popcount45_pvta_core_095 = popcount45_pvta_core_061 ^ popcount45_pvta_core_085;
  assign popcount45_pvta_core_096 = popcount45_pvta_core_061 & popcount45_pvta_core_085;
  assign popcount45_pvta_core_097 = popcount45_pvta_core_095 ^ popcount45_pvta_core_094;
  assign popcount45_pvta_core_098 = popcount45_pvta_core_095 & popcount45_pvta_core_094;
  assign popcount45_pvta_core_099 = popcount45_pvta_core_096 | popcount45_pvta_core_098;
  assign popcount45_pvta_core_101 = input_a[6] & popcount45_pvta_core_087;
  assign popcount45_pvta_core_102 = popcount45_pvta_core_087 ^ popcount45_pvta_core_099;
  assign popcount45_pvta_core_103 = popcount45_pvta_core_087 & popcount45_pvta_core_099;
  assign popcount45_pvta_core_104 = popcount45_pvta_core_101 | popcount45_pvta_core_103;
  assign popcount45_pvta_core_105 = ~(input_a[0] | input_a[12]);
  assign popcount45_pvta_core_106 = input_a[11] & input_a[12];
  assign popcount45_pvta_core_107 = ~(input_a[14] | input_a[15]);
  assign popcount45_pvta_core_108 = input_a[14] & input_a[15];
  assign popcount45_pvta_core_109 = input_a[13] ^ popcount45_pvta_core_107;
  assign popcount45_pvta_core_110 = input_a[13] & popcount45_pvta_core_107;
  assign popcount45_pvta_core_111 = ~popcount45_pvta_core_108;
  assign popcount45_pvta_core_112 = popcount45_pvta_core_108 & popcount45_pvta_core_110;
  assign popcount45_pvta_core_114 = popcount45_pvta_core_105 & input_a[31];
  assign popcount45_pvta_core_115 = popcount45_pvta_core_106 ^ popcount45_pvta_core_111;
  assign popcount45_pvta_core_116 = popcount45_pvta_core_106 & popcount45_pvta_core_111;
  assign popcount45_pvta_core_117 = input_a[30] ^ popcount45_pvta_core_114;
  assign popcount45_pvta_core_118 = popcount45_pvta_core_115 & popcount45_pvta_core_114;
  assign popcount45_pvta_core_122 = ~(input_a[17] & input_a[18]);
  assign popcount45_pvta_core_124 = input_a[25] ^ popcount45_pvta_core_122;
  assign popcount45_pvta_core_125 = ~(input_a[16] | popcount45_pvta_core_122);
  assign popcount45_pvta_core_126 = input_a[17] ^ popcount45_pvta_core_125;
  assign popcount45_pvta_core_127 = input_a[17] & popcount45_pvta_core_125;
  assign popcount45_pvta_core_128 = input_a[20] ^ input_a[21];
  assign popcount45_pvta_core_129 = input_a[20] & input_a[21];
  assign popcount45_pvta_core_134_not = ~popcount45_pvta_core_124;
  assign popcount45_pvta_core_136 = popcount45_pvta_core_126 ^ input_a[8];
  assign popcount45_pvta_core_137 = popcount45_pvta_core_126 & input_a[8];
  assign popcount45_pvta_core_138 = popcount45_pvta_core_136 ^ popcount45_pvta_core_124;
  assign popcount45_pvta_core_139 = popcount45_pvta_core_136 & popcount45_pvta_core_124;
  assign popcount45_pvta_core_140 = popcount45_pvta_core_137 | input_a[30];
  assign popcount45_pvta_core_143 = popcount45_pvta_core_127 ^ popcount45_pvta_core_140;
  assign popcount45_pvta_core_144 = popcount45_pvta_core_127 & popcount45_pvta_core_140;
  assign popcount45_pvta_core_149 = popcount45_pvta_core_117 & input_a[26];
  assign popcount45_pvta_core_152 = input_a[36] | input_a[17];
  assign popcount45_pvta_core_154 = popcount45_pvta_core_112 & popcount45_pvta_core_143;
  assign popcount45_pvta_core_155 = ~(popcount45_pvta_core_112 & popcount45_pvta_core_152);
  assign popcount45_pvta_core_156 = popcount45_pvta_core_112 & popcount45_pvta_core_152;
  assign popcount45_pvta_core_157 = popcount45_pvta_core_154 | popcount45_pvta_core_156;
  assign popcount45_pvta_core_158 = popcount45_pvta_core_112 ^ popcount45_pvta_core_144;
  assign popcount45_pvta_core_159 = popcount45_pvta_core_112 & popcount45_pvta_core_144;
  assign popcount45_pvta_core_160 = popcount45_pvta_core_158 ^ popcount45_pvta_core_157;
  assign popcount45_pvta_core_161 = popcount45_pvta_core_158 & popcount45_pvta_core_157;
  assign popcount45_pvta_core_164 = ~(input_a[24] | popcount45_pvta_core_134_not);
  assign popcount45_pvta_core_165 = input_a[31] ^ input_a[5];
  assign popcount45_pvta_core_166 = input_a[8] & input_a[5];
  assign popcount45_pvta_core_167 = input_a[29] ^ popcount45_pvta_core_164;
  assign popcount45_pvta_core_168 = popcount45_pvta_core_165 & popcount45_pvta_core_164;
  assign popcount45_pvta_core_169 = popcount45_pvta_core_166 | popcount45_pvta_core_168;
  assign popcount45_pvta_core_170 = popcount45_pvta_core_097 ^ popcount45_pvta_core_155;
  assign popcount45_pvta_core_171 = popcount45_pvta_core_097 & popcount45_pvta_core_155;
  assign popcount45_pvta_core_172 = popcount45_pvta_core_170 ^ popcount45_pvta_core_169;
  assign popcount45_pvta_core_173 = popcount45_pvta_core_170 & popcount45_pvta_core_169;
  assign popcount45_pvta_core_174 = popcount45_pvta_core_171 | popcount45_pvta_core_173;
  assign popcount45_pvta_core_175 = popcount45_pvta_core_102 ^ popcount45_pvta_core_160;
  assign popcount45_pvta_core_176 = popcount45_pvta_core_102 & popcount45_pvta_core_160;
  assign popcount45_pvta_core_177 = popcount45_pvta_core_175 ^ popcount45_pvta_core_174;
  assign popcount45_pvta_core_178 = popcount45_pvta_core_175 & popcount45_pvta_core_174;
  assign popcount45_pvta_core_179 = popcount45_pvta_core_176 | popcount45_pvta_core_178;
  assign popcount45_pvta_core_182 = popcount45_pvta_core_104 ^ popcount45_pvta_core_179;
  assign popcount45_pvta_core_183 = input_a[2] & popcount45_pvta_core_179;
  assign popcount45_pvta_core_185 = input_a[22] ^ input_a[23];
  assign popcount45_pvta_core_186 = input_a[22] & input_a[23];
  assign popcount45_pvta_core_189 = input_a[24] ^ input_a[5];
  assign popcount45_pvta_core_193 = popcount45_pvta_core_185 ^ popcount45_pvta_core_189;
  assign popcount45_pvta_core_194 = popcount45_pvta_core_185 & popcount45_pvta_core_189;
  assign popcount45_pvta_core_195 = popcount45_pvta_core_186 ^ input_a[24];
  assign popcount45_pvta_core_196 = popcount45_pvta_core_186 & input_a[24];
  assign popcount45_pvta_core_197 = popcount45_pvta_core_195 ^ popcount45_pvta_core_194;
  assign popcount45_pvta_core_198 = popcount45_pvta_core_195 & popcount45_pvta_core_194;
  assign popcount45_pvta_core_199 = input_a[24] | input_a[33];
  assign popcount45_pvta_core_203 = input_a[28] & input_a[29];
  assign popcount45_pvta_core_204 = ~input_a[27];
  assign popcount45_pvta_core_206 = popcount45_pvta_core_203 ^ input_a[27];
  assign popcount45_pvta_core_207 = popcount45_pvta_core_203 & input_a[28];
  assign popcount45_pvta_core_208 = ~(input_a[31] | input_a[32]);
  assign popcount45_pvta_core_209 = input_a[5] & input_a[32];
  assign popcount45_pvta_core_211 = input_a[30] & popcount45_pvta_core_208;
  assign popcount45_pvta_core_212 = popcount45_pvta_core_209 ^ popcount45_pvta_core_211;
  assign popcount45_pvta_core_213 = input_a[43] & popcount45_pvta_core_211;
  assign popcount45_pvta_core_214_not = ~popcount45_pvta_core_204;
  assign popcount45_pvta_core_216 = ~(popcount45_pvta_core_206 & popcount45_pvta_core_212);
  assign popcount45_pvta_core_217 = popcount45_pvta_core_206 & input_a[24];
  assign popcount45_pvta_core_219 = popcount45_pvta_core_216 & popcount45_pvta_core_204;
  assign popcount45_pvta_core_220 = popcount45_pvta_core_217 | input_a[36];
  assign popcount45_pvta_core_221 = popcount45_pvta_core_207 ^ popcount45_pvta_core_213;
  assign popcount45_pvta_core_222 = popcount45_pvta_core_207 & popcount45_pvta_core_213;
  assign popcount45_pvta_core_223 = ~(popcount45_pvta_core_221 & popcount45_pvta_core_220);
  assign popcount45_pvta_core_224 = popcount45_pvta_core_221 & popcount45_pvta_core_220;
  assign popcount45_pvta_core_225 = popcount45_pvta_core_222 | popcount45_pvta_core_224;
  assign popcount45_pvta_core_226 = popcount45_pvta_core_193 ^ popcount45_pvta_core_214_not;
  assign popcount45_pvta_core_227 = ~popcount45_pvta_core_193;
  assign popcount45_pvta_core_228_not = ~popcount45_pvta_core_197;
  assign popcount45_pvta_core_230 = popcount45_pvta_core_228_not ^ popcount45_pvta_core_227;
  assign popcount45_pvta_core_231 = popcount45_pvta_core_228_not & popcount45_pvta_core_227;
  assign popcount45_pvta_core_232 = input_a[30] | popcount45_pvta_core_231;
  assign popcount45_pvta_core_233_not = ~popcount45_pvta_core_223;
  assign popcount45_pvta_core_234 = input_a[32] & popcount45_pvta_core_223;
  assign popcount45_pvta_core_235 = popcount45_pvta_core_233_not ^ popcount45_pvta_core_232;
  assign popcount45_pvta_core_236 = popcount45_pvta_core_233_not & popcount45_pvta_core_232;
  assign popcount45_pvta_core_237 = popcount45_pvta_core_234 | popcount45_pvta_core_236;
  assign popcount45_pvta_core_240 = popcount45_pvta_core_225 ^ popcount45_pvta_core_237;
  assign popcount45_pvta_core_241 = popcount45_pvta_core_225 & popcount45_pvta_core_237;
  assign popcount45_pvta_core_243 = input_a[23] ^ input_a[35];
  assign popcount45_pvta_core_245 = ~(input_a[33] & popcount45_pvta_core_243);
  assign popcount45_pvta_core_246 = input_a[33] & popcount45_pvta_core_243;
  assign popcount45_pvta_core_249 = input_a[37] ^ input_a[38];
  assign popcount45_pvta_core_250 = input_a[37] & input_a[38];
  assign popcount45_pvta_core_251 = ~(input_a[36] | popcount45_pvta_core_249);
  assign popcount45_pvta_core_252 = input_a[24] & input_a[13];
  assign popcount45_pvta_core_253 = popcount45_pvta_core_250 ^ popcount45_pvta_core_252;
  assign popcount45_pvta_core_254 = popcount45_pvta_core_250 & popcount45_pvta_core_252;
  assign popcount45_pvta_core_255 = ~popcount45_pvta_core_245;
  assign popcount45_pvta_core_256 = input_a[33] & input_a[35];
  assign popcount45_pvta_core_259 = popcount45_pvta_core_253 ^ popcount45_pvta_core_256;
  assign popcount45_pvta_core_260 = input_a[0] & popcount45_pvta_core_256;
  assign popcount45_pvta_core_264 = input_a[11] ^ input_a[27];
  assign popcount45_pvta_core_265 = popcount45_pvta_core_254 & input_a[27];
  assign popcount45_pvta_core_267 = input_a[40] ^ input_a[41];
  assign popcount45_pvta_core_268 = input_a[40] & input_a[41];
  assign popcount45_pvta_core_269 = input_a[39] ^ popcount45_pvta_core_267;
  assign popcount45_pvta_core_270 = input_a[39] & popcount45_pvta_core_267;
  assign popcount45_pvta_core_271 = popcount45_pvta_core_268 ^ popcount45_pvta_core_270;
  assign popcount45_pvta_core_273 = input_a[43] ^ input_a[44];
  assign popcount45_pvta_core_274 = input_a[43] & input_a[44];
  assign popcount45_pvta_core_275 = input_a[42] ^ popcount45_pvta_core_273;
  assign popcount45_pvta_core_276 = input_a[30] & popcount45_pvta_core_273;
  assign popcount45_pvta_core_277 = input_a[27] ^ input_a[39];
  assign popcount45_pvta_core_278 = popcount45_pvta_core_274 & popcount45_pvta_core_276;
  assign popcount45_pvta_core_280 = popcount45_pvta_core_269 & popcount45_pvta_core_275;
  assign popcount45_pvta_core_281 = popcount45_pvta_core_271 ^ popcount45_pvta_core_277;
  assign popcount45_pvta_core_284 = popcount45_pvta_core_281 & popcount45_pvta_core_280;
  assign popcount45_pvta_core_288 = popcount45_pvta_core_278 | input_a[38];
  assign popcount45_pvta_core_292 = popcount45_pvta_core_255 & input_a[15];
  assign popcount45_pvta_core_295 = input_a[8] | popcount45_pvta_core_292;
  assign popcount45_pvta_core_296 = ~input_a[3];
  assign popcount45_pvta_core_298 = popcount45_pvta_core_264 ^ popcount45_pvta_core_288;
  assign popcount45_pvta_core_299 = popcount45_pvta_core_264 & popcount45_pvta_core_288;
  assign popcount45_pvta_core_303 = popcount45_pvta_core_265 ^ popcount45_pvta_core_278;
  assign popcount45_pvta_core_304 = popcount45_pvta_core_265 & popcount45_pvta_core_278;
  assign popcount45_pvta_core_305 = popcount45_pvta_core_303 ^ popcount45_pvta_core_299;
  assign popcount45_pvta_core_306 = popcount45_pvta_core_303 & popcount45_pvta_core_299;
  assign popcount45_pvta_core_308 = popcount45_pvta_core_226 & popcount45_pvta_core_255;
  assign popcount45_pvta_core_309 = popcount45_pvta_core_226 & popcount45_pvta_core_255;
  assign popcount45_pvta_core_310 = popcount45_pvta_core_230 ^ popcount45_pvta_core_295;
  assign popcount45_pvta_core_311 = popcount45_pvta_core_230 & popcount45_pvta_core_295;
  assign popcount45_pvta_core_315 = input_a[1] ^ input_a[11];
  assign popcount45_pvta_core_316 = popcount45_pvta_core_235 & input_a[11];
  assign popcount45_pvta_core_317_not = ~popcount45_pvta_core_315;
  assign popcount45_pvta_core_319 = ~popcount45_pvta_core_316;
  assign popcount45_pvta_core_320 = popcount45_pvta_core_240 ^ popcount45_pvta_core_305;
  assign popcount45_pvta_core_321 = popcount45_pvta_core_240 & popcount45_pvta_core_305;
  assign popcount45_pvta_core_322 = popcount45_pvta_core_320 ^ popcount45_pvta_core_319;
  assign popcount45_pvta_core_323 = popcount45_pvta_core_320 & popcount45_pvta_core_319;
  assign popcount45_pvta_core_324 = popcount45_pvta_core_321 | popcount45_pvta_core_323;
  assign popcount45_pvta_core_325 = popcount45_pvta_core_241 | popcount45_pvta_core_304;
  assign popcount45_pvta_core_326 = popcount45_pvta_core_241 & popcount45_pvta_core_304;
  assign popcount45_pvta_core_327 = popcount45_pvta_core_325 ^ popcount45_pvta_core_324;
  assign popcount45_pvta_core_328 = popcount45_pvta_core_325 & popcount45_pvta_core_324;
  assign popcount45_pvta_core_329 = popcount45_pvta_core_326 | popcount45_pvta_core_328;
  assign popcount45_pvta_core_332 = popcount45_pvta_core_167 ^ popcount45_pvta_core_310;
  assign popcount45_pvta_core_333 = ~(popcount45_pvta_core_167 & popcount45_pvta_core_310);
  assign popcount45_pvta_core_336 = input_a[44] & input_a[26];
  assign popcount45_pvta_core_337 = popcount45_pvta_core_172 ^ popcount45_pvta_core_317_not;
  assign popcount45_pvta_core_338 = popcount45_pvta_core_172 & popcount45_pvta_core_317_not;
  assign popcount45_pvta_core_339 = input_a[7] ^ popcount45_pvta_core_336;
  assign popcount45_pvta_core_340 = popcount45_pvta_core_337 & popcount45_pvta_core_336;
  assign popcount45_pvta_core_341 = popcount45_pvta_core_338 | input_a[38];
  assign popcount45_pvta_core_342 = popcount45_pvta_core_177 ^ popcount45_pvta_core_322;
  assign popcount45_pvta_core_343 = input_a[3] & popcount45_pvta_core_322;
  assign popcount45_pvta_core_344 = popcount45_pvta_core_342 ^ popcount45_pvta_core_341;
  assign popcount45_pvta_core_345 = popcount45_pvta_core_342 & popcount45_pvta_core_341;
  assign popcount45_pvta_core_346 = popcount45_pvta_core_343 | popcount45_pvta_core_345;
  assign popcount45_pvta_core_347 = popcount45_pvta_core_182 ^ popcount45_pvta_core_327;
  assign popcount45_pvta_core_348 = popcount45_pvta_core_182 & popcount45_pvta_core_327;
  assign popcount45_pvta_core_349 = ~(popcount45_pvta_core_347 & popcount45_pvta_core_346);
  assign popcount45_pvta_core_350 = popcount45_pvta_core_347 & popcount45_pvta_core_346;
  assign popcount45_pvta_core_351 = popcount45_pvta_core_348 | popcount45_pvta_core_350;
  assign popcount45_pvta_core_352 = popcount45_pvta_core_183 ^ popcount45_pvta_core_329;
  assign popcount45_pvta_core_353 = popcount45_pvta_core_183 & popcount45_pvta_core_329;
  assign popcount45_pvta_core_354 = popcount45_pvta_core_352 ^ popcount45_pvta_core_351;
  assign popcount45_pvta_core_355 = popcount45_pvta_core_352 & popcount45_pvta_core_351;
  assign popcount45_pvta_core_356 = popcount45_pvta_core_353 | popcount45_pvta_core_355;

  assign popcount45_pvta_out[0] = popcount45_pvta_core_308;
  assign popcount45_pvta_out[1] = popcount45_pvta_core_332;
  assign popcount45_pvta_out[2] = popcount45_pvta_core_339;
  assign popcount45_pvta_out[3] = popcount45_pvta_core_344;
  assign popcount45_pvta_out[4] = popcount45_pvta_core_349;
  assign popcount45_pvta_out[5] = popcount45_pvta_core_354;
endmodule