// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.41533
// WCE=12.0
// EP=0.875124%
// Printed PDK parameters:
//  Area=1576580.0
//  Delay=5889130.5
//  Power=61525.0

module popcount23_053y(input [22:0] input_a, output [4:0] popcount23_053y_out);
  wire popcount23_053y_core_025;
  wire popcount23_053y_core_026;
  wire popcount23_053y_core_027;
  wire popcount23_053y_core_028;
  wire popcount23_053y_core_030;
  wire popcount23_053y_core_032;
  wire popcount23_053y_core_034;
  wire popcount23_053y_core_035;
  wire popcount23_053y_core_038;
  wire popcount23_053y_core_039;
  wire popcount23_053y_core_040;
  wire popcount23_053y_core_042;
  wire popcount23_053y_core_043;
  wire popcount23_053y_core_044;
  wire popcount23_053y_core_045;
  wire popcount23_053y_core_046;
  wire popcount23_053y_core_047;
  wire popcount23_053y_core_049;
  wire popcount23_053y_core_052;
  wire popcount23_053y_core_054;
  wire popcount23_053y_core_055;
  wire popcount23_053y_core_056_not;
  wire popcount23_053y_core_061;
  wire popcount23_053y_core_063;
  wire popcount23_053y_core_068_not;
  wire popcount23_053y_core_070;
  wire popcount23_053y_core_072;
  wire popcount23_053y_core_073;
  wire popcount23_053y_core_076;
  wire popcount23_053y_core_078;
  wire popcount23_053y_core_080;
  wire popcount23_053y_core_081;
  wire popcount23_053y_core_084;
  wire popcount23_053y_core_088;
  wire popcount23_053y_core_089;
  wire popcount23_053y_core_090;
  wire popcount23_053y_core_091;
  wire popcount23_053y_core_092;
  wire popcount23_053y_core_093;
  wire popcount23_053y_core_094;
  wire popcount23_053y_core_095;
  wire popcount23_053y_core_096;
  wire popcount23_053y_core_097;
  wire popcount23_053y_core_098;
  wire popcount23_053y_core_099;
  wire popcount23_053y_core_100;
  wire popcount23_053y_core_102;
  wire popcount23_053y_core_103;
  wire popcount23_053y_core_104;
  wire popcount23_053y_core_105;
  wire popcount23_053y_core_106;
  wire popcount23_053y_core_107;
  wire popcount23_053y_core_108;
  wire popcount23_053y_core_110;
  wire popcount23_053y_core_111;
  wire popcount23_053y_core_113;
  wire popcount23_053y_core_114;
  wire popcount23_053y_core_115;
  wire popcount23_053y_core_116;
  wire popcount23_053y_core_117;
  wire popcount23_053y_core_118;
  wire popcount23_053y_core_119;
  wire popcount23_053y_core_120;
  wire popcount23_053y_core_121;
  wire popcount23_053y_core_126;
  wire popcount23_053y_core_128;
  wire popcount23_053y_core_134;
  wire popcount23_053y_core_136;
  wire popcount23_053y_core_137;
  wire popcount23_053y_core_138;
  wire popcount23_053y_core_144;
  wire popcount23_053y_core_145;
  wire popcount23_053y_core_146;
  wire popcount23_053y_core_147;
  wire popcount23_053y_core_150;
  wire popcount23_053y_core_154;
  wire popcount23_053y_core_155_not;
  wire popcount23_053y_core_157;
  wire popcount23_053y_core_159_not;
  wire popcount23_053y_core_160;
  wire popcount23_053y_core_161;
  wire popcount23_053y_core_162;
  wire popcount23_053y_core_163;
  wire popcount23_053y_core_164;
  wire popcount23_053y_core_165;
  wire popcount23_053y_core_166;
  wire popcount23_053y_core_168;
  wire popcount23_053y_core_169;

  assign popcount23_053y_core_025 = input_a[17] ^ input_a[19];
  assign popcount23_053y_core_026 = ~(input_a[5] ^ input_a[0]);
  assign popcount23_053y_core_027 = input_a[2] & input_a[17];
  assign popcount23_053y_core_028 = ~input_a[2];
  assign popcount23_053y_core_030 = input_a[2] & input_a[2];
  assign popcount23_053y_core_032 = input_a[21] & input_a[10];
  assign popcount23_053y_core_034 = ~(input_a[9] & input_a[18]);
  assign popcount23_053y_core_035 = input_a[21] & input_a[1];
  assign popcount23_053y_core_038 = input_a[20] ^ input_a[0];
  assign popcount23_053y_core_039 = ~(input_a[20] | input_a[16]);
  assign popcount23_053y_core_040 = input_a[16] & input_a[14];
  assign popcount23_053y_core_042 = ~(input_a[8] ^ input_a[18]);
  assign popcount23_053y_core_043 = input_a[10] & input_a[6];
  assign popcount23_053y_core_044 = ~(input_a[9] | input_a[20]);
  assign popcount23_053y_core_045 = input_a[21] & input_a[18];
  assign popcount23_053y_core_046 = popcount23_053y_core_043 | popcount23_053y_core_045;
  assign popcount23_053y_core_047 = input_a[2] & input_a[3];
  assign popcount23_053y_core_049 = ~input_a[15];
  assign popcount23_053y_core_052 = ~(input_a[2] | input_a[0]);
  assign popcount23_053y_core_054 = ~(input_a[21] ^ input_a[12]);
  assign popcount23_053y_core_055 = ~(input_a[12] ^ input_a[6]);
  assign popcount23_053y_core_056_not = ~input_a[18];
  assign popcount23_053y_core_061 = input_a[5] | input_a[2];
  assign popcount23_053y_core_063 = input_a[1] | popcount23_053y_core_046;
  assign popcount23_053y_core_068_not = ~input_a[9];
  assign popcount23_053y_core_070 = input_a[18] | input_a[12];
  assign popcount23_053y_core_072 = ~(input_a[13] & input_a[10]);
  assign popcount23_053y_core_073 = input_a[9] | popcount23_053y_core_063;
  assign popcount23_053y_core_076 = ~(input_a[1] & input_a[1]);
  assign popcount23_053y_core_078 = ~(input_a[17] & input_a[20]);
  assign popcount23_053y_core_080 = input_a[13] ^ input_a[3];
  assign popcount23_053y_core_081 = input_a[13] ^ input_a[1];
  assign popcount23_053y_core_084 = ~(input_a[11] & input_a[17]);
  assign popcount23_053y_core_088 = input_a[7] ^ input_a[20];
  assign popcount23_053y_core_089 = ~(input_a[15] ^ input_a[9]);
  assign popcount23_053y_core_090 = input_a[20] ^ input_a[1];
  assign popcount23_053y_core_091 = ~(input_a[13] ^ input_a[0]);
  assign popcount23_053y_core_092 = ~input_a[22];
  assign popcount23_053y_core_093 = ~(input_a[6] ^ input_a[8]);
  assign popcount23_053y_core_094 = ~(input_a[20] ^ input_a[22]);
  assign popcount23_053y_core_095 = input_a[2] | input_a[9];
  assign popcount23_053y_core_096 = ~input_a[18];
  assign popcount23_053y_core_097 = ~input_a[1];
  assign popcount23_053y_core_098 = input_a[12] | input_a[13];
  assign popcount23_053y_core_099 = ~(input_a[7] & input_a[20]);
  assign popcount23_053y_core_100 = ~(input_a[11] ^ input_a[8]);
  assign popcount23_053y_core_102 = ~(input_a[1] ^ input_a[19]);
  assign popcount23_053y_core_103 = ~(input_a[21] & input_a[11]);
  assign popcount23_053y_core_104 = ~input_a[7];
  assign popcount23_053y_core_105 = input_a[9] | input_a[1];
  assign popcount23_053y_core_106 = ~(input_a[14] ^ input_a[6]);
  assign popcount23_053y_core_107 = ~(input_a[9] ^ input_a[12]);
  assign popcount23_053y_core_108 = ~(input_a[13] & input_a[11]);
  assign popcount23_053y_core_110 = input_a[16] | input_a[13];
  assign popcount23_053y_core_111 = input_a[11] | input_a[13];
  assign popcount23_053y_core_113 = input_a[16] | input_a[0];
  assign popcount23_053y_core_114 = ~(input_a[14] | input_a[18]);
  assign popcount23_053y_core_115 = ~(input_a[0] ^ input_a[9]);
  assign popcount23_053y_core_116 = ~(input_a[0] ^ input_a[20]);
  assign popcount23_053y_core_117 = input_a[17] ^ input_a[16];
  assign popcount23_053y_core_118 = ~(input_a[7] ^ input_a[6]);
  assign popcount23_053y_core_119 = ~(input_a[9] | input_a[14]);
  assign popcount23_053y_core_120 = ~(input_a[18] & input_a[21]);
  assign popcount23_053y_core_121 = input_a[12] & input_a[13];
  assign popcount23_053y_core_126 = ~input_a[18];
  assign popcount23_053y_core_128 = input_a[21] ^ input_a[4];
  assign popcount23_053y_core_134 = ~input_a[0];
  assign popcount23_053y_core_136 = input_a[22] & input_a[15];
  assign popcount23_053y_core_137 = input_a[7] & input_a[8];
  assign popcount23_053y_core_138 = ~(input_a[6] & input_a[20]);
  assign popcount23_053y_core_144 = input_a[20] ^ input_a[11];
  assign popcount23_053y_core_145 = ~(input_a[9] | input_a[1]);
  assign popcount23_053y_core_146 = input_a[3] ^ input_a[10];
  assign popcount23_053y_core_147 = input_a[12] ^ input_a[2];
  assign popcount23_053y_core_150 = ~input_a[19];
  assign popcount23_053y_core_154 = ~input_a[15];
  assign popcount23_053y_core_155_not = ~input_a[10];
  assign popcount23_053y_core_157 = ~input_a[2];
  assign popcount23_053y_core_159_not = ~input_a[20];
  assign popcount23_053y_core_160 = ~(input_a[10] | input_a[0]);
  assign popcount23_053y_core_161 = ~(input_a[9] ^ input_a[15]);
  assign popcount23_053y_core_162 = ~(input_a[15] ^ input_a[22]);
  assign popcount23_053y_core_163 = ~(input_a[9] | input_a[6]);
  assign popcount23_053y_core_164 = ~(input_a[3] & input_a[4]);
  assign popcount23_053y_core_165 = ~(input_a[18] & input_a[5]);
  assign popcount23_053y_core_166 = ~input_a[4];
  assign popcount23_053y_core_168 = input_a[13] ^ input_a[21];
  assign popcount23_053y_core_169 = ~input_a[18];

  assign popcount23_053y_out[0] = input_a[14];
  assign popcount23_053y_out[1] = 1'b1;
  assign popcount23_053y_out[2] = popcount23_053y_core_145;
  assign popcount23_053y_out[3] = popcount23_053y_core_073;
  assign popcount23_053y_out[4] = 1'b0;
endmodule