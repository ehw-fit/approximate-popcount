// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.17559
// WCE=16.0
// EP=0.991379%
// Printed PDK parameters:
//  Area=25471038.0
//  Delay=32281666.0
//  Power=1068000.0

module popcount31_4js4(input [30:0] input_a, output [4:0] popcount31_4js4_out);
  wire popcount31_4js4_core_033;
  wire popcount31_4js4_core_034;
  wire popcount31_4js4_core_035;
  wire popcount31_4js4_core_037;
  wire popcount31_4js4_core_038;
  wire popcount31_4js4_core_040;
  wire popcount31_4js4_core_041;
  wire popcount31_4js4_core_042;
  wire popcount31_4js4_core_044;
  wire popcount31_4js4_core_045;
  wire popcount31_4js4_core_046;
  wire popcount31_4js4_core_048;
  wire popcount31_4js4_core_049;
  wire popcount31_4js4_core_051;
  wire popcount31_4js4_core_052;
  wire popcount31_4js4_core_053;
  wire popcount31_4js4_core_055;
  wire popcount31_4js4_core_056;
  wire popcount31_4js4_core_060;
  wire popcount31_4js4_core_062;
  wire popcount31_4js4_core_063;
  wire popcount31_4js4_core_064;
  wire popcount31_4js4_core_065;
  wire popcount31_4js4_core_066;
  wire popcount31_4js4_core_067;
  wire popcount31_4js4_core_068;
  wire popcount31_4js4_core_069;
  wire popcount31_4js4_core_073;
  wire popcount31_4js4_core_074;
  wire popcount31_4js4_core_075;
  wire popcount31_4js4_core_076;
  wire popcount31_4js4_core_077;
  wire popcount31_4js4_core_079;
  wire popcount31_4js4_core_080;
  wire popcount31_4js4_core_082;
  wire popcount31_4js4_core_084;
  wire popcount31_4js4_core_085;
  wire popcount31_4js4_core_086;
  wire popcount31_4js4_core_087;
  wire popcount31_4js4_core_089;
  wire popcount31_4js4_core_090;
  wire popcount31_4js4_core_091;
  wire popcount31_4js4_core_092;
  wire popcount31_4js4_core_093;
  wire popcount31_4js4_core_096;
  wire popcount31_4js4_core_099;
  wire popcount31_4js4_core_101;
  wire popcount31_4js4_core_103;
  wire popcount31_4js4_core_104;
  wire popcount31_4js4_core_105;
  wire popcount31_4js4_core_106;
  wire popcount31_4js4_core_107;
  wire popcount31_4js4_core_109;
  wire popcount31_4js4_core_110;
  wire popcount31_4js4_core_112;
  wire popcount31_4js4_core_114;
  wire popcount31_4js4_core_115;
  wire popcount31_4js4_core_117;
  wire popcount31_4js4_core_120;
  wire popcount31_4js4_core_121;
  wire popcount31_4js4_core_122;
  wire popcount31_4js4_core_123;
  wire popcount31_4js4_core_125;
  wire popcount31_4js4_core_126;
  wire popcount31_4js4_core_127;
  wire popcount31_4js4_core_129;
  wire popcount31_4js4_core_131;
  wire popcount31_4js4_core_133;
  wire popcount31_4js4_core_134;
  wire popcount31_4js4_core_135;
  wire popcount31_4js4_core_138;
  wire popcount31_4js4_core_139;
  wire popcount31_4js4_core_141;
  wire popcount31_4js4_core_143;
  wire popcount31_4js4_core_145;
  wire popcount31_4js4_core_146;
  wire popcount31_4js4_core_149;
  wire popcount31_4js4_core_153;
  wire popcount31_4js4_core_155;
  wire popcount31_4js4_core_156;
  wire popcount31_4js4_core_158;
  wire popcount31_4js4_core_161;
  wire popcount31_4js4_core_162;
  wire popcount31_4js4_core_166;
  wire popcount31_4js4_core_169_not;
  wire popcount31_4js4_core_170;
  wire popcount31_4js4_core_171;
  wire popcount31_4js4_core_172;
  wire popcount31_4js4_core_173;
  wire popcount31_4js4_core_174;
  wire popcount31_4js4_core_177;
  wire popcount31_4js4_core_178;
  wire popcount31_4js4_core_179;
  wire popcount31_4js4_core_182_not;
  wire popcount31_4js4_core_183;
  wire popcount31_4js4_core_184;
  wire popcount31_4js4_core_186;
  wire popcount31_4js4_core_187;
  wire popcount31_4js4_core_188;
  wire popcount31_4js4_core_189;
  wire popcount31_4js4_core_190;
  wire popcount31_4js4_core_191;
  wire popcount31_4js4_core_192;
  wire popcount31_4js4_core_196;
  wire popcount31_4js4_core_197;
  wire popcount31_4js4_core_198;
  wire popcount31_4js4_core_199;
  wire popcount31_4js4_core_201;
  wire popcount31_4js4_core_202;
  wire popcount31_4js4_core_203;
  wire popcount31_4js4_core_204;
  wire popcount31_4js4_core_205;
  wire popcount31_4js4_core_206;
  wire popcount31_4js4_core_208;
  wire popcount31_4js4_core_210;
  wire popcount31_4js4_core_211;
  wire popcount31_4js4_core_212;
  wire popcount31_4js4_core_213;
  wire popcount31_4js4_core_214;
  wire popcount31_4js4_core_215;
  wire popcount31_4js4_core_217;
  wire popcount31_4js4_core_219;

  assign popcount31_4js4_core_033 = input_a[19] & input_a[5];
  assign popcount31_4js4_core_034 = ~(input_a[2] & input_a[18]);
  assign popcount31_4js4_core_035 = input_a[16] & input_a[8];
  assign popcount31_4js4_core_037 = input_a[24] | input_a[10];
  assign popcount31_4js4_core_038 = ~(input_a[22] | input_a[26]);
  assign popcount31_4js4_core_040 = input_a[5] & input_a[30];
  assign popcount31_4js4_core_041 = ~(input_a[25] & input_a[15]);
  assign popcount31_4js4_core_042 = input_a[22] & input_a[6];
  assign popcount31_4js4_core_044 = input_a[11] | input_a[21];
  assign popcount31_4js4_core_045 = popcount31_4js4_core_040 | popcount31_4js4_core_042;
  assign popcount31_4js4_core_046 = ~(input_a[1] | input_a[4]);
  assign popcount31_4js4_core_048 = input_a[7] | input_a[20];
  assign popcount31_4js4_core_049 = input_a[10] & input_a[17];
  assign popcount31_4js4_core_051 = input_a[23] & input_a[9];
  assign popcount31_4js4_core_052 = input_a[14] & input_a[16];
  assign popcount31_4js4_core_053 = popcount31_4js4_core_037 & popcount31_4js4_core_045;
  assign popcount31_4js4_core_055 = input_a[26] & popcount31_4js4_core_051;
  assign popcount31_4js4_core_056 = popcount31_4js4_core_053 | popcount31_4js4_core_055;
  assign popcount31_4js4_core_060 = input_a[4] & input_a[28];
  assign popcount31_4js4_core_062 = ~(input_a[19] | input_a[24]);
  assign popcount31_4js4_core_063 = input_a[17] & input_a[20];
  assign popcount31_4js4_core_064 = input_a[15] & input_a[12];
  assign popcount31_4js4_core_065 = input_a[1] & input_a[3];
  assign popcount31_4js4_core_066 = ~input_a[8];
  assign popcount31_4js4_core_067 = input_a[22] ^ input_a[13];
  assign popcount31_4js4_core_068 = popcount31_4js4_core_063 ^ popcount31_4js4_core_065;
  assign popcount31_4js4_core_069 = popcount31_4js4_core_063 & popcount31_4js4_core_065;
  assign popcount31_4js4_core_073 = input_a[11] ^ input_a[12];
  assign popcount31_4js4_core_074 = input_a[11] & input_a[12];
  assign popcount31_4js4_core_075 = input_a[13] ^ input_a[14];
  assign popcount31_4js4_core_076 = input_a[13] & input_a[14];
  assign popcount31_4js4_core_077 = popcount31_4js4_core_073 | popcount31_4js4_core_075;
  assign popcount31_4js4_core_079 = popcount31_4js4_core_074 ^ popcount31_4js4_core_076;
  assign popcount31_4js4_core_080 = popcount31_4js4_core_074 & popcount31_4js4_core_076;
  assign popcount31_4js4_core_082 = ~(input_a[27] & input_a[9]);
  assign popcount31_4js4_core_084 = ~(input_a[23] ^ input_a[2]);
  assign popcount31_4js4_core_085 = input_a[4] & popcount31_4js4_core_077;
  assign popcount31_4js4_core_086 = popcount31_4js4_core_068 | popcount31_4js4_core_079;
  assign popcount31_4js4_core_087 = popcount31_4js4_core_068 & popcount31_4js4_core_079;
  assign popcount31_4js4_core_089 = input_a[0] & popcount31_4js4_core_085;
  assign popcount31_4js4_core_090 = popcount31_4js4_core_087 | popcount31_4js4_core_089;
  assign popcount31_4js4_core_091 = popcount31_4js4_core_069 ^ popcount31_4js4_core_080;
  assign popcount31_4js4_core_092 = popcount31_4js4_core_069 & popcount31_4js4_core_080;
  assign popcount31_4js4_core_093 = popcount31_4js4_core_091 | popcount31_4js4_core_090;
  assign popcount31_4js4_core_096 = ~(input_a[17] ^ input_a[5]);
  assign popcount31_4js4_core_099 = input_a[15] & popcount31_4js4_core_086;
  assign popcount31_4js4_core_101 = input_a[4] & input_a[26];
  assign popcount31_4js4_core_103 = popcount31_4js4_core_056 ^ popcount31_4js4_core_093;
  assign popcount31_4js4_core_104 = popcount31_4js4_core_056 & popcount31_4js4_core_093;
  assign popcount31_4js4_core_105 = popcount31_4js4_core_103 ^ popcount31_4js4_core_099;
  assign popcount31_4js4_core_106 = popcount31_4js4_core_103 & popcount31_4js4_core_099;
  assign popcount31_4js4_core_107 = popcount31_4js4_core_104 | popcount31_4js4_core_106;
  assign popcount31_4js4_core_109 = input_a[0] & input_a[10];
  assign popcount31_4js4_core_110 = popcount31_4js4_core_092 | popcount31_4js4_core_107;
  assign popcount31_4js4_core_112 = ~(input_a[29] ^ input_a[23]);
  assign popcount31_4js4_core_114 = ~(input_a[23] ^ input_a[22]);
  assign popcount31_4js4_core_115 = ~input_a[30];
  assign popcount31_4js4_core_117 = ~input_a[25];
  assign popcount31_4js4_core_120 = input_a[8] | input_a[20];
  assign popcount31_4js4_core_121 = ~(input_a[12] ^ input_a[28]);
  assign popcount31_4js4_core_122 = input_a[5] & input_a[6];
  assign popcount31_4js4_core_123 = ~(input_a[4] | input_a[26]);
  assign popcount31_4js4_core_125 = ~input_a[27];
  assign popcount31_4js4_core_126 = ~(input_a[18] ^ input_a[4]);
  assign popcount31_4js4_core_127 = ~(input_a[4] & input_a[16]);
  assign popcount31_4js4_core_129 = input_a[25] ^ input_a[4];
  assign popcount31_4js4_core_131 = ~(input_a[16] ^ input_a[20]);
  assign popcount31_4js4_core_133 = ~(input_a[29] & input_a[23]);
  assign popcount31_4js4_core_134 = ~input_a[0];
  assign popcount31_4js4_core_135 = ~(input_a[11] & input_a[27]);
  assign popcount31_4js4_core_138 = input_a[19] & input_a[21];
  assign popcount31_4js4_core_139 = ~input_a[7];
  assign popcount31_4js4_core_141 = popcount31_4js4_core_138 | popcount31_4js4_core_117;
  assign popcount31_4js4_core_143 = ~input_a[21];
  assign popcount31_4js4_core_145 = ~(input_a[17] | input_a[21]);
  assign popcount31_4js4_core_146 = input_a[8] & input_a[16];
  assign popcount31_4js4_core_149 = input_a[26] ^ input_a[5];
  assign popcount31_4js4_core_153 = ~(input_a[18] ^ input_a[2]);
  assign popcount31_4js4_core_155 = input_a[28] | input_a[7];
  assign popcount31_4js4_core_156 = input_a[24] ^ input_a[10];
  assign popcount31_4js4_core_158 = ~(input_a[15] ^ input_a[2]);
  assign popcount31_4js4_core_161 = input_a[8] & input_a[27];
  assign popcount31_4js4_core_162 = input_a[24] ^ input_a[9];
  assign popcount31_4js4_core_166 = input_a[29] | input_a[16];
  assign popcount31_4js4_core_169_not = ~input_a[18];
  assign popcount31_4js4_core_170 = ~(input_a[11] ^ input_a[23]);
  assign popcount31_4js4_core_171 = ~(input_a[11] ^ input_a[6]);
  assign popcount31_4js4_core_172 = popcount31_4js4_core_155 & popcount31_4js4_core_166;
  assign popcount31_4js4_core_173 = input_a[20] | input_a[18];
  assign popcount31_4js4_core_174 = ~(input_a[26] & input_a[8]);
  assign popcount31_4js4_core_177 = ~(input_a[25] | input_a[21]);
  assign popcount31_4js4_core_178 = popcount31_4js4_core_161 | popcount31_4js4_core_172;
  assign popcount31_4js4_core_179 = ~input_a[2];
  assign popcount31_4js4_core_182_not = ~input_a[19];
  assign popcount31_4js4_core_183 = ~input_a[10];
  assign popcount31_4js4_core_184 = input_a[3] ^ input_a[15];
  assign popcount31_4js4_core_186 = input_a[3] ^ input_a[27];
  assign popcount31_4js4_core_187 = input_a[2] | input_a[18];
  assign popcount31_4js4_core_188 = popcount31_4js4_core_141 ^ popcount31_4js4_core_178;
  assign popcount31_4js4_core_189 = popcount31_4js4_core_141 & popcount31_4js4_core_178;
  assign popcount31_4js4_core_190 = popcount31_4js4_core_188 ^ popcount31_4js4_core_187;
  assign popcount31_4js4_core_191 = popcount31_4js4_core_188 & popcount31_4js4_core_187;
  assign popcount31_4js4_core_192 = popcount31_4js4_core_189 | popcount31_4js4_core_191;
  assign popcount31_4js4_core_196 = ~(input_a[28] | input_a[9]);
  assign popcount31_4js4_core_197 = input_a[17] ^ input_a[19];
  assign popcount31_4js4_core_198 = ~(input_a[25] | input_a[3]);
  assign popcount31_4js4_core_199 = input_a[30] ^ input_a[25];
  assign popcount31_4js4_core_201 = input_a[23] | input_a[16];
  assign popcount31_4js4_core_202 = input_a[19] & input_a[15];
  assign popcount31_4js4_core_203 = ~(input_a[27] | input_a[27]);
  assign popcount31_4js4_core_204 = input_a[28] ^ input_a[11];
  assign popcount31_4js4_core_205 = ~input_a[16];
  assign popcount31_4js4_core_206 = popcount31_4js4_core_105 & popcount31_4js4_core_190;
  assign popcount31_4js4_core_208 = ~(input_a[12] ^ input_a[20]);
  assign popcount31_4js4_core_210 = popcount31_4js4_core_110 | popcount31_4js4_core_192;
  assign popcount31_4js4_core_211 = popcount31_4js4_core_110 & popcount31_4js4_core_192;
  assign popcount31_4js4_core_212 = input_a[27] & input_a[21];
  assign popcount31_4js4_core_213 = popcount31_4js4_core_210 & popcount31_4js4_core_206;
  assign popcount31_4js4_core_214 = popcount31_4js4_core_211 | popcount31_4js4_core_213;
  assign popcount31_4js4_core_215 = input_a[14] | input_a[15];
  assign popcount31_4js4_core_217 = ~(input_a[4] | input_a[0]);
  assign popcount31_4js4_core_219 = input_a[20] | input_a[28];

  assign popcount31_4js4_out[0] = popcount31_4js4_core_117;
  assign popcount31_4js4_out[1] = popcount31_4js4_core_153;
  assign popcount31_4js4_out[2] = popcount31_4js4_core_117;
  assign popcount31_4js4_out[3] = input_a[25];
  assign popcount31_4js4_out[4] = popcount31_4js4_core_214;
endmodule