// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.47828
// WCE=23.0
// EP=0.936354%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_hs5j(input [29:0] input_a, output [4:0] popcount30_hs5j_out);
  wire popcount30_hs5j_core_033;
  wire popcount30_hs5j_core_034;
  wire popcount30_hs5j_core_035;
  wire popcount30_hs5j_core_036;
  wire popcount30_hs5j_core_040;
  wire popcount30_hs5j_core_041;
  wire popcount30_hs5j_core_042;
  wire popcount30_hs5j_core_044;
  wire popcount30_hs5j_core_046;
  wire popcount30_hs5j_core_047;
  wire popcount30_hs5j_core_049;
  wire popcount30_hs5j_core_051;
  wire popcount30_hs5j_core_053;
  wire popcount30_hs5j_core_055;
  wire popcount30_hs5j_core_056;
  wire popcount30_hs5j_core_057;
  wire popcount30_hs5j_core_059;
  wire popcount30_hs5j_core_063;
  wire popcount30_hs5j_core_064;
  wire popcount30_hs5j_core_066;
  wire popcount30_hs5j_core_068;
  wire popcount30_hs5j_core_069;
  wire popcount30_hs5j_core_070;
  wire popcount30_hs5j_core_071;
  wire popcount30_hs5j_core_072;
  wire popcount30_hs5j_core_073;
  wire popcount30_hs5j_core_075;
  wire popcount30_hs5j_core_077;
  wire popcount30_hs5j_core_079;
  wire popcount30_hs5j_core_080;
  wire popcount30_hs5j_core_082;
  wire popcount30_hs5j_core_083;
  wire popcount30_hs5j_core_084;
  wire popcount30_hs5j_core_085;
  wire popcount30_hs5j_core_086;
  wire popcount30_hs5j_core_087;
  wire popcount30_hs5j_core_088;
  wire popcount30_hs5j_core_089;
  wire popcount30_hs5j_core_090;
  wire popcount30_hs5j_core_091;
  wire popcount30_hs5j_core_093;
  wire popcount30_hs5j_core_095;
  wire popcount30_hs5j_core_097;
  wire popcount30_hs5j_core_102;
  wire popcount30_hs5j_core_103;
  wire popcount30_hs5j_core_104;
  wire popcount30_hs5j_core_105;
  wire popcount30_hs5j_core_107;
  wire popcount30_hs5j_core_112;
  wire popcount30_hs5j_core_113;
  wire popcount30_hs5j_core_115;
  wire popcount30_hs5j_core_116;
  wire popcount30_hs5j_core_117;
  wire popcount30_hs5j_core_118;
  wire popcount30_hs5j_core_120;
  wire popcount30_hs5j_core_121;
  wire popcount30_hs5j_core_122;
  wire popcount30_hs5j_core_123;
  wire popcount30_hs5j_core_125;
  wire popcount30_hs5j_core_126;
  wire popcount30_hs5j_core_127;
  wire popcount30_hs5j_core_129;
  wire popcount30_hs5j_core_130;
  wire popcount30_hs5j_core_131;
  wire popcount30_hs5j_core_135;
  wire popcount30_hs5j_core_137;
  wire popcount30_hs5j_core_138;
  wire popcount30_hs5j_core_139;
  wire popcount30_hs5j_core_141;
  wire popcount30_hs5j_core_142;
  wire popcount30_hs5j_core_143;
  wire popcount30_hs5j_core_146;
  wire popcount30_hs5j_core_150;
  wire popcount30_hs5j_core_151;
  wire popcount30_hs5j_core_152;
  wire popcount30_hs5j_core_153;
  wire popcount30_hs5j_core_154;
  wire popcount30_hs5j_core_156;
  wire popcount30_hs5j_core_157;
  wire popcount30_hs5j_core_158;
  wire popcount30_hs5j_core_161;
  wire popcount30_hs5j_core_163;
  wire popcount30_hs5j_core_164;
  wire popcount30_hs5j_core_165;
  wire popcount30_hs5j_core_166;
  wire popcount30_hs5j_core_168;
  wire popcount30_hs5j_core_169;
  wire popcount30_hs5j_core_173;
  wire popcount30_hs5j_core_175;
  wire popcount30_hs5j_core_177;
  wire popcount30_hs5j_core_178;
  wire popcount30_hs5j_core_181;
  wire popcount30_hs5j_core_182;
  wire popcount30_hs5j_core_183;
  wire popcount30_hs5j_core_184;
  wire popcount30_hs5j_core_185;
  wire popcount30_hs5j_core_186;
  wire popcount30_hs5j_core_187;
  wire popcount30_hs5j_core_188;
  wire popcount30_hs5j_core_193;
  wire popcount30_hs5j_core_195;
  wire popcount30_hs5j_core_197;
  wire popcount30_hs5j_core_198;
  wire popcount30_hs5j_core_199;
  wire popcount30_hs5j_core_200;
  wire popcount30_hs5j_core_201;
  wire popcount30_hs5j_core_202;
  wire popcount30_hs5j_core_205;
  wire popcount30_hs5j_core_207;
  wire popcount30_hs5j_core_213;

  assign popcount30_hs5j_core_033 = input_a[1] & input_a[6];
  assign popcount30_hs5j_core_034 = ~input_a[19];
  assign popcount30_hs5j_core_035 = input_a[20] ^ input_a[28];
  assign popcount30_hs5j_core_036 = input_a[16] & input_a[18];
  assign popcount30_hs5j_core_040 = ~input_a[20];
  assign popcount30_hs5j_core_041 = ~(input_a[17] | input_a[13]);
  assign popcount30_hs5j_core_042 = input_a[10] ^ input_a[26];
  assign popcount30_hs5j_core_044 = input_a[20] & input_a[29];
  assign popcount30_hs5j_core_046 = input_a[24] | input_a[21];
  assign popcount30_hs5j_core_047 = input_a[21] & input_a[2];
  assign popcount30_hs5j_core_049 = input_a[22] | input_a[9];
  assign popcount30_hs5j_core_051 = ~(input_a[6] & input_a[16]);
  assign popcount30_hs5j_core_053 = ~(input_a[6] ^ input_a[25]);
  assign popcount30_hs5j_core_055 = input_a[3] ^ input_a[24];
  assign popcount30_hs5j_core_056 = ~(input_a[23] & input_a[26]);
  assign popcount30_hs5j_core_057 = ~(input_a[10] ^ input_a[25]);
  assign popcount30_hs5j_core_059 = input_a[16] & input_a[29];
  assign popcount30_hs5j_core_063 = ~(input_a[9] & input_a[13]);
  assign popcount30_hs5j_core_064 = input_a[8] ^ input_a[12];
  assign popcount30_hs5j_core_066 = input_a[9] ^ input_a[11];
  assign popcount30_hs5j_core_068 = ~input_a[4];
  assign popcount30_hs5j_core_069 = input_a[21] & input_a[29];
  assign popcount30_hs5j_core_070 = input_a[11] & input_a[7];
  assign popcount30_hs5j_core_071 = input_a[7] ^ input_a[18];
  assign popcount30_hs5j_core_072 = input_a[23] ^ input_a[1];
  assign popcount30_hs5j_core_073 = input_a[17] & input_a[2];
  assign popcount30_hs5j_core_075 = input_a[8] | input_a[28];
  assign popcount30_hs5j_core_077 = ~input_a[21];
  assign popcount30_hs5j_core_079 = input_a[18] | input_a[29];
  assign popcount30_hs5j_core_080 = input_a[11] ^ input_a[27];
  assign popcount30_hs5j_core_082 = ~input_a[17];
  assign popcount30_hs5j_core_083 = ~input_a[1];
  assign popcount30_hs5j_core_084 = ~(input_a[4] & input_a[22]);
  assign popcount30_hs5j_core_085 = ~(input_a[13] | input_a[8]);
  assign popcount30_hs5j_core_086 = input_a[5] ^ input_a[21];
  assign popcount30_hs5j_core_087 = input_a[27] | input_a[28];
  assign popcount30_hs5j_core_088 = ~(input_a[17] & input_a[3]);
  assign popcount30_hs5j_core_089 = ~input_a[29];
  assign popcount30_hs5j_core_090 = input_a[0] | input_a[4];
  assign popcount30_hs5j_core_091 = ~(input_a[10] & input_a[18]);
  assign popcount30_hs5j_core_093 = ~(input_a[24] & input_a[27]);
  assign popcount30_hs5j_core_095 = ~(input_a[7] & input_a[9]);
  assign popcount30_hs5j_core_097 = ~input_a[4];
  assign popcount30_hs5j_core_102 = ~(input_a[13] & input_a[5]);
  assign popcount30_hs5j_core_103 = ~input_a[21];
  assign popcount30_hs5j_core_104 = ~input_a[5];
  assign popcount30_hs5j_core_105 = ~(input_a[7] & input_a[5]);
  assign popcount30_hs5j_core_107 = ~input_a[20];
  assign popcount30_hs5j_core_112 = input_a[8] & input_a[4];
  assign popcount30_hs5j_core_113 = ~(input_a[4] ^ input_a[12]);
  assign popcount30_hs5j_core_115 = ~(input_a[10] & input_a[21]);
  assign popcount30_hs5j_core_116 = ~(input_a[0] | input_a[2]);
  assign popcount30_hs5j_core_117 = input_a[29] | input_a[16];
  assign popcount30_hs5j_core_118 = input_a[23] | input_a[25];
  assign popcount30_hs5j_core_120 = input_a[26] ^ input_a[10];
  assign popcount30_hs5j_core_121 = ~(input_a[1] & input_a[18]);
  assign popcount30_hs5j_core_122 = input_a[16] ^ input_a[13];
  assign popcount30_hs5j_core_123 = ~(input_a[10] ^ input_a[11]);
  assign popcount30_hs5j_core_125 = input_a[1] ^ input_a[13];
  assign popcount30_hs5j_core_126 = input_a[7] ^ input_a[29];
  assign popcount30_hs5j_core_127 = ~(input_a[2] & input_a[2]);
  assign popcount30_hs5j_core_129 = ~(input_a[28] & input_a[4]);
  assign popcount30_hs5j_core_130 = input_a[11] ^ input_a[26];
  assign popcount30_hs5j_core_131 = ~input_a[4];
  assign popcount30_hs5j_core_135 = input_a[10] ^ input_a[11];
  assign popcount30_hs5j_core_137 = ~input_a[14];
  assign popcount30_hs5j_core_138 = ~(input_a[28] & input_a[0]);
  assign popcount30_hs5j_core_139 = input_a[15] | input_a[17];
  assign popcount30_hs5j_core_141 = input_a[17] | input_a[20];
  assign popcount30_hs5j_core_142 = ~(input_a[10] & input_a[0]);
  assign popcount30_hs5j_core_143 = ~(input_a[11] | input_a[26]);
  assign popcount30_hs5j_core_146 = input_a[24] ^ input_a[13];
  assign popcount30_hs5j_core_150 = ~(input_a[24] ^ input_a[12]);
  assign popcount30_hs5j_core_151 = ~(input_a[8] | input_a[11]);
  assign popcount30_hs5j_core_152 = ~input_a[25];
  assign popcount30_hs5j_core_153 = input_a[11] & input_a[22];
  assign popcount30_hs5j_core_154 = ~(input_a[10] | input_a[16]);
  assign popcount30_hs5j_core_156 = ~(input_a[17] | input_a[18]);
  assign popcount30_hs5j_core_157 = ~input_a[9];
  assign popcount30_hs5j_core_158 = input_a[13] & input_a[26];
  assign popcount30_hs5j_core_161 = input_a[13] ^ input_a[23];
  assign popcount30_hs5j_core_163 = input_a[22] | input_a[22];
  assign popcount30_hs5j_core_164 = input_a[27] ^ input_a[10];
  assign popcount30_hs5j_core_165 = ~(input_a[3] | input_a[6]);
  assign popcount30_hs5j_core_166 = ~(input_a[9] & input_a[17]);
  assign popcount30_hs5j_core_168 = ~(input_a[26] & input_a[0]);
  assign popcount30_hs5j_core_169 = ~(input_a[0] | input_a[15]);
  assign popcount30_hs5j_core_173 = ~(input_a[10] & input_a[15]);
  assign popcount30_hs5j_core_175 = input_a[10] ^ input_a[6];
  assign popcount30_hs5j_core_177 = ~(input_a[1] | input_a[25]);
  assign popcount30_hs5j_core_178 = input_a[16] & input_a[25];
  assign popcount30_hs5j_core_181 = ~input_a[7];
  assign popcount30_hs5j_core_182 = ~(input_a[18] | input_a[12]);
  assign popcount30_hs5j_core_183 = input_a[21] ^ input_a[29];
  assign popcount30_hs5j_core_184 = input_a[9] | input_a[16];
  assign popcount30_hs5j_core_185 = ~(input_a[3] | input_a[7]);
  assign popcount30_hs5j_core_186 = ~(input_a[8] & input_a[20]);
  assign popcount30_hs5j_core_187 = ~input_a[1];
  assign popcount30_hs5j_core_188 = ~(input_a[6] | input_a[6]);
  assign popcount30_hs5j_core_193 = ~input_a[13];
  assign popcount30_hs5j_core_195 = input_a[13] | input_a[13];
  assign popcount30_hs5j_core_197 = ~(input_a[9] & input_a[25]);
  assign popcount30_hs5j_core_198 = ~input_a[7];
  assign popcount30_hs5j_core_199 = ~(input_a[12] & input_a[1]);
  assign popcount30_hs5j_core_200 = ~input_a[13];
  assign popcount30_hs5j_core_201 = input_a[0] ^ input_a[10];
  assign popcount30_hs5j_core_202 = ~(input_a[21] & input_a[3]);
  assign popcount30_hs5j_core_205 = input_a[0] | input_a[7];
  assign popcount30_hs5j_core_207 = input_a[14] ^ input_a[1];
  assign popcount30_hs5j_core_213 = ~(input_a[7] & input_a[0]);

  assign popcount30_hs5j_out[0] = 1'b0;
  assign popcount30_hs5j_out[1] = 1'b0;
  assign popcount30_hs5j_out[2] = 1'b0;
  assign popcount30_hs5j_out[3] = input_a[23];
  assign popcount30_hs5j_out[4] = 1'b1;
endmodule