// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.62886
// WCE=28.0
// EP=0.966115%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_h738(input [20:0] input_a, output [4:0] popcount21_h738_out);
  wire popcount21_h738_core_023;
  wire popcount21_h738_core_024;
  wire popcount21_h738_core_025;
  wire popcount21_h738_core_026;
  wire popcount21_h738_core_027;
  wire popcount21_h738_core_028;
  wire popcount21_h738_core_029;
  wire popcount21_h738_core_030;
  wire popcount21_h738_core_031;
  wire popcount21_h738_core_033;
  wire popcount21_h738_core_034;
  wire popcount21_h738_core_035;
  wire popcount21_h738_core_036;
  wire popcount21_h738_core_039;
  wire popcount21_h738_core_040;
  wire popcount21_h738_core_044;
  wire popcount21_h738_core_045;
  wire popcount21_h738_core_046;
  wire popcount21_h738_core_049;
  wire popcount21_h738_core_050;
  wire popcount21_h738_core_051;
  wire popcount21_h738_core_052;
  wire popcount21_h738_core_053;
  wire popcount21_h738_core_054;
  wire popcount21_h738_core_055_not;
  wire popcount21_h738_core_056;
  wire popcount21_h738_core_057;
  wire popcount21_h738_core_058;
  wire popcount21_h738_core_061;
  wire popcount21_h738_core_063;
  wire popcount21_h738_core_064;
  wire popcount21_h738_core_065;
  wire popcount21_h738_core_066;
  wire popcount21_h738_core_069;
  wire popcount21_h738_core_071;
  wire popcount21_h738_core_073;
  wire popcount21_h738_core_075;
  wire popcount21_h738_core_076;
  wire popcount21_h738_core_077;
  wire popcount21_h738_core_078;
  wire popcount21_h738_core_080;
  wire popcount21_h738_core_082;
  wire popcount21_h738_core_083;
  wire popcount21_h738_core_084;
  wire popcount21_h738_core_085;
  wire popcount21_h738_core_087;
  wire popcount21_h738_core_088;
  wire popcount21_h738_core_089;
  wire popcount21_h738_core_090_not;
  wire popcount21_h738_core_091;
  wire popcount21_h738_core_092;
  wire popcount21_h738_core_093;
  wire popcount21_h738_core_094;
  wire popcount21_h738_core_096;
  wire popcount21_h738_core_097;
  wire popcount21_h738_core_099;
  wire popcount21_h738_core_100;
  wire popcount21_h738_core_101;
  wire popcount21_h738_core_102;
  wire popcount21_h738_core_103;
  wire popcount21_h738_core_104;
  wire popcount21_h738_core_105;
  wire popcount21_h738_core_106;
  wire popcount21_h738_core_107;
  wire popcount21_h738_core_108;
  wire popcount21_h738_core_109;
  wire popcount21_h738_core_110;
  wire popcount21_h738_core_113;
  wire popcount21_h738_core_114;
  wire popcount21_h738_core_115;
  wire popcount21_h738_core_117;
  wire popcount21_h738_core_118_not;
  wire popcount21_h738_core_120;
  wire popcount21_h738_core_123;
  wire popcount21_h738_core_126;
  wire popcount21_h738_core_127;
  wire popcount21_h738_core_130;
  wire popcount21_h738_core_131;
  wire popcount21_h738_core_132;
  wire popcount21_h738_core_133;
  wire popcount21_h738_core_136;
  wire popcount21_h738_core_139;
  wire popcount21_h738_core_141;
  wire popcount21_h738_core_143;
  wire popcount21_h738_core_144;
  wire popcount21_h738_core_145;
  wire popcount21_h738_core_146;
  wire popcount21_h738_core_148;
  wire popcount21_h738_core_150;
  wire popcount21_h738_core_151;

  assign popcount21_h738_core_023 = input_a[17] & input_a[12];
  assign popcount21_h738_core_024 = ~(input_a[12] ^ input_a[20]);
  assign popcount21_h738_core_025 = input_a[18] | input_a[20];
  assign popcount21_h738_core_026 = input_a[8] & input_a[20];
  assign popcount21_h738_core_027 = ~(input_a[0] & input_a[11]);
  assign popcount21_h738_core_028 = ~(input_a[6] | input_a[1]);
  assign popcount21_h738_core_029 = input_a[16] ^ input_a[0];
  assign popcount21_h738_core_030 = ~(input_a[12] & input_a[17]);
  assign popcount21_h738_core_031 = ~input_a[11];
  assign popcount21_h738_core_033 = ~input_a[13];
  assign popcount21_h738_core_034 = ~(input_a[5] & input_a[7]);
  assign popcount21_h738_core_035 = ~(input_a[2] & input_a[8]);
  assign popcount21_h738_core_036 = ~input_a[2];
  assign popcount21_h738_core_039 = ~input_a[18];
  assign popcount21_h738_core_040 = ~(input_a[18] ^ input_a[18]);
  assign popcount21_h738_core_044 = ~input_a[20];
  assign popcount21_h738_core_045 = input_a[3] | input_a[7];
  assign popcount21_h738_core_046 = ~(input_a[1] ^ input_a[3]);
  assign popcount21_h738_core_049 = input_a[18] | input_a[18];
  assign popcount21_h738_core_050 = input_a[17] | input_a[20];
  assign popcount21_h738_core_051 = ~(input_a[18] | input_a[13]);
  assign popcount21_h738_core_052 = input_a[10] ^ input_a[18];
  assign popcount21_h738_core_053 = ~(input_a[6] ^ input_a[11]);
  assign popcount21_h738_core_054 = ~input_a[10];
  assign popcount21_h738_core_055_not = ~input_a[6];
  assign popcount21_h738_core_056 = input_a[8] ^ input_a[2];
  assign popcount21_h738_core_057 = input_a[4] | input_a[7];
  assign popcount21_h738_core_058 = ~(input_a[7] & input_a[18]);
  assign popcount21_h738_core_061 = ~(input_a[4] | input_a[13]);
  assign popcount21_h738_core_063 = ~(input_a[3] | input_a[8]);
  assign popcount21_h738_core_064 = input_a[19] | input_a[16];
  assign popcount21_h738_core_065 = ~input_a[7];
  assign popcount21_h738_core_066 = input_a[17] ^ input_a[7];
  assign popcount21_h738_core_069 = ~(input_a[7] | input_a[17]);
  assign popcount21_h738_core_071 = input_a[1] ^ input_a[17];
  assign popcount21_h738_core_073 = input_a[4] | input_a[7];
  assign popcount21_h738_core_075 = ~input_a[0];
  assign popcount21_h738_core_076 = input_a[3] ^ input_a[8];
  assign popcount21_h738_core_077 = input_a[19] | input_a[19];
  assign popcount21_h738_core_078 = input_a[19] ^ input_a[12];
  assign popcount21_h738_core_080 = ~input_a[5];
  assign popcount21_h738_core_082 = ~(input_a[18] | input_a[2]);
  assign popcount21_h738_core_083 = ~(input_a[10] | input_a[1]);
  assign popcount21_h738_core_084 = ~(input_a[10] ^ input_a[9]);
  assign popcount21_h738_core_085 = ~(input_a[17] & input_a[2]);
  assign popcount21_h738_core_087 = input_a[17] & input_a[0];
  assign popcount21_h738_core_088 = ~input_a[1];
  assign popcount21_h738_core_089 = ~(input_a[6] & input_a[9]);
  assign popcount21_h738_core_090_not = ~input_a[11];
  assign popcount21_h738_core_091 = ~input_a[9];
  assign popcount21_h738_core_092 = ~input_a[16];
  assign popcount21_h738_core_093 = ~(input_a[5] | input_a[17]);
  assign popcount21_h738_core_094 = ~(input_a[17] & input_a[1]);
  assign popcount21_h738_core_096 = ~(input_a[10] ^ input_a[12]);
  assign popcount21_h738_core_097 = ~(input_a[19] & input_a[6]);
  assign popcount21_h738_core_099 = ~input_a[15];
  assign popcount21_h738_core_100 = ~(input_a[15] & input_a[10]);
  assign popcount21_h738_core_101 = ~(input_a[17] & input_a[13]);
  assign popcount21_h738_core_102 = input_a[15] | input_a[16];
  assign popcount21_h738_core_103 = input_a[20] & input_a[8];
  assign popcount21_h738_core_104 = input_a[19] & input_a[7];
  assign popcount21_h738_core_105 = input_a[2] | input_a[1];
  assign popcount21_h738_core_106 = ~input_a[7];
  assign popcount21_h738_core_107 = ~input_a[13];
  assign popcount21_h738_core_108 = input_a[9] ^ input_a[16];
  assign popcount21_h738_core_109 = input_a[4] | input_a[9];
  assign popcount21_h738_core_110 = input_a[3] ^ input_a[4];
  assign popcount21_h738_core_113 = input_a[12] ^ input_a[1];
  assign popcount21_h738_core_114 = ~(input_a[16] & input_a[14]);
  assign popcount21_h738_core_115 = ~(input_a[2] | input_a[13]);
  assign popcount21_h738_core_117 = input_a[12] ^ input_a[13];
  assign popcount21_h738_core_118_not = ~input_a[13];
  assign popcount21_h738_core_120 = ~(input_a[18] | input_a[17]);
  assign popcount21_h738_core_123 = ~(input_a[18] & input_a[16]);
  assign popcount21_h738_core_126 = ~(input_a[11] ^ input_a[17]);
  assign popcount21_h738_core_127 = ~input_a[11];
  assign popcount21_h738_core_130 = ~(input_a[11] | input_a[13]);
  assign popcount21_h738_core_131 = ~(input_a[6] ^ input_a[6]);
  assign popcount21_h738_core_132 = ~input_a[20];
  assign popcount21_h738_core_133 = ~input_a[1];
  assign popcount21_h738_core_136 = ~input_a[16];
  assign popcount21_h738_core_139 = ~(input_a[15] | input_a[19]);
  assign popcount21_h738_core_141 = ~(input_a[20] & input_a[6]);
  assign popcount21_h738_core_143 = input_a[6] ^ input_a[14];
  assign popcount21_h738_core_144 = ~input_a[9];
  assign popcount21_h738_core_145 = input_a[11] | input_a[11];
  assign popcount21_h738_core_146 = ~(input_a[19] ^ input_a[10]);
  assign popcount21_h738_core_148 = ~(input_a[4] | input_a[18]);
  assign popcount21_h738_core_150 = input_a[19] | input_a[8];
  assign popcount21_h738_core_151 = ~input_a[13];

  assign popcount21_h738_out[0] = 1'b1;
  assign popcount21_h738_out[1] = input_a[6];
  assign popcount21_h738_out[2] = input_a[6];
  assign popcount21_h738_out[3] = input_a[13];
  assign popcount21_h738_out[4] = input_a[15];
endmodule