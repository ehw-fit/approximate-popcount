// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=0.0
// WCE=0.0
// EP=0.0%
// Printed PDK parameters:
//  Area=58065925.0
//  Delay=68229544.0
//  Power=3011000.0

module popcount18_ldz5(input [17:0] input_a, output [4:0] popcount18_ldz5_out);
  wire popcount18_ldz5_core_020;
  wire popcount18_ldz5_core_021;
  wire popcount18_ldz5_core_022;
  wire popcount18_ldz5_core_023;
  wire popcount18_ldz5_core_024;
  wire popcount18_ldz5_core_025;
  wire popcount18_ldz5_core_026;
  wire popcount18_ldz5_core_027;
  wire popcount18_ldz5_core_028;
  wire popcount18_ldz5_core_031;
  wire popcount18_ldz5_core_032;
  wire popcount18_ldz5_core_033;
  wire popcount18_ldz5_core_034;
  wire popcount18_ldz5_core_035;
  wire popcount18_ldz5_core_036;
  wire popcount18_ldz5_core_037;
  wire popcount18_ldz5_core_039;
  wire popcount18_ldz5_core_040;
  wire popcount18_ldz5_core_041;
  wire popcount18_ldz5_core_042;
  wire popcount18_ldz5_core_043;
  wire popcount18_ldz5_core_044;
  wire popcount18_ldz5_core_045;
  wire popcount18_ldz5_core_048;
  wire popcount18_ldz5_core_049;
  wire popcount18_ldz5_core_050;
  wire popcount18_ldz5_core_051;
  wire popcount18_ldz5_core_052;
  wire popcount18_ldz5_core_053;
  wire popcount18_ldz5_core_054;
  wire popcount18_ldz5_core_055;
  wire popcount18_ldz5_core_056;
  wire popcount18_ldz5_core_057;
  wire popcount18_ldz5_core_058;
  wire popcount18_ldz5_core_059;
  wire popcount18_ldz5_core_062;
  wire popcount18_ldz5_core_063;
  wire popcount18_ldz5_core_064;
  wire popcount18_ldz5_core_065;
  wire popcount18_ldz5_core_066;
  wire popcount18_ldz5_core_067;
  wire popcount18_ldz5_core_068;
  wire popcount18_ldz5_core_069;
  wire popcount18_ldz5_core_070;
  wire popcount18_ldz5_core_073;
  wire popcount18_ldz5_core_074;
  wire popcount18_ldz5_core_075;
  wire popcount18_ldz5_core_076;
  wire popcount18_ldz5_core_077;
  wire popcount18_ldz5_core_078;
  wire popcount18_ldz5_core_079;
  wire popcount18_ldz5_core_081;
  wire popcount18_ldz5_core_082;
  wire popcount18_ldz5_core_083;
  wire popcount18_ldz5_core_084;
  wire popcount18_ldz5_core_085;
  wire popcount18_ldz5_core_086;
  wire popcount18_ldz5_core_087;
  wire popcount18_ldz5_core_090;
  wire popcount18_ldz5_core_091;
  wire popcount18_ldz5_core_092;
  wire popcount18_ldz5_core_093;
  wire popcount18_ldz5_core_094;
  wire popcount18_ldz5_core_095;
  wire popcount18_ldz5_core_096;
  wire popcount18_ldz5_core_097;
  wire popcount18_ldz5_core_098;
  wire popcount18_ldz5_core_099;
  wire popcount18_ldz5_core_100;
  wire popcount18_ldz5_core_101;
  wire popcount18_ldz5_core_103;
  wire popcount18_ldz5_core_104;
  wire popcount18_ldz5_core_105;
  wire popcount18_ldz5_core_106;
  wire popcount18_ldz5_core_107;
  wire popcount18_ldz5_core_108;
  wire popcount18_ldz5_core_109;
  wire popcount18_ldz5_core_110;
  wire popcount18_ldz5_core_111;
  wire popcount18_ldz5_core_112;
  wire popcount18_ldz5_core_113;
  wire popcount18_ldz5_core_114;
  wire popcount18_ldz5_core_115;
  wire popcount18_ldz5_core_116;
  wire popcount18_ldz5_core_117;
  wire popcount18_ldz5_core_118;
  wire popcount18_ldz5_core_119;
  wire popcount18_ldz5_core_120;
  wire popcount18_ldz5_core_123;
  wire popcount18_ldz5_core_124;

  assign popcount18_ldz5_core_020 = input_a[0] ^ input_a[1];
  assign popcount18_ldz5_core_021 = input_a[0] & input_a[1];
  assign popcount18_ldz5_core_022 = input_a[2] ^ input_a[3];
  assign popcount18_ldz5_core_023 = input_a[2] & input_a[3];
  assign popcount18_ldz5_core_024 = popcount18_ldz5_core_020 ^ popcount18_ldz5_core_022;
  assign popcount18_ldz5_core_025 = popcount18_ldz5_core_020 & popcount18_ldz5_core_022;
  assign popcount18_ldz5_core_026 = popcount18_ldz5_core_021 ^ popcount18_ldz5_core_023;
  assign popcount18_ldz5_core_027 = popcount18_ldz5_core_021 & popcount18_ldz5_core_023;
  assign popcount18_ldz5_core_028 = popcount18_ldz5_core_026 | popcount18_ldz5_core_025;
  assign popcount18_ldz5_core_031 = input_a[4] ^ input_a[5];
  assign popcount18_ldz5_core_032 = input_a[4] & input_a[5];
  assign popcount18_ldz5_core_033 = input_a[7] ^ input_a[8];
  assign popcount18_ldz5_core_034 = input_a[7] & input_a[8];
  assign popcount18_ldz5_core_035 = input_a[6] ^ popcount18_ldz5_core_033;
  assign popcount18_ldz5_core_036 = input_a[6] & popcount18_ldz5_core_033;
  assign popcount18_ldz5_core_037 = popcount18_ldz5_core_034 | popcount18_ldz5_core_036;
  assign popcount18_ldz5_core_039 = popcount18_ldz5_core_031 ^ popcount18_ldz5_core_035;
  assign popcount18_ldz5_core_040 = popcount18_ldz5_core_031 & popcount18_ldz5_core_035;
  assign popcount18_ldz5_core_041 = popcount18_ldz5_core_032 ^ popcount18_ldz5_core_037;
  assign popcount18_ldz5_core_042 = popcount18_ldz5_core_032 & popcount18_ldz5_core_037;
  assign popcount18_ldz5_core_043 = popcount18_ldz5_core_041 ^ popcount18_ldz5_core_040;
  assign popcount18_ldz5_core_044 = popcount18_ldz5_core_041 & popcount18_ldz5_core_040;
  assign popcount18_ldz5_core_045 = popcount18_ldz5_core_042 | popcount18_ldz5_core_044;
  assign popcount18_ldz5_core_048 = popcount18_ldz5_core_024 ^ popcount18_ldz5_core_039;
  assign popcount18_ldz5_core_049 = popcount18_ldz5_core_024 & popcount18_ldz5_core_039;
  assign popcount18_ldz5_core_050 = popcount18_ldz5_core_028 ^ popcount18_ldz5_core_043;
  assign popcount18_ldz5_core_051 = popcount18_ldz5_core_028 & popcount18_ldz5_core_043;
  assign popcount18_ldz5_core_052 = popcount18_ldz5_core_050 ^ popcount18_ldz5_core_049;
  assign popcount18_ldz5_core_053 = popcount18_ldz5_core_050 & popcount18_ldz5_core_049;
  assign popcount18_ldz5_core_054 = popcount18_ldz5_core_051 | popcount18_ldz5_core_053;
  assign popcount18_ldz5_core_055 = popcount18_ldz5_core_027 ^ popcount18_ldz5_core_045;
  assign popcount18_ldz5_core_056 = popcount18_ldz5_core_027 & popcount18_ldz5_core_045;
  assign popcount18_ldz5_core_057 = popcount18_ldz5_core_055 ^ popcount18_ldz5_core_054;
  assign popcount18_ldz5_core_058 = popcount18_ldz5_core_055 & popcount18_ldz5_core_054;
  assign popcount18_ldz5_core_059 = popcount18_ldz5_core_056 | popcount18_ldz5_core_058;
  assign popcount18_ldz5_core_062 = input_a[9] ^ input_a[10];
  assign popcount18_ldz5_core_063 = input_a[9] & input_a[10];
  assign popcount18_ldz5_core_064 = input_a[11] ^ input_a[12];
  assign popcount18_ldz5_core_065 = input_a[11] & input_a[12];
  assign popcount18_ldz5_core_066 = popcount18_ldz5_core_062 ^ popcount18_ldz5_core_064;
  assign popcount18_ldz5_core_067 = popcount18_ldz5_core_062 & popcount18_ldz5_core_064;
  assign popcount18_ldz5_core_068 = popcount18_ldz5_core_063 ^ popcount18_ldz5_core_065;
  assign popcount18_ldz5_core_069 = popcount18_ldz5_core_063 & popcount18_ldz5_core_065;
  assign popcount18_ldz5_core_070 = popcount18_ldz5_core_068 | popcount18_ldz5_core_067;
  assign popcount18_ldz5_core_073 = input_a[13] ^ input_a[14];
  assign popcount18_ldz5_core_074 = input_a[13] & input_a[14];
  assign popcount18_ldz5_core_075 = input_a[16] ^ input_a[17];
  assign popcount18_ldz5_core_076 = input_a[16] & input_a[17];
  assign popcount18_ldz5_core_077 = input_a[15] ^ popcount18_ldz5_core_075;
  assign popcount18_ldz5_core_078 = input_a[15] & popcount18_ldz5_core_075;
  assign popcount18_ldz5_core_079 = popcount18_ldz5_core_076 | popcount18_ldz5_core_078;
  assign popcount18_ldz5_core_081 = popcount18_ldz5_core_073 ^ popcount18_ldz5_core_077;
  assign popcount18_ldz5_core_082 = popcount18_ldz5_core_073 & popcount18_ldz5_core_077;
  assign popcount18_ldz5_core_083 = popcount18_ldz5_core_074 ^ popcount18_ldz5_core_079;
  assign popcount18_ldz5_core_084 = popcount18_ldz5_core_074 & popcount18_ldz5_core_079;
  assign popcount18_ldz5_core_085 = popcount18_ldz5_core_083 ^ popcount18_ldz5_core_082;
  assign popcount18_ldz5_core_086 = popcount18_ldz5_core_083 & popcount18_ldz5_core_082;
  assign popcount18_ldz5_core_087 = popcount18_ldz5_core_084 | popcount18_ldz5_core_086;
  assign popcount18_ldz5_core_090 = popcount18_ldz5_core_066 ^ popcount18_ldz5_core_081;
  assign popcount18_ldz5_core_091 = popcount18_ldz5_core_066 & popcount18_ldz5_core_081;
  assign popcount18_ldz5_core_092 = popcount18_ldz5_core_070 ^ popcount18_ldz5_core_085;
  assign popcount18_ldz5_core_093 = popcount18_ldz5_core_070 & popcount18_ldz5_core_085;
  assign popcount18_ldz5_core_094 = popcount18_ldz5_core_092 ^ popcount18_ldz5_core_091;
  assign popcount18_ldz5_core_095 = popcount18_ldz5_core_092 & popcount18_ldz5_core_091;
  assign popcount18_ldz5_core_096 = popcount18_ldz5_core_093 | popcount18_ldz5_core_095;
  assign popcount18_ldz5_core_097 = popcount18_ldz5_core_069 ^ popcount18_ldz5_core_087;
  assign popcount18_ldz5_core_098 = popcount18_ldz5_core_069 & popcount18_ldz5_core_087;
  assign popcount18_ldz5_core_099 = popcount18_ldz5_core_097 ^ popcount18_ldz5_core_096;
  assign popcount18_ldz5_core_100 = popcount18_ldz5_core_097 & popcount18_ldz5_core_096;
  assign popcount18_ldz5_core_101 = popcount18_ldz5_core_098 | popcount18_ldz5_core_100;
  assign popcount18_ldz5_core_103 = input_a[15] | input_a[7];
  assign popcount18_ldz5_core_104 = popcount18_ldz5_core_048 ^ popcount18_ldz5_core_090;
  assign popcount18_ldz5_core_105 = popcount18_ldz5_core_048 & popcount18_ldz5_core_090;
  assign popcount18_ldz5_core_106 = popcount18_ldz5_core_052 ^ popcount18_ldz5_core_094;
  assign popcount18_ldz5_core_107 = popcount18_ldz5_core_052 & popcount18_ldz5_core_094;
  assign popcount18_ldz5_core_108 = popcount18_ldz5_core_106 ^ popcount18_ldz5_core_105;
  assign popcount18_ldz5_core_109 = popcount18_ldz5_core_106 & popcount18_ldz5_core_105;
  assign popcount18_ldz5_core_110 = popcount18_ldz5_core_107 | popcount18_ldz5_core_109;
  assign popcount18_ldz5_core_111 = popcount18_ldz5_core_057 ^ popcount18_ldz5_core_099;
  assign popcount18_ldz5_core_112 = popcount18_ldz5_core_057 & popcount18_ldz5_core_099;
  assign popcount18_ldz5_core_113 = popcount18_ldz5_core_111 ^ popcount18_ldz5_core_110;
  assign popcount18_ldz5_core_114 = popcount18_ldz5_core_111 & popcount18_ldz5_core_110;
  assign popcount18_ldz5_core_115 = popcount18_ldz5_core_112 | popcount18_ldz5_core_114;
  assign popcount18_ldz5_core_116 = popcount18_ldz5_core_059 ^ popcount18_ldz5_core_101;
  assign popcount18_ldz5_core_117 = popcount18_ldz5_core_059 & popcount18_ldz5_core_101;
  assign popcount18_ldz5_core_118 = popcount18_ldz5_core_116 ^ popcount18_ldz5_core_115;
  assign popcount18_ldz5_core_119 = popcount18_ldz5_core_116 & popcount18_ldz5_core_115;
  assign popcount18_ldz5_core_120 = popcount18_ldz5_core_117 | popcount18_ldz5_core_119;
  assign popcount18_ldz5_core_123 = ~input_a[14];
  assign popcount18_ldz5_core_124 = ~(input_a[10] ^ input_a[7]);

  assign popcount18_ldz5_out[0] = popcount18_ldz5_core_104;
  assign popcount18_ldz5_out[1] = popcount18_ldz5_core_108;
  assign popcount18_ldz5_out[2] = popcount18_ldz5_core_113;
  assign popcount18_ldz5_out[3] = popcount18_ldz5_core_118;
  assign popcount18_ldz5_out[4] = popcount18_ldz5_core_120;
endmodule