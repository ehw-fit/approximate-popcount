// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.93124
// WCE=21.0
// EP=0.930097%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_en6z(input [32:0] input_a, output [5:0] popcount33_en6z_out);
  wire popcount33_en6z_core_036;
  wire popcount33_en6z_core_037;
  wire popcount33_en6z_core_038;
  wire popcount33_en6z_core_040;
  wire popcount33_en6z_core_041;
  wire popcount33_en6z_core_042;
  wire popcount33_en6z_core_043_not;
  wire popcount33_en6z_core_045;
  wire popcount33_en6z_core_047;
  wire popcount33_en6z_core_048;
  wire popcount33_en6z_core_049;
  wire popcount33_en6z_core_051;
  wire popcount33_en6z_core_052;
  wire popcount33_en6z_core_055;
  wire popcount33_en6z_core_056;
  wire popcount33_en6z_core_057;
  wire popcount33_en6z_core_059;
  wire popcount33_en6z_core_060;
  wire popcount33_en6z_core_061;
  wire popcount33_en6z_core_062;
  wire popcount33_en6z_core_063;
  wire popcount33_en6z_core_065;
  wire popcount33_en6z_core_067;
  wire popcount33_en6z_core_072;
  wire popcount33_en6z_core_073;
  wire popcount33_en6z_core_075;
  wire popcount33_en6z_core_080;
  wire popcount33_en6z_core_082;
  wire popcount33_en6z_core_086;
  wire popcount33_en6z_core_087;
  wire popcount33_en6z_core_088;
  wire popcount33_en6z_core_089;
  wire popcount33_en6z_core_090;
  wire popcount33_en6z_core_091;
  wire popcount33_en6z_core_092;
  wire popcount33_en6z_core_093;
  wire popcount33_en6z_core_095;
  wire popcount33_en6z_core_097;
  wire popcount33_en6z_core_101;
  wire popcount33_en6z_core_104;
  wire popcount33_en6z_core_107;
  wire popcount33_en6z_core_110;
  wire popcount33_en6z_core_111;
  wire popcount33_en6z_core_112;
  wire popcount33_en6z_core_113;
  wire popcount33_en6z_core_114;
  wire popcount33_en6z_core_117;
  wire popcount33_en6z_core_119;
  wire popcount33_en6z_core_121;
  wire popcount33_en6z_core_122;
  wire popcount33_en6z_core_124;
  wire popcount33_en6z_core_125;
  wire popcount33_en6z_core_126;
  wire popcount33_en6z_core_127;
  wire popcount33_en6z_core_128;
  wire popcount33_en6z_core_129;
  wire popcount33_en6z_core_131;
  wire popcount33_en6z_core_133;
  wire popcount33_en6z_core_135;
  wire popcount33_en6z_core_136;
  wire popcount33_en6z_core_137;
  wire popcount33_en6z_core_138;
  wire popcount33_en6z_core_139;
  wire popcount33_en6z_core_140;
  wire popcount33_en6z_core_141;
  wire popcount33_en6z_core_142;
  wire popcount33_en6z_core_143;
  wire popcount33_en6z_core_146;
  wire popcount33_en6z_core_147;
  wire popcount33_en6z_core_148;
  wire popcount33_en6z_core_150;
  wire popcount33_en6z_core_152;
  wire popcount33_en6z_core_154;
  wire popcount33_en6z_core_156;
  wire popcount33_en6z_core_157;
  wire popcount33_en6z_core_158;
  wire popcount33_en6z_core_160;
  wire popcount33_en6z_core_162;
  wire popcount33_en6z_core_163;
  wire popcount33_en6z_core_164;
  wire popcount33_en6z_core_166;
  wire popcount33_en6z_core_167;
  wire popcount33_en6z_core_168;
  wire popcount33_en6z_core_170;
  wire popcount33_en6z_core_173;
  wire popcount33_en6z_core_176;
  wire popcount33_en6z_core_180;
  wire popcount33_en6z_core_182;
  wire popcount33_en6z_core_183;
  wire popcount33_en6z_core_186;
  wire popcount33_en6z_core_187;
  wire popcount33_en6z_core_188;
  wire popcount33_en6z_core_189;
  wire popcount33_en6z_core_193;
  wire popcount33_en6z_core_194;
  wire popcount33_en6z_core_195;
  wire popcount33_en6z_core_196;
  wire popcount33_en6z_core_197;
  wire popcount33_en6z_core_198;
  wire popcount33_en6z_core_199;
  wire popcount33_en6z_core_200_not;
  wire popcount33_en6z_core_203;
  wire popcount33_en6z_core_204;
  wire popcount33_en6z_core_205;
  wire popcount33_en6z_core_206;
  wire popcount33_en6z_core_207;
  wire popcount33_en6z_core_209;
  wire popcount33_en6z_core_210;
  wire popcount33_en6z_core_212;
  wire popcount33_en6z_core_213;
  wire popcount33_en6z_core_214;
  wire popcount33_en6z_core_215;
  wire popcount33_en6z_core_218;
  wire popcount33_en6z_core_219;
  wire popcount33_en6z_core_221;
  wire popcount33_en6z_core_222;
  wire popcount33_en6z_core_223;
  wire popcount33_en6z_core_224;
  wire popcount33_en6z_core_225;
  wire popcount33_en6z_core_226_not;
  wire popcount33_en6z_core_228;
  wire popcount33_en6z_core_229;
  wire popcount33_en6z_core_230;
  wire popcount33_en6z_core_231;
  wire popcount33_en6z_core_233;
  wire popcount33_en6z_core_234;
  wire popcount33_en6z_core_237;

  assign popcount33_en6z_core_036 = input_a[17] | input_a[5];
  assign popcount33_en6z_core_037 = ~(input_a[25] & input_a[30]);
  assign popcount33_en6z_core_038 = ~input_a[3];
  assign popcount33_en6z_core_040 = input_a[2] & input_a[17];
  assign popcount33_en6z_core_041 = ~(input_a[23] ^ input_a[12]);
  assign popcount33_en6z_core_042 = input_a[0] & input_a[32];
  assign popcount33_en6z_core_043_not = ~input_a[8];
  assign popcount33_en6z_core_045 = ~input_a[4];
  assign popcount33_en6z_core_047 = ~input_a[25];
  assign popcount33_en6z_core_048 = input_a[15] | input_a[0];
  assign popcount33_en6z_core_049 = ~(input_a[28] & input_a[1]);
  assign popcount33_en6z_core_051 = ~input_a[2];
  assign popcount33_en6z_core_052 = input_a[2] & input_a[17];
  assign popcount33_en6z_core_055 = input_a[14] & input_a[18];
  assign popcount33_en6z_core_056 = ~input_a[30];
  assign popcount33_en6z_core_057 = ~input_a[12];
  assign popcount33_en6z_core_059 = input_a[18] & input_a[9];
  assign popcount33_en6z_core_060 = input_a[14] | input_a[31];
  assign popcount33_en6z_core_061 = ~(input_a[15] ^ input_a[7]);
  assign popcount33_en6z_core_062 = ~(input_a[7] & input_a[0]);
  assign popcount33_en6z_core_063 = ~input_a[26];
  assign popcount33_en6z_core_065 = ~(input_a[9] | input_a[22]);
  assign popcount33_en6z_core_067 = ~(input_a[27] & input_a[32]);
  assign popcount33_en6z_core_072 = input_a[13] & input_a[0];
  assign popcount33_en6z_core_073 = ~(input_a[21] & input_a[20]);
  assign popcount33_en6z_core_075 = ~input_a[27];
  assign popcount33_en6z_core_080 = ~(input_a[10] ^ input_a[18]);
  assign popcount33_en6z_core_082 = ~(input_a[27] & input_a[20]);
  assign popcount33_en6z_core_086 = ~input_a[3];
  assign popcount33_en6z_core_087 = ~(input_a[6] & input_a[19]);
  assign popcount33_en6z_core_088 = ~(input_a[32] & input_a[0]);
  assign popcount33_en6z_core_089 = ~(input_a[16] & input_a[5]);
  assign popcount33_en6z_core_090 = input_a[4] | input_a[9];
  assign popcount33_en6z_core_091 = ~(input_a[22] ^ input_a[23]);
  assign popcount33_en6z_core_092 = ~(input_a[6] | input_a[14]);
  assign popcount33_en6z_core_093 = input_a[8] ^ input_a[8];
  assign popcount33_en6z_core_095 = input_a[17] ^ input_a[6];
  assign popcount33_en6z_core_097 = input_a[12] ^ input_a[14];
  assign popcount33_en6z_core_101 = ~(input_a[24] | input_a[18]);
  assign popcount33_en6z_core_104 = ~(input_a[5] ^ input_a[13]);
  assign popcount33_en6z_core_107 = input_a[24] | input_a[22];
  assign popcount33_en6z_core_110 = ~input_a[14];
  assign popcount33_en6z_core_111 = input_a[3] | input_a[13];
  assign popcount33_en6z_core_112 = ~(input_a[14] | input_a[8]);
  assign popcount33_en6z_core_113 = input_a[20] ^ input_a[22];
  assign popcount33_en6z_core_114 = ~input_a[26];
  assign popcount33_en6z_core_117 = input_a[31] ^ input_a[1];
  assign popcount33_en6z_core_119 = ~(input_a[29] | input_a[6]);
  assign popcount33_en6z_core_121 = ~input_a[5];
  assign popcount33_en6z_core_122 = ~(input_a[2] ^ input_a[13]);
  assign popcount33_en6z_core_124 = ~(input_a[9] ^ input_a[25]);
  assign popcount33_en6z_core_125 = input_a[7] | input_a[23];
  assign popcount33_en6z_core_126 = input_a[0] ^ input_a[15];
  assign popcount33_en6z_core_127 = input_a[15] ^ input_a[32];
  assign popcount33_en6z_core_128 = ~input_a[5];
  assign popcount33_en6z_core_129 = ~(input_a[9] ^ input_a[29]);
  assign popcount33_en6z_core_131 = input_a[3] ^ input_a[21];
  assign popcount33_en6z_core_133 = ~(input_a[10] | input_a[5]);
  assign popcount33_en6z_core_135 = ~(input_a[9] ^ input_a[26]);
  assign popcount33_en6z_core_136 = input_a[23] ^ input_a[27];
  assign popcount33_en6z_core_137 = input_a[6] & input_a[1];
  assign popcount33_en6z_core_138 = ~(input_a[5] ^ input_a[2]);
  assign popcount33_en6z_core_139 = input_a[16] | input_a[9];
  assign popcount33_en6z_core_140 = ~(input_a[32] & input_a[28]);
  assign popcount33_en6z_core_141 = input_a[13] | input_a[25];
  assign popcount33_en6z_core_142 = ~input_a[28];
  assign popcount33_en6z_core_143 = ~input_a[16];
  assign popcount33_en6z_core_146 = input_a[3] & input_a[9];
  assign popcount33_en6z_core_147 = ~(input_a[22] | input_a[3]);
  assign popcount33_en6z_core_148 = ~(input_a[12] ^ input_a[18]);
  assign popcount33_en6z_core_150 = input_a[29] ^ input_a[0];
  assign popcount33_en6z_core_152 = ~input_a[4];
  assign popcount33_en6z_core_154 = input_a[0] & input_a[22];
  assign popcount33_en6z_core_156 = ~input_a[20];
  assign popcount33_en6z_core_157 = input_a[32] ^ input_a[26];
  assign popcount33_en6z_core_158 = input_a[2] | input_a[31];
  assign popcount33_en6z_core_160 = input_a[8] ^ input_a[29];
  assign popcount33_en6z_core_162 = input_a[4] | input_a[28];
  assign popcount33_en6z_core_163 = input_a[29] | input_a[11];
  assign popcount33_en6z_core_164 = input_a[0] & input_a[28];
  assign popcount33_en6z_core_166 = ~(input_a[4] ^ input_a[4]);
  assign popcount33_en6z_core_167 = ~(input_a[23] & input_a[11]);
  assign popcount33_en6z_core_168 = ~input_a[32];
  assign popcount33_en6z_core_170 = input_a[26] | input_a[19];
  assign popcount33_en6z_core_173 = input_a[5] | input_a[1];
  assign popcount33_en6z_core_176 = input_a[21] & input_a[32];
  assign popcount33_en6z_core_180 = input_a[16] & input_a[8];
  assign popcount33_en6z_core_182 = ~input_a[16];
  assign popcount33_en6z_core_183 = input_a[22] & input_a[6];
  assign popcount33_en6z_core_186 = input_a[15] ^ input_a[30];
  assign popcount33_en6z_core_187 = input_a[8] ^ input_a[15];
  assign popcount33_en6z_core_188 = input_a[2] & input_a[16];
  assign popcount33_en6z_core_189 = input_a[29] ^ input_a[20];
  assign popcount33_en6z_core_193 = ~input_a[11];
  assign popcount33_en6z_core_194 = input_a[11] | input_a[17];
  assign popcount33_en6z_core_195 = input_a[30] ^ input_a[10];
  assign popcount33_en6z_core_196 = ~(input_a[23] & input_a[2]);
  assign popcount33_en6z_core_197 = ~(input_a[26] | input_a[14]);
  assign popcount33_en6z_core_198 = ~(input_a[2] & input_a[7]);
  assign popcount33_en6z_core_199 = ~(input_a[12] | input_a[2]);
  assign popcount33_en6z_core_200_not = ~input_a[8];
  assign popcount33_en6z_core_203 = ~input_a[19];
  assign popcount33_en6z_core_204 = input_a[0] ^ input_a[14];
  assign popcount33_en6z_core_205 = input_a[1] ^ input_a[4];
  assign popcount33_en6z_core_206 = input_a[23] | input_a[15];
  assign popcount33_en6z_core_207 = input_a[27] ^ input_a[28];
  assign popcount33_en6z_core_209 = ~(input_a[16] | input_a[21]);
  assign popcount33_en6z_core_210 = input_a[6] | input_a[8];
  assign popcount33_en6z_core_212 = input_a[18] & input_a[4];
  assign popcount33_en6z_core_213 = ~(input_a[12] & input_a[21]);
  assign popcount33_en6z_core_214 = input_a[12] | input_a[17];
  assign popcount33_en6z_core_215 = input_a[26] ^ input_a[29];
  assign popcount33_en6z_core_218 = ~(input_a[9] | input_a[23]);
  assign popcount33_en6z_core_219 = input_a[20] & input_a[30];
  assign popcount33_en6z_core_221 = ~input_a[22];
  assign popcount33_en6z_core_222 = input_a[10] & input_a[22];
  assign popcount33_en6z_core_223 = input_a[31] ^ input_a[30];
  assign popcount33_en6z_core_224 = ~(input_a[24] & input_a[23]);
  assign popcount33_en6z_core_225 = input_a[1] | input_a[26];
  assign popcount33_en6z_core_226_not = ~input_a[0];
  assign popcount33_en6z_core_228 = ~(input_a[4] ^ input_a[1]);
  assign popcount33_en6z_core_229 = ~input_a[1];
  assign popcount33_en6z_core_230 = ~(input_a[13] ^ input_a[31]);
  assign popcount33_en6z_core_231 = input_a[10] | input_a[29];
  assign popcount33_en6z_core_233 = ~(input_a[0] | input_a[6]);
  assign popcount33_en6z_core_234 = ~(input_a[29] & input_a[27]);
  assign popcount33_en6z_core_237 = ~(input_a[25] & input_a[21]);

  assign popcount33_en6z_out[0] = 1'b1;
  assign popcount33_en6z_out[1] = input_a[28];
  assign popcount33_en6z_out[2] = input_a[17];
  assign popcount33_en6z_out[3] = 1'b0;
  assign popcount33_en6z_out[4] = 1'b1;
  assign popcount33_en6z_out[5] = 1'b0;
endmodule