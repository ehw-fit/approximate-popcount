// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.43472
// WCE=12.0
// EP=0.879866%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount20_py96(input [19:0] input_a, output [4:0] popcount20_py96_out);
  wire popcount20_py96_core_022;
  wire popcount20_py96_core_023;
  wire popcount20_py96_core_024;
  wire popcount20_py96_core_029;
  wire popcount20_py96_core_030;
  wire popcount20_py96_core_032;
  wire popcount20_py96_core_033;
  wire popcount20_py96_core_034;
  wire popcount20_py96_core_035;
  wire popcount20_py96_core_037;
  wire popcount20_py96_core_038;
  wire popcount20_py96_core_041_not;
  wire popcount20_py96_core_043;
  wire popcount20_py96_core_046;
  wire popcount20_py96_core_047;
  wire popcount20_py96_core_050;
  wire popcount20_py96_core_051;
  wire popcount20_py96_core_052;
  wire popcount20_py96_core_053;
  wire popcount20_py96_core_055;
  wire popcount20_py96_core_058;
  wire popcount20_py96_core_060;
  wire popcount20_py96_core_061;
  wire popcount20_py96_core_062;
  wire popcount20_py96_core_065;
  wire popcount20_py96_core_066;
  wire popcount20_py96_core_069;
  wire popcount20_py96_core_070;
  wire popcount20_py96_core_071;
  wire popcount20_py96_core_072;
  wire popcount20_py96_core_073;
  wire popcount20_py96_core_075;
  wire popcount20_py96_core_076;
  wire popcount20_py96_core_078;
  wire popcount20_py96_core_081;
  wire popcount20_py96_core_082;
  wire popcount20_py96_core_083;
  wire popcount20_py96_core_084;
  wire popcount20_py96_core_085;
  wire popcount20_py96_core_086;
  wire popcount20_py96_core_089;
  wire popcount20_py96_core_090;
  wire popcount20_py96_core_092;
  wire popcount20_py96_core_093;
  wire popcount20_py96_core_096;
  wire popcount20_py96_core_097;
  wire popcount20_py96_core_098;
  wire popcount20_py96_core_099;
  wire popcount20_py96_core_100;
  wire popcount20_py96_core_101;
  wire popcount20_py96_core_104_not;
  wire popcount20_py96_core_106;
  wire popcount20_py96_core_107;
  wire popcount20_py96_core_109_not;
  wire popcount20_py96_core_112;
  wire popcount20_py96_core_113;
  wire popcount20_py96_core_114;
  wire popcount20_py96_core_115;
  wire popcount20_py96_core_120;
  wire popcount20_py96_core_121;
  wire popcount20_py96_core_122;
  wire popcount20_py96_core_123;
  wire popcount20_py96_core_124;
  wire popcount20_py96_core_125_not;
  wire popcount20_py96_core_126;
  wire popcount20_py96_core_130;
  wire popcount20_py96_core_132;
  wire popcount20_py96_core_133;
  wire popcount20_py96_core_135;
  wire popcount20_py96_core_140;
  wire popcount20_py96_core_144;
  wire popcount20_py96_core_145;

  assign popcount20_py96_core_022 = input_a[6] ^ input_a[15];
  assign popcount20_py96_core_023 = ~input_a[16];
  assign popcount20_py96_core_024 = input_a[2] | input_a[10];
  assign popcount20_py96_core_029 = input_a[10] | input_a[7];
  assign popcount20_py96_core_030 = ~input_a[7];
  assign popcount20_py96_core_032 = input_a[3] & input_a[1];
  assign popcount20_py96_core_033 = ~(input_a[3] | input_a[3]);
  assign popcount20_py96_core_034 = input_a[8] | input_a[19];
  assign popcount20_py96_core_035 = ~(input_a[7] & input_a[10]);
  assign popcount20_py96_core_037 = ~(input_a[6] & input_a[0]);
  assign popcount20_py96_core_038 = ~(input_a[4] ^ input_a[3]);
  assign popcount20_py96_core_041_not = ~input_a[4];
  assign popcount20_py96_core_043 = input_a[14] ^ input_a[2];
  assign popcount20_py96_core_046 = input_a[0] | input_a[0];
  assign popcount20_py96_core_047 = input_a[11] & input_a[16];
  assign popcount20_py96_core_050 = input_a[1] ^ input_a[17];
  assign popcount20_py96_core_051 = input_a[19] & input_a[11];
  assign popcount20_py96_core_052 = input_a[14] | input_a[0];
  assign popcount20_py96_core_053 = ~input_a[10];
  assign popcount20_py96_core_055 = ~(input_a[9] | input_a[11]);
  assign popcount20_py96_core_058 = ~(input_a[16] & input_a[1]);
  assign popcount20_py96_core_060 = input_a[18] & input_a[3];
  assign popcount20_py96_core_061 = ~(input_a[19] | input_a[4]);
  assign popcount20_py96_core_062 = input_a[8] ^ input_a[14];
  assign popcount20_py96_core_065 = input_a[17] | input_a[2];
  assign popcount20_py96_core_066 = ~(input_a[4] | input_a[4]);
  assign popcount20_py96_core_069 = ~(input_a[15] | input_a[4]);
  assign popcount20_py96_core_070 = ~(input_a[7] & input_a[14]);
  assign popcount20_py96_core_071 = ~(input_a[18] & input_a[8]);
  assign popcount20_py96_core_072 = ~(input_a[18] ^ input_a[0]);
  assign popcount20_py96_core_073 = input_a[6] & input_a[3];
  assign popcount20_py96_core_075 = input_a[0] ^ input_a[10];
  assign popcount20_py96_core_076 = input_a[0] & input_a[8];
  assign popcount20_py96_core_078 = ~input_a[3];
  assign popcount20_py96_core_081 = input_a[6] & input_a[0];
  assign popcount20_py96_core_082 = input_a[19] | input_a[10];
  assign popcount20_py96_core_083 = input_a[16] ^ input_a[13];
  assign popcount20_py96_core_084 = ~(input_a[19] ^ input_a[12]);
  assign popcount20_py96_core_085 = ~input_a[4];
  assign popcount20_py96_core_086 = input_a[2] | input_a[17];
  assign popcount20_py96_core_089 = ~input_a[8];
  assign popcount20_py96_core_090 = input_a[18] & input_a[9];
  assign popcount20_py96_core_092 = input_a[3] | input_a[15];
  assign popcount20_py96_core_093 = ~(input_a[11] & input_a[7]);
  assign popcount20_py96_core_096 = input_a[0] & input_a[14];
  assign popcount20_py96_core_097 = input_a[3] & input_a[17];
  assign popcount20_py96_core_098 = ~(input_a[15] ^ input_a[18]);
  assign popcount20_py96_core_099 = input_a[9] ^ input_a[17];
  assign popcount20_py96_core_100 = input_a[2] | input_a[4];
  assign popcount20_py96_core_101 = input_a[8] & input_a[4];
  assign popcount20_py96_core_104_not = ~input_a[17];
  assign popcount20_py96_core_106 = ~input_a[8];
  assign popcount20_py96_core_107 = input_a[1] & input_a[19];
  assign popcount20_py96_core_109_not = ~input_a[14];
  assign popcount20_py96_core_112 = input_a[12] ^ input_a[15];
  assign popcount20_py96_core_113 = ~(input_a[18] | input_a[4]);
  assign popcount20_py96_core_114 = ~(input_a[11] | input_a[11]);
  assign popcount20_py96_core_115 = ~(input_a[7] & input_a[18]);
  assign popcount20_py96_core_120 = ~(input_a[17] ^ input_a[19]);
  assign popcount20_py96_core_121 = ~(input_a[1] | input_a[16]);
  assign popcount20_py96_core_122 = ~(input_a[10] | input_a[5]);
  assign popcount20_py96_core_123 = ~(input_a[10] | input_a[1]);
  assign popcount20_py96_core_124 = input_a[17] & input_a[18];
  assign popcount20_py96_core_125_not = ~input_a[15];
  assign popcount20_py96_core_126 = ~(input_a[4] & input_a[8]);
  assign popcount20_py96_core_130 = ~(input_a[0] & input_a[17]);
  assign popcount20_py96_core_132 = input_a[0] & input_a[11];
  assign popcount20_py96_core_133 = ~(input_a[16] & input_a[8]);
  assign popcount20_py96_core_135 = input_a[3] & input_a[12];
  assign popcount20_py96_core_140 = ~(input_a[3] | input_a[16]);
  assign popcount20_py96_core_144 = ~(input_a[0] | input_a[1]);
  assign popcount20_py96_core_145 = input_a[15] & input_a[12];

  assign popcount20_py96_out[0] = input_a[12];
  assign popcount20_py96_out[1] = 1'b0;
  assign popcount20_py96_out[2] = 1'b0;
  assign popcount20_py96_out[3] = 1'b1;
  assign popcount20_py96_out[4] = 1'b0;
endmodule