// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.29536
// WCE=38.0
// EP=0.925179%
// Printed PDK parameters:
//  Area=120648059.0
//  Delay=90558128.0
//  Power=7136000.0

module popcount43_r54b(input [42:0] input_a, output [5:0] popcount43_r54b_out);
  wire popcount43_r54b_core_046;
  wire popcount43_r54b_core_047;
  wire popcount43_r54b_core_048;
  wire popcount43_r54b_core_049;
  wire popcount43_r54b_core_050;
  wire popcount43_r54b_core_051;
  wire popcount43_r54b_core_055;
  wire popcount43_r54b_core_057;
  wire popcount43_r54b_core_062;
  wire popcount43_r54b_core_064;
  wire popcount43_r54b_core_065;
  wire popcount43_r54b_core_067;
  wire popcount43_r54b_core_068;
  wire popcount43_r54b_core_069;
  wire popcount43_r54b_core_080;
  wire popcount43_r54b_core_081;
  wire popcount43_r54b_core_082;
  wire popcount43_r54b_core_084;
  wire popcount43_r54b_core_096;
  wire popcount43_r54b_core_098;
  wire popcount43_r54b_core_099;
  wire popcount43_r54b_core_100;
  wire popcount43_r54b_core_101;
  wire popcount43_r54b_core_102;
  wire popcount43_r54b_core_103;
  wire popcount43_r54b_core_104;
  wire popcount43_r54b_core_105;
  wire popcount43_r54b_core_106;
  wire popcount43_r54b_core_107;
  wire popcount43_r54b_core_108;
  wire popcount43_r54b_core_109;
  wire popcount43_r54b_core_110;
  wire popcount43_r54b_core_111;
  wire popcount43_r54b_core_112;
  wire popcount43_r54b_core_113;
  wire popcount43_r54b_core_114;
  wire popcount43_r54b_core_115;
  wire popcount43_r54b_core_116;
  wire popcount43_r54b_core_117;
  wire popcount43_r54b_core_118;
  wire popcount43_r54b_core_119;
  wire popcount43_r54b_core_120;
  wire popcount43_r54b_core_121;
  wire popcount43_r54b_core_122;
  wire popcount43_r54b_core_123;
  wire popcount43_r54b_core_124;
  wire popcount43_r54b_core_125;
  wire popcount43_r54b_core_126;
  wire popcount43_r54b_core_127;
  wire popcount43_r54b_core_128;
  wire popcount43_r54b_core_129;
  wire popcount43_r54b_core_130;
  wire popcount43_r54b_core_131;
  wire popcount43_r54b_core_132;
  wire popcount43_r54b_core_133;
  wire popcount43_r54b_core_134;
  wire popcount43_r54b_core_135;
  wire popcount43_r54b_core_136;
  wire popcount43_r54b_core_137;
  wire popcount43_r54b_core_138;
  wire popcount43_r54b_core_139;
  wire popcount43_r54b_core_140;
  wire popcount43_r54b_core_141;
  wire popcount43_r54b_core_142;
  wire popcount43_r54b_core_143;
  wire popcount43_r54b_core_144;
  wire popcount43_r54b_core_145;
  wire popcount43_r54b_core_146;
  wire popcount43_r54b_core_147;
  wire popcount43_r54b_core_148;
  wire popcount43_r54b_core_149;
  wire popcount43_r54b_core_151;
  wire popcount43_r54b_core_152;
  wire popcount43_r54b_core_154;
  wire popcount43_r54b_core_155;
  wire popcount43_r54b_core_156;
  wire popcount43_r54b_core_157;
  wire popcount43_r54b_core_158;
  wire popcount43_r54b_core_159;
  wire popcount43_r54b_core_160;
  wire popcount43_r54b_core_161;
  wire popcount43_r54b_core_162;
  wire popcount43_r54b_core_163;
  wire popcount43_r54b_core_164;
  wire popcount43_r54b_core_165;
  wire popcount43_r54b_core_168;
  wire popcount43_r54b_core_169;
  wire popcount43_r54b_core_174;
  wire popcount43_r54b_core_176;
  wire popcount43_r54b_core_177;
  wire popcount43_r54b_core_178;
  wire popcount43_r54b_core_180;
  wire popcount43_r54b_core_181;
  wire popcount43_r54b_core_182;
  wire popcount43_r54b_core_183;
  wire popcount43_r54b_core_184;
  wire popcount43_r54b_core_185;
  wire popcount43_r54b_core_187;
  wire popcount43_r54b_core_188;
  wire popcount43_r54b_core_189;
  wire popcount43_r54b_core_190;
  wire popcount43_r54b_core_191;
  wire popcount43_r54b_core_192;
  wire popcount43_r54b_core_193;
  wire popcount43_r54b_core_195;
  wire popcount43_r54b_core_196;
  wire popcount43_r54b_core_199;
  wire popcount43_r54b_core_200;
  wire popcount43_r54b_core_201;
  wire popcount43_r54b_core_202;
  wire popcount43_r54b_core_203;
  wire popcount43_r54b_core_204;
  wire popcount43_r54b_core_205;
  wire popcount43_r54b_core_206;
  wire popcount43_r54b_core_207;
  wire popcount43_r54b_core_208;
  wire popcount43_r54b_core_210;
  wire popcount43_r54b_core_211;
  wire popcount43_r54b_core_214;
  wire popcount43_r54b_core_215;
  wire popcount43_r54b_core_217;
  wire popcount43_r54b_core_218;
  wire popcount43_r54b_core_221;
  wire popcount43_r54b_core_222;
  wire popcount43_r54b_core_224;
  wire popcount43_r54b_core_225;
  wire popcount43_r54b_core_226;
  wire popcount43_r54b_core_227;
  wire popcount43_r54b_core_228;
  wire popcount43_r54b_core_229;
  wire popcount43_r54b_core_231;
  wire popcount43_r54b_core_234;
  wire popcount43_r54b_core_235;
  wire popcount43_r54b_core_236;
  wire popcount43_r54b_core_238;
  wire popcount43_r54b_core_239;
  wire popcount43_r54b_core_242;
  wire popcount43_r54b_core_243;
  wire popcount43_r54b_core_244;
  wire popcount43_r54b_core_245;
  wire popcount43_r54b_core_246;
  wire popcount43_r54b_core_247;
  wire popcount43_r54b_core_248;
  wire popcount43_r54b_core_251;
  wire popcount43_r54b_core_252;
  wire popcount43_r54b_core_255;
  wire popcount43_r54b_core_256;
  wire popcount43_r54b_core_257;
  wire popcount43_r54b_core_258;
  wire popcount43_r54b_core_259;
  wire popcount43_r54b_core_260;
  wire popcount43_r54b_core_261;
  wire popcount43_r54b_core_262;
  wire popcount43_r54b_core_264;
  wire popcount43_r54b_core_265;
  wire popcount43_r54b_core_266;
  wire popcount43_r54b_core_267;
  wire popcount43_r54b_core_270;
  wire popcount43_r54b_core_271;
  wire popcount43_r54b_core_272;
  wire popcount43_r54b_core_273;
  wire popcount43_r54b_core_274;
  wire popcount43_r54b_core_275;
  wire popcount43_r54b_core_276;
  wire popcount43_r54b_core_277;
  wire popcount43_r54b_core_278;
  wire popcount43_r54b_core_279;
  wire popcount43_r54b_core_280;
  wire popcount43_r54b_core_281;
  wire popcount43_r54b_core_282;
  wire popcount43_r54b_core_283;
  wire popcount43_r54b_core_284;
  wire popcount43_r54b_core_285;
  wire popcount43_r54b_core_286;
  wire popcount43_r54b_core_289;
  wire popcount43_r54b_core_290;
  wire popcount43_r54b_core_292;
  wire popcount43_r54b_core_293;
  wire popcount43_r54b_core_294;
  wire popcount43_r54b_core_295;
  wire popcount43_r54b_core_296;
  wire popcount43_r54b_core_297;
  wire popcount43_r54b_core_298;
  wire popcount43_r54b_core_299;
  wire popcount43_r54b_core_300;
  wire popcount43_r54b_core_301;
  wire popcount43_r54b_core_302;
  wire popcount43_r54b_core_303;
  wire popcount43_r54b_core_304;
  wire popcount43_r54b_core_305;
  wire popcount43_r54b_core_306;
  wire popcount43_r54b_core_307;
  wire popcount43_r54b_core_308;
  wire popcount43_r54b_core_312;
  wire popcount43_r54b_core_313;
  wire popcount43_r54b_core_314;
  wire popcount43_r54b_core_315;
  wire popcount43_r54b_core_317;
  wire popcount43_r54b_core_318;
  wire popcount43_r54b_core_319;
  wire popcount43_r54b_core_320;
  wire popcount43_r54b_core_321;
  wire popcount43_r54b_core_322;
  wire popcount43_r54b_core_323;
  wire popcount43_r54b_core_324;
  wire popcount43_r54b_core_325;
  wire popcount43_r54b_core_326;
  wire popcount43_r54b_core_327;
  wire popcount43_r54b_core_328;
  wire popcount43_r54b_core_329;
  wire popcount43_r54b_core_330;
  wire popcount43_r54b_core_331;
  wire popcount43_r54b_core_332;
  wire popcount43_r54b_core_333;
  wire popcount43_r54b_core_334;
  wire popcount43_r54b_core_335;
  wire popcount43_r54b_core_337;

  assign popcount43_r54b_core_046 = input_a[0] & input_a[1];
  assign popcount43_r54b_core_047 = input_a[3] | input_a[4];
  assign popcount43_r54b_core_048 = input_a[3] & input_a[41];
  assign popcount43_r54b_core_049 = input_a[2] | popcount43_r54b_core_047;
  assign popcount43_r54b_core_050 = input_a[2] & popcount43_r54b_core_047;
  assign popcount43_r54b_core_051 = popcount43_r54b_core_048 ^ popcount43_r54b_core_050;
  assign popcount43_r54b_core_055 = input_a[23] ^ popcount43_r54b_core_051;
  assign popcount43_r54b_core_057 = popcount43_r54b_core_055 ^ input_a[34];
  assign popcount43_r54b_core_062 = input_a[5] ^ input_a[6];
  assign popcount43_r54b_core_064 = input_a[15] ^ input_a[4];
  assign popcount43_r54b_core_065 = input_a[8] & input_a[9];
  assign popcount43_r54b_core_067 = input_a[7] & input_a[9];
  assign popcount43_r54b_core_068 = popcount43_r54b_core_065 ^ popcount43_r54b_core_067;
  assign popcount43_r54b_core_069 = popcount43_r54b_core_065 & popcount43_r54b_core_067;
  assign popcount43_r54b_core_080 = input_a[8] & input_a[12];
  assign popcount43_r54b_core_081 = popcount43_r54b_core_057 ^ input_a[25];
  assign popcount43_r54b_core_082 = popcount43_r54b_core_057 & input_a[25];
  assign popcount43_r54b_core_084 = input_a[19] & popcount43_r54b_core_080;
  assign popcount43_r54b_core_096 = input_a[10] ^ input_a[11];
  assign popcount43_r54b_core_098 = input_a[13] ^ input_a[14];
  assign popcount43_r54b_core_099 = ~(input_a[13] | input_a[14]);
  assign popcount43_r54b_core_100 = input_a[12] ^ popcount43_r54b_core_098;
  assign popcount43_r54b_core_101 = input_a[12] & popcount43_r54b_core_098;
  assign popcount43_r54b_core_102 = popcount43_r54b_core_099 ^ popcount43_r54b_core_101;
  assign popcount43_r54b_core_103 = popcount43_r54b_core_099 & popcount43_r54b_core_101;
  assign popcount43_r54b_core_104 = ~popcount43_r54b_core_096;
  assign popcount43_r54b_core_105 = ~(popcount43_r54b_core_096 | popcount43_r54b_core_100);
  assign popcount43_r54b_core_106 = input_a[11] ^ popcount43_r54b_core_102;
  assign popcount43_r54b_core_107 = input_a[11] & popcount43_r54b_core_102;
  assign popcount43_r54b_core_108 = popcount43_r54b_core_106 ^ popcount43_r54b_core_105;
  assign popcount43_r54b_core_109 = popcount43_r54b_core_106 & popcount43_r54b_core_105;
  assign popcount43_r54b_core_110 = popcount43_r54b_core_107 | popcount43_r54b_core_109;
  assign popcount43_r54b_core_111 = popcount43_r54b_core_103 ^ popcount43_r54b_core_110;
  assign popcount43_r54b_core_112 = popcount43_r54b_core_103 & popcount43_r54b_core_110;
  assign popcount43_r54b_core_113 = input_a[16] ^ input_a[17];
  assign popcount43_r54b_core_114 = input_a[16] & input_a[17];
  assign popcount43_r54b_core_115 = input_a[15] ^ popcount43_r54b_core_113;
  assign popcount43_r54b_core_116 = input_a[15] & popcount43_r54b_core_113;
  assign popcount43_r54b_core_117 = popcount43_r54b_core_114 ^ popcount43_r54b_core_116;
  assign popcount43_r54b_core_118 = popcount43_r54b_core_114 & popcount43_r54b_core_116;
  assign popcount43_r54b_core_119 = input_a[19] ^ input_a[20];
  assign popcount43_r54b_core_120 = input_a[19] & input_a[20];
  assign popcount43_r54b_core_121 = input_a[18] ^ popcount43_r54b_core_119;
  assign popcount43_r54b_core_122 = input_a[18] & popcount43_r54b_core_119;
  assign popcount43_r54b_core_123 = popcount43_r54b_core_120 ^ popcount43_r54b_core_122;
  assign popcount43_r54b_core_124 = popcount43_r54b_core_120 & popcount43_r54b_core_122;
  assign popcount43_r54b_core_125 = popcount43_r54b_core_115 ^ popcount43_r54b_core_121;
  assign popcount43_r54b_core_126 = popcount43_r54b_core_115 & popcount43_r54b_core_121;
  assign popcount43_r54b_core_127 = popcount43_r54b_core_117 ^ popcount43_r54b_core_123;
  assign popcount43_r54b_core_128 = popcount43_r54b_core_117 & popcount43_r54b_core_123;
  assign popcount43_r54b_core_129 = popcount43_r54b_core_127 ^ popcount43_r54b_core_126;
  assign popcount43_r54b_core_130 = popcount43_r54b_core_127 & popcount43_r54b_core_126;
  assign popcount43_r54b_core_131 = popcount43_r54b_core_128 | popcount43_r54b_core_130;
  assign popcount43_r54b_core_132 = popcount43_r54b_core_118 ^ popcount43_r54b_core_124;
  assign popcount43_r54b_core_133 = popcount43_r54b_core_118 & popcount43_r54b_core_124;
  assign popcount43_r54b_core_134 = popcount43_r54b_core_132 ^ popcount43_r54b_core_131;
  assign popcount43_r54b_core_135 = popcount43_r54b_core_132 & popcount43_r54b_core_131;
  assign popcount43_r54b_core_136 = popcount43_r54b_core_133 | popcount43_r54b_core_135;
  assign popcount43_r54b_core_137 = popcount43_r54b_core_104 ^ popcount43_r54b_core_125;
  assign popcount43_r54b_core_138 = popcount43_r54b_core_104 & popcount43_r54b_core_125;
  assign popcount43_r54b_core_139 = popcount43_r54b_core_108 ^ popcount43_r54b_core_129;
  assign popcount43_r54b_core_140 = popcount43_r54b_core_108 & popcount43_r54b_core_129;
  assign popcount43_r54b_core_141 = popcount43_r54b_core_139 ^ popcount43_r54b_core_138;
  assign popcount43_r54b_core_142 = input_a[7] & popcount43_r54b_core_138;
  assign popcount43_r54b_core_143 = popcount43_r54b_core_140 | popcount43_r54b_core_142;
  assign popcount43_r54b_core_144 = popcount43_r54b_core_111 ^ popcount43_r54b_core_134;
  assign popcount43_r54b_core_145 = popcount43_r54b_core_111 & popcount43_r54b_core_134;
  assign popcount43_r54b_core_146 = popcount43_r54b_core_144 ^ popcount43_r54b_core_143;
  assign popcount43_r54b_core_147 = popcount43_r54b_core_144 & popcount43_r54b_core_143;
  assign popcount43_r54b_core_148 = popcount43_r54b_core_145 | popcount43_r54b_core_147;
  assign popcount43_r54b_core_149 = popcount43_r54b_core_112 ^ popcount43_r54b_core_136;
  assign popcount43_r54b_core_151 = popcount43_r54b_core_149 | popcount43_r54b_core_148;
  assign popcount43_r54b_core_152 = popcount43_r54b_core_149 & popcount43_r54b_core_148;
  assign popcount43_r54b_core_154 = input_a[13] ^ popcount43_r54b_core_137;
  assign popcount43_r54b_core_155 = input_a[13] & popcount43_r54b_core_137;
  assign popcount43_r54b_core_156 = popcount43_r54b_core_081 ^ popcount43_r54b_core_141;
  assign popcount43_r54b_core_157 = popcount43_r54b_core_081 & popcount43_r54b_core_141;
  assign popcount43_r54b_core_158 = popcount43_r54b_core_156 ^ popcount43_r54b_core_155;
  assign popcount43_r54b_core_159 = popcount43_r54b_core_156 & popcount43_r54b_core_155;
  assign popcount43_r54b_core_160 = popcount43_r54b_core_157 | popcount43_r54b_core_159;
  assign popcount43_r54b_core_161 = popcount43_r54b_core_069 ^ popcount43_r54b_core_146;
  assign popcount43_r54b_core_162 = popcount43_r54b_core_069 & popcount43_r54b_core_146;
  assign popcount43_r54b_core_163 = popcount43_r54b_core_161 ^ popcount43_r54b_core_160;
  assign popcount43_r54b_core_164 = popcount43_r54b_core_161 & popcount43_r54b_core_160;
  assign popcount43_r54b_core_165 = popcount43_r54b_core_162 | popcount43_r54b_core_164;
  assign popcount43_r54b_core_168 = popcount43_r54b_core_151 ^ popcount43_r54b_core_165;
  assign popcount43_r54b_core_169 = popcount43_r54b_core_151 & popcount43_r54b_core_165;
  assign popcount43_r54b_core_174 = popcount43_r54b_core_152 | popcount43_r54b_core_169;
  assign popcount43_r54b_core_176 = input_a[21] ^ input_a[22];
  assign popcount43_r54b_core_177 = input_a[21] & input_a[22];
  assign popcount43_r54b_core_178 = input_a[24] ^ input_a[25];
  assign popcount43_r54b_core_180 = input_a[23] ^ popcount43_r54b_core_178;
  assign popcount43_r54b_core_181 = input_a[23] & popcount43_r54b_core_178;
  assign popcount43_r54b_core_182 = input_a[24] ^ popcount43_r54b_core_181;
  assign popcount43_r54b_core_183 = input_a[24] & popcount43_r54b_core_181;
  assign popcount43_r54b_core_184 = popcount43_r54b_core_176 ^ popcount43_r54b_core_180;
  assign popcount43_r54b_core_185 = popcount43_r54b_core_176 & popcount43_r54b_core_180;
  assign popcount43_r54b_core_187 = ~input_a[20];
  assign popcount43_r54b_core_188 = popcount43_r54b_core_177 ^ popcount43_r54b_core_185;
  assign popcount43_r54b_core_189 = popcount43_r54b_core_177 & popcount43_r54b_core_185;
  assign popcount43_r54b_core_190 = input_a[42] | input_a[16];
  assign popcount43_r54b_core_191 = popcount43_r54b_core_183 ^ popcount43_r54b_core_190;
  assign popcount43_r54b_core_192 = popcount43_r54b_core_183 & popcount43_r54b_core_190;
  assign popcount43_r54b_core_193 = input_a[9] ^ input_a[28];
  assign popcount43_r54b_core_195 = input_a[26] ^ popcount43_r54b_core_193;
  assign popcount43_r54b_core_196 = input_a[26] & popcount43_r54b_core_193;
  assign popcount43_r54b_core_199 = input_a[27] ^ input_a[31];
  assign popcount43_r54b_core_200 = input_a[30] & input_a[31];
  assign popcount43_r54b_core_201 = input_a[29] ^ popcount43_r54b_core_199;
  assign popcount43_r54b_core_202 = input_a[29] & popcount43_r54b_core_199;
  assign popcount43_r54b_core_203 = input_a[5] ^ popcount43_r54b_core_202;
  assign popcount43_r54b_core_204 = popcount43_r54b_core_200 & input_a[38];
  assign popcount43_r54b_core_205 = popcount43_r54b_core_195 ^ popcount43_r54b_core_201;
  assign popcount43_r54b_core_206 = popcount43_r54b_core_195 & popcount43_r54b_core_201;
  assign popcount43_r54b_core_207 = popcount43_r54b_core_196 ^ popcount43_r54b_core_203;
  assign popcount43_r54b_core_208 = popcount43_r54b_core_196 & popcount43_r54b_core_203;
  assign popcount43_r54b_core_210 = popcount43_r54b_core_207 & popcount43_r54b_core_206;
  assign popcount43_r54b_core_211 = input_a[13] | popcount43_r54b_core_210;
  assign popcount43_r54b_core_214 = input_a[7] ^ popcount43_r54b_core_211;
  assign popcount43_r54b_core_215 = input_a[7] & popcount43_r54b_core_211;
  assign popcount43_r54b_core_217 = popcount43_r54b_core_184 ^ popcount43_r54b_core_205;
  assign popcount43_r54b_core_218 = popcount43_r54b_core_184 & popcount43_r54b_core_205;
  assign popcount43_r54b_core_221 = popcount43_r54b_core_188 ^ popcount43_r54b_core_218;
  assign popcount43_r54b_core_222 = popcount43_r54b_core_188 & popcount43_r54b_core_218;
  assign popcount43_r54b_core_224 = popcount43_r54b_core_191 ^ popcount43_r54b_core_214;
  assign popcount43_r54b_core_225 = popcount43_r54b_core_191 & popcount43_r54b_core_214;
  assign popcount43_r54b_core_226 = popcount43_r54b_core_224 ^ popcount43_r54b_core_222;
  assign popcount43_r54b_core_227 = popcount43_r54b_core_224 & popcount43_r54b_core_222;
  assign popcount43_r54b_core_228 = popcount43_r54b_core_225 | popcount43_r54b_core_227;
  assign popcount43_r54b_core_229 = popcount43_r54b_core_192 ^ popcount43_r54b_core_215;
  assign popcount43_r54b_core_231 = popcount43_r54b_core_229 ^ popcount43_r54b_core_228;
  assign popcount43_r54b_core_234 = input_a[32] ^ input_a[28];
  assign popcount43_r54b_core_235 = input_a[38] & input_a[30];
  assign popcount43_r54b_core_236 = input_a[35] ^ input_a[36];
  assign popcount43_r54b_core_238 = input_a[34] ^ input_a[33];
  assign popcount43_r54b_core_239 = input_a[34] & input_a[0];
  assign popcount43_r54b_core_242 = input_a[10] ^ popcount43_r54b_core_238;
  assign popcount43_r54b_core_243 = input_a[2] & popcount43_r54b_core_238;
  assign popcount43_r54b_core_244 = popcount43_r54b_core_235 ^ input_a[14];
  assign popcount43_r54b_core_245 = popcount43_r54b_core_235 & popcount43_r54b_core_239;
  assign popcount43_r54b_core_246 = popcount43_r54b_core_244 ^ popcount43_r54b_core_243;
  assign popcount43_r54b_core_247 = popcount43_r54b_core_244 & popcount43_r54b_core_243;
  assign popcount43_r54b_core_248 = popcount43_r54b_core_245 | popcount43_r54b_core_247;
  assign popcount43_r54b_core_251 = input_a[38] ^ input_a[39];
  assign popcount43_r54b_core_252 = input_a[38] & input_a[39];
  assign popcount43_r54b_core_255 = popcount43_r54b_core_252 ^ input_a[37];
  assign popcount43_r54b_core_256 = popcount43_r54b_core_252 & input_a[37];
  assign popcount43_r54b_core_257 = input_a[41] ^ input_a[42];
  assign popcount43_r54b_core_258 = input_a[41] & input_a[42];
  assign popcount43_r54b_core_259 = input_a[40] ^ input_a[40];
  assign popcount43_r54b_core_260 = input_a[40] & popcount43_r54b_core_257;
  assign popcount43_r54b_core_261 = popcount43_r54b_core_258 ^ popcount43_r54b_core_260;
  assign popcount43_r54b_core_262 = popcount43_r54b_core_258 & popcount43_r54b_core_260;
  assign popcount43_r54b_core_264 = input_a[19] & popcount43_r54b_core_259;
  assign popcount43_r54b_core_265 = popcount43_r54b_core_255 ^ popcount43_r54b_core_261;
  assign popcount43_r54b_core_266 = popcount43_r54b_core_255 & popcount43_r54b_core_261;
  assign popcount43_r54b_core_267 = popcount43_r54b_core_265 ^ popcount43_r54b_core_264;
  assign popcount43_r54b_core_270 = popcount43_r54b_core_256 ^ popcount43_r54b_core_262;
  assign popcount43_r54b_core_271 = popcount43_r54b_core_256 & popcount43_r54b_core_262;
  assign popcount43_r54b_core_272 = popcount43_r54b_core_270 ^ popcount43_r54b_core_266;
  assign popcount43_r54b_core_273 = popcount43_r54b_core_270 & popcount43_r54b_core_266;
  assign popcount43_r54b_core_274 = popcount43_r54b_core_271 | popcount43_r54b_core_273;
  assign popcount43_r54b_core_275 = popcount43_r54b_core_242 ^ popcount43_r54b_core_259;
  assign popcount43_r54b_core_276 = popcount43_r54b_core_242 & popcount43_r54b_core_259;
  assign popcount43_r54b_core_277 = popcount43_r54b_core_246 ^ popcount43_r54b_core_267;
  assign popcount43_r54b_core_278 = popcount43_r54b_core_246 & popcount43_r54b_core_267;
  assign popcount43_r54b_core_279 = popcount43_r54b_core_277 ^ popcount43_r54b_core_276;
  assign popcount43_r54b_core_280 = popcount43_r54b_core_277 & popcount43_r54b_core_276;
  assign popcount43_r54b_core_281 = popcount43_r54b_core_278 | popcount43_r54b_core_280;
  assign popcount43_r54b_core_282 = popcount43_r54b_core_248 ^ popcount43_r54b_core_272;
  assign popcount43_r54b_core_283 = popcount43_r54b_core_248 & popcount43_r54b_core_272;
  assign popcount43_r54b_core_284 = popcount43_r54b_core_282 ^ popcount43_r54b_core_281;
  assign popcount43_r54b_core_285 = popcount43_r54b_core_282 & popcount43_r54b_core_281;
  assign popcount43_r54b_core_286 = popcount43_r54b_core_283 | popcount43_r54b_core_285;
  assign popcount43_r54b_core_289 = popcount43_r54b_core_274 ^ popcount43_r54b_core_286;
  assign popcount43_r54b_core_290 = popcount43_r54b_core_274 & popcount43_r54b_core_286;
  assign popcount43_r54b_core_292 = popcount43_r54b_core_217 ^ input_a[36];
  assign popcount43_r54b_core_293 = popcount43_r54b_core_217 & popcount43_r54b_core_275;
  assign popcount43_r54b_core_294 = popcount43_r54b_core_221 ^ popcount43_r54b_core_279;
  assign popcount43_r54b_core_295 = popcount43_r54b_core_221 & popcount43_r54b_core_279;
  assign popcount43_r54b_core_296 = popcount43_r54b_core_294 ^ popcount43_r54b_core_293;
  assign popcount43_r54b_core_297 = popcount43_r54b_core_294 & popcount43_r54b_core_293;
  assign popcount43_r54b_core_298 = popcount43_r54b_core_295 | popcount43_r54b_core_297;
  assign popcount43_r54b_core_299 = popcount43_r54b_core_226 ^ popcount43_r54b_core_284;
  assign popcount43_r54b_core_300 = popcount43_r54b_core_226 & popcount43_r54b_core_284;
  assign popcount43_r54b_core_301 = popcount43_r54b_core_299 ^ popcount43_r54b_core_298;
  assign popcount43_r54b_core_302 = popcount43_r54b_core_299 & popcount43_r54b_core_298;
  assign popcount43_r54b_core_303 = popcount43_r54b_core_300 | popcount43_r54b_core_302;
  assign popcount43_r54b_core_304 = popcount43_r54b_core_231 ^ popcount43_r54b_core_289;
  assign popcount43_r54b_core_305 = popcount43_r54b_core_231 & popcount43_r54b_core_289;
  assign popcount43_r54b_core_306 = popcount43_r54b_core_304 ^ popcount43_r54b_core_303;
  assign popcount43_r54b_core_307 = popcount43_r54b_core_304 & popcount43_r54b_core_303;
  assign popcount43_r54b_core_308 = popcount43_r54b_core_305 | popcount43_r54b_core_307;
  assign popcount43_r54b_core_312 = input_a[35] & popcount43_r54b_core_308;
  assign popcount43_r54b_core_313 = input_a[12] | popcount43_r54b_core_312;
  assign popcount43_r54b_core_314 = popcount43_r54b_core_154 ^ popcount43_r54b_core_292;
  assign popcount43_r54b_core_315 = popcount43_r54b_core_154 & input_a[6];
  assign popcount43_r54b_core_317 = popcount43_r54b_core_158 & popcount43_r54b_core_296;
  assign popcount43_r54b_core_318 = popcount43_r54b_core_158 ^ popcount43_r54b_core_315;
  assign popcount43_r54b_core_319 = popcount43_r54b_core_158 & popcount43_r54b_core_315;
  assign popcount43_r54b_core_320 = popcount43_r54b_core_317 | popcount43_r54b_core_319;
  assign popcount43_r54b_core_321 = popcount43_r54b_core_163 ^ popcount43_r54b_core_301;
  assign popcount43_r54b_core_322 = popcount43_r54b_core_163 & popcount43_r54b_core_301;
  assign popcount43_r54b_core_323 = popcount43_r54b_core_321 ^ popcount43_r54b_core_320;
  assign popcount43_r54b_core_324 = popcount43_r54b_core_321 & popcount43_r54b_core_320;
  assign popcount43_r54b_core_325 = popcount43_r54b_core_322 | popcount43_r54b_core_324;
  assign popcount43_r54b_core_326 = popcount43_r54b_core_168 ^ popcount43_r54b_core_306;
  assign popcount43_r54b_core_327 = popcount43_r54b_core_168 & popcount43_r54b_core_306;
  assign popcount43_r54b_core_328 = popcount43_r54b_core_326 ^ popcount43_r54b_core_325;
  assign popcount43_r54b_core_329 = popcount43_r54b_core_326 & popcount43_r54b_core_325;
  assign popcount43_r54b_core_330 = popcount43_r54b_core_327 | popcount43_r54b_core_329;
  assign popcount43_r54b_core_331 = popcount43_r54b_core_152 ^ popcount43_r54b_core_308;
  assign popcount43_r54b_core_332 = popcount43_r54b_core_152 & popcount43_r54b_core_308;
  assign popcount43_r54b_core_333 = popcount43_r54b_core_331 ^ popcount43_r54b_core_330;
  assign popcount43_r54b_core_334 = popcount43_r54b_core_331 & popcount43_r54b_core_330;
  assign popcount43_r54b_core_335 = popcount43_r54b_core_332 | popcount43_r54b_core_334;
  assign popcount43_r54b_core_337 = popcount43_r54b_core_174 & input_a[22];

  assign popcount43_r54b_out[0] = popcount43_r54b_core_314;
  assign popcount43_r54b_out[1] = popcount43_r54b_core_318;
  assign popcount43_r54b_out[2] = popcount43_r54b_core_323;
  assign popcount43_r54b_out[3] = popcount43_r54b_core_328;
  assign popcount43_r54b_out[4] = popcount43_r54b_core_333;
  assign popcount43_r54b_out[5] = popcount43_r54b_core_335;
endmodule