// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.32517
// WCE=17.0
// EP=0.920002%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_g3eh(input [28:0] input_a, output [4:0] popcount29_g3eh_out);
  wire popcount29_g3eh_core_031;
  wire popcount29_g3eh_core_033;
  wire popcount29_g3eh_core_034;
  wire popcount29_g3eh_core_035;
  wire popcount29_g3eh_core_036;
  wire popcount29_g3eh_core_037;
  wire popcount29_g3eh_core_038;
  wire popcount29_g3eh_core_040;
  wire popcount29_g3eh_core_041;
  wire popcount29_g3eh_core_042;
  wire popcount29_g3eh_core_045;
  wire popcount29_g3eh_core_046;
  wire popcount29_g3eh_core_048;
  wire popcount29_g3eh_core_052;
  wire popcount29_g3eh_core_053;
  wire popcount29_g3eh_core_056;
  wire popcount29_g3eh_core_057;
  wire popcount29_g3eh_core_063;
  wire popcount29_g3eh_core_064;
  wire popcount29_g3eh_core_065;
  wire popcount29_g3eh_core_067;
  wire popcount29_g3eh_core_071_not;
  wire popcount29_g3eh_core_072;
  wire popcount29_g3eh_core_074;
  wire popcount29_g3eh_core_075;
  wire popcount29_g3eh_core_078;
  wire popcount29_g3eh_core_079;
  wire popcount29_g3eh_core_080;
  wire popcount29_g3eh_core_084;
  wire popcount29_g3eh_core_086;
  wire popcount29_g3eh_core_090;
  wire popcount29_g3eh_core_091;
  wire popcount29_g3eh_core_093;
  wire popcount29_g3eh_core_095;
  wire popcount29_g3eh_core_097;
  wire popcount29_g3eh_core_100;
  wire popcount29_g3eh_core_101;
  wire popcount29_g3eh_core_102;
  wire popcount29_g3eh_core_104;
  wire popcount29_g3eh_core_105;
  wire popcount29_g3eh_core_106;
  wire popcount29_g3eh_core_107;
  wire popcount29_g3eh_core_110;
  wire popcount29_g3eh_core_115;
  wire popcount29_g3eh_core_119;
  wire popcount29_g3eh_core_122;
  wire popcount29_g3eh_core_123;
  wire popcount29_g3eh_core_126;
  wire popcount29_g3eh_core_128;
  wire popcount29_g3eh_core_129;
  wire popcount29_g3eh_core_131;
  wire popcount29_g3eh_core_132;
  wire popcount29_g3eh_core_134;
  wire popcount29_g3eh_core_136;
  wire popcount29_g3eh_core_138;
  wire popcount29_g3eh_core_141;
  wire popcount29_g3eh_core_143;
  wire popcount29_g3eh_core_144;
  wire popcount29_g3eh_core_145;
  wire popcount29_g3eh_core_147;
  wire popcount29_g3eh_core_149;
  wire popcount29_g3eh_core_150;
  wire popcount29_g3eh_core_151;
  wire popcount29_g3eh_core_153;
  wire popcount29_g3eh_core_154;
  wire popcount29_g3eh_core_155_not;
  wire popcount29_g3eh_core_156;
  wire popcount29_g3eh_core_157_not;
  wire popcount29_g3eh_core_158;
  wire popcount29_g3eh_core_159;
  wire popcount29_g3eh_core_160;
  wire popcount29_g3eh_core_162;
  wire popcount29_g3eh_core_163;
  wire popcount29_g3eh_core_165;
  wire popcount29_g3eh_core_166;
  wire popcount29_g3eh_core_168;
  wire popcount29_g3eh_core_169;
  wire popcount29_g3eh_core_171;
  wire popcount29_g3eh_core_172;
  wire popcount29_g3eh_core_173;
  wire popcount29_g3eh_core_175;
  wire popcount29_g3eh_core_176;
  wire popcount29_g3eh_core_177;
  wire popcount29_g3eh_core_178;
  wire popcount29_g3eh_core_185;
  wire popcount29_g3eh_core_189;
  wire popcount29_g3eh_core_190;
  wire popcount29_g3eh_core_191;
  wire popcount29_g3eh_core_192;
  wire popcount29_g3eh_core_195;
  wire popcount29_g3eh_core_196;
  wire popcount29_g3eh_core_197;
  wire popcount29_g3eh_core_199;
  wire popcount29_g3eh_core_200;
  wire popcount29_g3eh_core_202;
  wire popcount29_g3eh_core_203;
  wire popcount29_g3eh_core_204;
  wire popcount29_g3eh_core_205;
  wire popcount29_g3eh_core_207;

  assign popcount29_g3eh_core_031 = input_a[1] | input_a[3];
  assign popcount29_g3eh_core_033 = ~(input_a[17] & input_a[10]);
  assign popcount29_g3eh_core_034 = input_a[7] & input_a[0];
  assign popcount29_g3eh_core_035 = ~(input_a[10] | input_a[20]);
  assign popcount29_g3eh_core_036 = input_a[1] | input_a[13];
  assign popcount29_g3eh_core_037 = input_a[0] & input_a[23];
  assign popcount29_g3eh_core_038 = input_a[27] ^ input_a[22];
  assign popcount29_g3eh_core_040 = input_a[17] ^ input_a[15];
  assign popcount29_g3eh_core_041 = ~(input_a[9] ^ input_a[14]);
  assign popcount29_g3eh_core_042 = input_a[3] & input_a[4];
  assign popcount29_g3eh_core_045 = ~input_a[26];
  assign popcount29_g3eh_core_046 = ~(input_a[27] | input_a[7]);
  assign popcount29_g3eh_core_048 = input_a[28] | input_a[21];
  assign popcount29_g3eh_core_052 = ~input_a[2];
  assign popcount29_g3eh_core_053 = input_a[26] | input_a[7];
  assign popcount29_g3eh_core_056 = input_a[27] & input_a[18];
  assign popcount29_g3eh_core_057 = ~(input_a[19] ^ input_a[3]);
  assign popcount29_g3eh_core_063 = ~(input_a[22] & input_a[8]);
  assign popcount29_g3eh_core_064 = input_a[18] & input_a[26];
  assign popcount29_g3eh_core_065 = input_a[2] ^ input_a[8];
  assign popcount29_g3eh_core_067 = ~input_a[3];
  assign popcount29_g3eh_core_071_not = ~input_a[11];
  assign popcount29_g3eh_core_072 = input_a[20] & input_a[28];
  assign popcount29_g3eh_core_074 = ~(input_a[23] | input_a[13]);
  assign popcount29_g3eh_core_075 = input_a[15] & input_a[9];
  assign popcount29_g3eh_core_078 = input_a[14] | input_a[12];
  assign popcount29_g3eh_core_079 = input_a[6] & input_a[10];
  assign popcount29_g3eh_core_080 = input_a[0] ^ input_a[11];
  assign popcount29_g3eh_core_084 = input_a[6] ^ input_a[8];
  assign popcount29_g3eh_core_086 = ~(input_a[20] | input_a[19]);
  assign popcount29_g3eh_core_090 = input_a[6] & input_a[18];
  assign popcount29_g3eh_core_091 = ~input_a[11];
  assign popcount29_g3eh_core_093 = ~input_a[9];
  assign popcount29_g3eh_core_095 = ~(input_a[0] & input_a[26]);
  assign popcount29_g3eh_core_097 = ~input_a[27];
  assign popcount29_g3eh_core_100 = input_a[23] & input_a[5];
  assign popcount29_g3eh_core_101 = ~(input_a[16] | input_a[24]);
  assign popcount29_g3eh_core_102 = ~(input_a[6] | input_a[18]);
  assign popcount29_g3eh_core_104 = input_a[10] | input_a[14];
  assign popcount29_g3eh_core_105 = ~(input_a[19] | input_a[15]);
  assign popcount29_g3eh_core_106 = input_a[3] & input_a[19];
  assign popcount29_g3eh_core_107 = ~input_a[12];
  assign popcount29_g3eh_core_110 = ~(input_a[21] ^ input_a[16]);
  assign popcount29_g3eh_core_115 = ~input_a[8];
  assign popcount29_g3eh_core_119 = ~(input_a[15] ^ input_a[14]);
  assign popcount29_g3eh_core_122 = ~(input_a[7] ^ input_a[18]);
  assign popcount29_g3eh_core_123 = ~(input_a[21] & input_a[18]);
  assign popcount29_g3eh_core_126 = ~(input_a[21] ^ input_a[10]);
  assign popcount29_g3eh_core_128 = input_a[7] ^ input_a[20];
  assign popcount29_g3eh_core_129 = ~(input_a[0] & input_a[8]);
  assign popcount29_g3eh_core_131 = input_a[23] ^ input_a[11];
  assign popcount29_g3eh_core_132 = ~(input_a[14] | input_a[9]);
  assign popcount29_g3eh_core_134 = ~(input_a[20] ^ input_a[21]);
  assign popcount29_g3eh_core_136 = input_a[17] & input_a[27];
  assign popcount29_g3eh_core_138 = ~(input_a[24] ^ input_a[11]);
  assign popcount29_g3eh_core_141 = ~(input_a[5] & input_a[7]);
  assign popcount29_g3eh_core_143 = ~input_a[2];
  assign popcount29_g3eh_core_144 = input_a[17] & input_a[12];
  assign popcount29_g3eh_core_145 = ~(input_a[20] & input_a[25]);
  assign popcount29_g3eh_core_147 = input_a[10] & input_a[11];
  assign popcount29_g3eh_core_149 = input_a[5] & input_a[4];
  assign popcount29_g3eh_core_150 = ~(input_a[19] | input_a[26]);
  assign popcount29_g3eh_core_151 = ~(input_a[16] ^ input_a[10]);
  assign popcount29_g3eh_core_153 = input_a[13] | input_a[9];
  assign popcount29_g3eh_core_154 = input_a[12] | input_a[9];
  assign popcount29_g3eh_core_155_not = ~input_a[10];
  assign popcount29_g3eh_core_156 = input_a[11] & input_a[12];
  assign popcount29_g3eh_core_157_not = ~input_a[18];
  assign popcount29_g3eh_core_158 = ~input_a[26];
  assign popcount29_g3eh_core_159 = input_a[2] ^ input_a[11];
  assign popcount29_g3eh_core_160 = ~(input_a[7] | input_a[3]);
  assign popcount29_g3eh_core_162 = ~input_a[15];
  assign popcount29_g3eh_core_163 = ~(input_a[16] | input_a[4]);
  assign popcount29_g3eh_core_165 = ~(input_a[10] & input_a[27]);
  assign popcount29_g3eh_core_166 = ~(input_a[3] & input_a[12]);
  assign popcount29_g3eh_core_168 = ~input_a[26];
  assign popcount29_g3eh_core_169 = ~(input_a[8] ^ input_a[6]);
  assign popcount29_g3eh_core_171 = input_a[22] | input_a[7];
  assign popcount29_g3eh_core_172 = ~(input_a[3] ^ input_a[10]);
  assign popcount29_g3eh_core_173 = ~(input_a[12] & input_a[27]);
  assign popcount29_g3eh_core_175 = input_a[12] & input_a[26];
  assign popcount29_g3eh_core_176 = input_a[3] & input_a[13];
  assign popcount29_g3eh_core_177 = ~input_a[0];
  assign popcount29_g3eh_core_178 = ~(input_a[24] | input_a[24]);
  assign popcount29_g3eh_core_185 = input_a[27] & input_a[23];
  assign popcount29_g3eh_core_189 = ~(input_a[11] ^ input_a[3]);
  assign popcount29_g3eh_core_190 = ~input_a[22];
  assign popcount29_g3eh_core_191 = input_a[16] ^ input_a[22];
  assign popcount29_g3eh_core_192 = input_a[27] ^ input_a[23];
  assign popcount29_g3eh_core_195 = ~input_a[3];
  assign popcount29_g3eh_core_196 = ~(input_a[20] ^ input_a[4]);
  assign popcount29_g3eh_core_197 = input_a[10] ^ input_a[0];
  assign popcount29_g3eh_core_199 = ~(input_a[0] ^ input_a[6]);
  assign popcount29_g3eh_core_200 = ~(input_a[22] & input_a[22]);
  assign popcount29_g3eh_core_202 = ~(input_a[12] ^ input_a[27]);
  assign popcount29_g3eh_core_203 = input_a[16] | input_a[22];
  assign popcount29_g3eh_core_204 = ~(input_a[0] | input_a[2]);
  assign popcount29_g3eh_core_205 = ~(input_a[12] & input_a[0]);
  assign popcount29_g3eh_core_207 = ~input_a[18];

  assign popcount29_g3eh_out[0] = input_a[22];
  assign popcount29_g3eh_out[1] = input_a[3];
  assign popcount29_g3eh_out[2] = 1'b0;
  assign popcount29_g3eh_out[3] = 1'b0;
  assign popcount29_g3eh_out[4] = 1'b1;
endmodule