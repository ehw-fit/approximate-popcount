// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=0.5
// WCE=1.0
// EP=0.5%
// Printed PDK parameters:
//  Area=1619360.0
//  Delay=5217426.0
//  Power=64244.0

module popcount04_zpp2(input [3:0] input_a, output [2:0] popcount04_zpp2_out);
  wire popcount04_zpp2_core_006;
  wire popcount04_zpp2_core_008;
  wire popcount04_zpp2_core_009;
  wire popcount04_zpp2_core_011;
  wire popcount04_zpp2_core_012;
  wire popcount04_zpp2_core_013;
  wire popcount04_zpp2_core_014;
  wire popcount04_zpp2_core_016;

  assign popcount04_zpp2_core_006 = input_a[1] | input_a[3];
  assign popcount04_zpp2_core_008 = ~input_a[0];
  assign popcount04_zpp2_core_009 = input_a[2] & input_a[3];
  assign popcount04_zpp2_core_011 = input_a[3] & popcount04_zpp2_core_008;
  assign popcount04_zpp2_core_012 = input_a[3] ^ input_a[2];
  assign popcount04_zpp2_core_013 = input_a[0] & popcount04_zpp2_core_009;
  assign popcount04_zpp2_core_014 = popcount04_zpp2_core_012 | popcount04_zpp2_core_011;
  assign popcount04_zpp2_core_016 = input_a[0] ^ input_a[0];

  assign popcount04_zpp2_out[0] = input_a[1];
  assign popcount04_zpp2_out[1] = popcount04_zpp2_core_014;
  assign popcount04_zpp2_out[2] = popcount04_zpp2_core_013;
endmodule