// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.12099
// WCE=24.0
// EP=0.928801%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_k4qz(input [31:0] input_a, output [5:0] popcount32_k4qz_out);
  wire popcount32_k4qz_core_034;
  wire popcount32_k4qz_core_035;
  wire popcount32_k4qz_core_036;
  wire popcount32_k4qz_core_037;
  wire popcount32_k4qz_core_038;
  wire popcount32_k4qz_core_039;
  wire popcount32_k4qz_core_040;
  wire popcount32_k4qz_core_043;
  wire popcount32_k4qz_core_044;
  wire popcount32_k4qz_core_046;
  wire popcount32_k4qz_core_047;
  wire popcount32_k4qz_core_048;
  wire popcount32_k4qz_core_049;
  wire popcount32_k4qz_core_051;
  wire popcount32_k4qz_core_052;
  wire popcount32_k4qz_core_055;
  wire popcount32_k4qz_core_056;
  wire popcount32_k4qz_core_058;
  wire popcount32_k4qz_core_061;
  wire popcount32_k4qz_core_063;
  wire popcount32_k4qz_core_065;
  wire popcount32_k4qz_core_068;
  wire popcount32_k4qz_core_069;
  wire popcount32_k4qz_core_071;
  wire popcount32_k4qz_core_072;
  wire popcount32_k4qz_core_073;
  wire popcount32_k4qz_core_077;
  wire popcount32_k4qz_core_078;
  wire popcount32_k4qz_core_080_not;
  wire popcount32_k4qz_core_082;
  wire popcount32_k4qz_core_083;
  wire popcount32_k4qz_core_087;
  wire popcount32_k4qz_core_088;
  wire popcount32_k4qz_core_089;
  wire popcount32_k4qz_core_091;
  wire popcount32_k4qz_core_092;
  wire popcount32_k4qz_core_093;
  wire popcount32_k4qz_core_094;
  wire popcount32_k4qz_core_096;
  wire popcount32_k4qz_core_098;
  wire popcount32_k4qz_core_099;
  wire popcount32_k4qz_core_100;
  wire popcount32_k4qz_core_101;
  wire popcount32_k4qz_core_103;
  wire popcount32_k4qz_core_107;
  wire popcount32_k4qz_core_111;
  wire popcount32_k4qz_core_115;
  wire popcount32_k4qz_core_116;
  wire popcount32_k4qz_core_120;
  wire popcount32_k4qz_core_122;
  wire popcount32_k4qz_core_123_not;
  wire popcount32_k4qz_core_126;
  wire popcount32_k4qz_core_128_not;
  wire popcount32_k4qz_core_130;
  wire popcount32_k4qz_core_131;
  wire popcount32_k4qz_core_132;
  wire popcount32_k4qz_core_136_not;
  wire popcount32_k4qz_core_137;
  wire popcount32_k4qz_core_138;
  wire popcount32_k4qz_core_139;
  wire popcount32_k4qz_core_140;
  wire popcount32_k4qz_core_141;
  wire popcount32_k4qz_core_144;
  wire popcount32_k4qz_core_145;
  wire popcount32_k4qz_core_146;
  wire popcount32_k4qz_core_147;
  wire popcount32_k4qz_core_148;
  wire popcount32_k4qz_core_149;
  wire popcount32_k4qz_core_150;
  wire popcount32_k4qz_core_151;
  wire popcount32_k4qz_core_152;
  wire popcount32_k4qz_core_153;
  wire popcount32_k4qz_core_154;
  wire popcount32_k4qz_core_155;
  wire popcount32_k4qz_core_158;
  wire popcount32_k4qz_core_160;
  wire popcount32_k4qz_core_161;
  wire popcount32_k4qz_core_162;
  wire popcount32_k4qz_core_163;
  wire popcount32_k4qz_core_165;
  wire popcount32_k4qz_core_166;
  wire popcount32_k4qz_core_167;
  wire popcount32_k4qz_core_168;
  wire popcount32_k4qz_core_169;
  wire popcount32_k4qz_core_170;
  wire popcount32_k4qz_core_171;
  wire popcount32_k4qz_core_172;
  wire popcount32_k4qz_core_173;
  wire popcount32_k4qz_core_175;
  wire popcount32_k4qz_core_176;
  wire popcount32_k4qz_core_177;
  wire popcount32_k4qz_core_179;
  wire popcount32_k4qz_core_182;
  wire popcount32_k4qz_core_184;
  wire popcount32_k4qz_core_186_not;
  wire popcount32_k4qz_core_188;
  wire popcount32_k4qz_core_191;
  wire popcount32_k4qz_core_192;
  wire popcount32_k4qz_core_193;
  wire popcount32_k4qz_core_194;
  wire popcount32_k4qz_core_195;
  wire popcount32_k4qz_core_196;
  wire popcount32_k4qz_core_198;
  wire popcount32_k4qz_core_200;
  wire popcount32_k4qz_core_201;
  wire popcount32_k4qz_core_203;
  wire popcount32_k4qz_core_205;
  wire popcount32_k4qz_core_209;
  wire popcount32_k4qz_core_211;
  wire popcount32_k4qz_core_212;
  wire popcount32_k4qz_core_214;
  wire popcount32_k4qz_core_218;
  wire popcount32_k4qz_core_219;
  wire popcount32_k4qz_core_221;
  wire popcount32_k4qz_core_222;
  wire popcount32_k4qz_core_223;
  wire popcount32_k4qz_core_224;
  wire popcount32_k4qz_core_225;

  assign popcount32_k4qz_core_034 = ~(input_a[8] | input_a[10]);
  assign popcount32_k4qz_core_035 = input_a[16] & input_a[7];
  assign popcount32_k4qz_core_036 = ~input_a[19];
  assign popcount32_k4qz_core_037 = ~input_a[18];
  assign popcount32_k4qz_core_038 = input_a[22] | input_a[31];
  assign popcount32_k4qz_core_039 = input_a[11] ^ input_a[26];
  assign popcount32_k4qz_core_040 = ~input_a[21];
  assign popcount32_k4qz_core_043 = ~(input_a[22] ^ input_a[14]);
  assign popcount32_k4qz_core_044 = ~(input_a[16] & input_a[10]);
  assign popcount32_k4qz_core_046 = ~(input_a[13] ^ input_a[11]);
  assign popcount32_k4qz_core_047 = ~input_a[15];
  assign popcount32_k4qz_core_048 = input_a[18] | input_a[5];
  assign popcount32_k4qz_core_049 = ~(input_a[29] ^ input_a[26]);
  assign popcount32_k4qz_core_051 = ~(input_a[14] | input_a[13]);
  assign popcount32_k4qz_core_052 = ~input_a[30];
  assign popcount32_k4qz_core_055 = input_a[28] ^ input_a[18];
  assign popcount32_k4qz_core_056 = input_a[2] ^ input_a[5];
  assign popcount32_k4qz_core_058 = input_a[14] ^ input_a[10];
  assign popcount32_k4qz_core_061 = input_a[19] | input_a[7];
  assign popcount32_k4qz_core_063 = ~(input_a[14] ^ input_a[27]);
  assign popcount32_k4qz_core_065 = ~(input_a[6] & input_a[25]);
  assign popcount32_k4qz_core_068 = ~input_a[25];
  assign popcount32_k4qz_core_069 = input_a[23] | input_a[9];
  assign popcount32_k4qz_core_071 = input_a[4] & input_a[23];
  assign popcount32_k4qz_core_072 = ~input_a[31];
  assign popcount32_k4qz_core_073 = input_a[7] & input_a[19];
  assign popcount32_k4qz_core_077 = ~(input_a[11] & input_a[25]);
  assign popcount32_k4qz_core_078 = input_a[21] ^ input_a[16];
  assign popcount32_k4qz_core_080_not = ~input_a[1];
  assign popcount32_k4qz_core_082 = ~input_a[30];
  assign popcount32_k4qz_core_083 = input_a[12] ^ input_a[2];
  assign popcount32_k4qz_core_087 = input_a[16] ^ input_a[2];
  assign popcount32_k4qz_core_088 = input_a[10] ^ input_a[9];
  assign popcount32_k4qz_core_089 = ~(input_a[1] | input_a[9]);
  assign popcount32_k4qz_core_091 = ~(input_a[15] | input_a[6]);
  assign popcount32_k4qz_core_092 = input_a[13] | input_a[7];
  assign popcount32_k4qz_core_093 = ~(input_a[9] ^ input_a[18]);
  assign popcount32_k4qz_core_094 = ~input_a[28];
  assign popcount32_k4qz_core_096 = input_a[23] & input_a[17];
  assign popcount32_k4qz_core_098 = input_a[16] ^ input_a[18];
  assign popcount32_k4qz_core_099 = ~input_a[18];
  assign popcount32_k4qz_core_100 = ~(input_a[4] | input_a[13]);
  assign popcount32_k4qz_core_101 = ~(input_a[30] ^ input_a[26]);
  assign popcount32_k4qz_core_103 = ~(input_a[0] & input_a[26]);
  assign popcount32_k4qz_core_107 = ~input_a[0];
  assign popcount32_k4qz_core_111 = input_a[26] ^ input_a[5];
  assign popcount32_k4qz_core_115 = input_a[2] & input_a[8];
  assign popcount32_k4qz_core_116 = ~(input_a[13] ^ input_a[6]);
  assign popcount32_k4qz_core_120 = input_a[1] | input_a[17];
  assign popcount32_k4qz_core_122 = ~(input_a[0] & input_a[28]);
  assign popcount32_k4qz_core_123_not = ~input_a[22];
  assign popcount32_k4qz_core_126 = ~(input_a[19] ^ input_a[13]);
  assign popcount32_k4qz_core_128_not = ~input_a[18];
  assign popcount32_k4qz_core_130 = ~(input_a[26] | input_a[14]);
  assign popcount32_k4qz_core_131 = input_a[1] | input_a[25];
  assign popcount32_k4qz_core_132 = ~(input_a[21] & input_a[24]);
  assign popcount32_k4qz_core_136_not = ~input_a[28];
  assign popcount32_k4qz_core_137 = ~(input_a[6] ^ input_a[24]);
  assign popcount32_k4qz_core_138 = ~(input_a[14] | input_a[0]);
  assign popcount32_k4qz_core_139 = input_a[8] ^ input_a[22];
  assign popcount32_k4qz_core_140 = ~(input_a[19] & input_a[8]);
  assign popcount32_k4qz_core_141 = input_a[30] | input_a[22];
  assign popcount32_k4qz_core_144 = input_a[9] | input_a[18];
  assign popcount32_k4qz_core_145 = ~(input_a[26] ^ input_a[4]);
  assign popcount32_k4qz_core_146 = input_a[21] | input_a[18];
  assign popcount32_k4qz_core_147 = input_a[23] ^ input_a[27];
  assign popcount32_k4qz_core_148 = ~input_a[28];
  assign popcount32_k4qz_core_149 = input_a[1] ^ input_a[29];
  assign popcount32_k4qz_core_150 = ~(input_a[3] & input_a[7]);
  assign popcount32_k4qz_core_151 = ~input_a[17];
  assign popcount32_k4qz_core_152 = ~(input_a[9] ^ input_a[8]);
  assign popcount32_k4qz_core_153 = ~(input_a[21] ^ input_a[8]);
  assign popcount32_k4qz_core_154 = input_a[31] & input_a[7];
  assign popcount32_k4qz_core_155 = ~(input_a[10] ^ input_a[27]);
  assign popcount32_k4qz_core_158 = ~(input_a[20] ^ input_a[21]);
  assign popcount32_k4qz_core_160 = ~(input_a[14] ^ input_a[5]);
  assign popcount32_k4qz_core_161 = ~input_a[30];
  assign popcount32_k4qz_core_162 = input_a[23] & input_a[14];
  assign popcount32_k4qz_core_163 = input_a[26] ^ input_a[21];
  assign popcount32_k4qz_core_165 = input_a[23] | input_a[6];
  assign popcount32_k4qz_core_166 = ~(input_a[5] | input_a[0]);
  assign popcount32_k4qz_core_167 = input_a[3] ^ input_a[28];
  assign popcount32_k4qz_core_168 = input_a[30] ^ input_a[19];
  assign popcount32_k4qz_core_169 = input_a[4] & input_a[17];
  assign popcount32_k4qz_core_170 = ~(input_a[28] ^ input_a[2]);
  assign popcount32_k4qz_core_171 = ~(input_a[29] | input_a[2]);
  assign popcount32_k4qz_core_172 = ~(input_a[6] ^ input_a[15]);
  assign popcount32_k4qz_core_173 = input_a[4] ^ input_a[26];
  assign popcount32_k4qz_core_175 = input_a[20] | input_a[9];
  assign popcount32_k4qz_core_176 = input_a[19] ^ input_a[14];
  assign popcount32_k4qz_core_177 = ~(input_a[6] | input_a[28]);
  assign popcount32_k4qz_core_179 = input_a[10] | input_a[29];
  assign popcount32_k4qz_core_182 = ~(input_a[5] | input_a[15]);
  assign popcount32_k4qz_core_184 = input_a[16] ^ input_a[19];
  assign popcount32_k4qz_core_186_not = ~input_a[0];
  assign popcount32_k4qz_core_188 = ~(input_a[6] | input_a[20]);
  assign popcount32_k4qz_core_191 = ~(input_a[15] ^ input_a[14]);
  assign popcount32_k4qz_core_192 = ~(input_a[23] ^ input_a[8]);
  assign popcount32_k4qz_core_193 = ~(input_a[2] ^ input_a[23]);
  assign popcount32_k4qz_core_194 = input_a[1] & input_a[2];
  assign popcount32_k4qz_core_195 = ~input_a[19];
  assign popcount32_k4qz_core_196 = input_a[31] & input_a[8];
  assign popcount32_k4qz_core_198 = input_a[31] & input_a[28];
  assign popcount32_k4qz_core_200 = input_a[10] ^ input_a[31];
  assign popcount32_k4qz_core_201 = ~(input_a[6] ^ input_a[23]);
  assign popcount32_k4qz_core_203 = ~input_a[5];
  assign popcount32_k4qz_core_205 = ~(input_a[3] | input_a[27]);
  assign popcount32_k4qz_core_209 = ~(input_a[10] ^ input_a[22]);
  assign popcount32_k4qz_core_211 = input_a[20] ^ input_a[20];
  assign popcount32_k4qz_core_212 = ~(input_a[20] | input_a[1]);
  assign popcount32_k4qz_core_214 = ~(input_a[21] ^ input_a[25]);
  assign popcount32_k4qz_core_218 = ~input_a[2];
  assign popcount32_k4qz_core_219 = ~input_a[27];
  assign popcount32_k4qz_core_221 = input_a[13] ^ input_a[5];
  assign popcount32_k4qz_core_222 = ~(input_a[12] | input_a[12]);
  assign popcount32_k4qz_core_223 = ~(input_a[22] | input_a[3]);
  assign popcount32_k4qz_core_224 = ~(input_a[23] ^ input_a[11]);
  assign popcount32_k4qz_core_225 = ~input_a[22];

  assign popcount32_k4qz_out[0] = 1'b0;
  assign popcount32_k4qz_out[1] = 1'b0;
  assign popcount32_k4qz_out[2] = 1'b0;
  assign popcount32_k4qz_out[3] = 1'b1;
  assign popcount32_k4qz_out[4] = 1'b1;
  assign popcount32_k4qz_out[5] = 1'b0;
endmodule