// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.25671
// WCE=4.0
// EP=0.766312%
// Printed PDK parameters:
//  Area=111667772.0
//  Delay=91282784.0
//  Power=5080200.0

module popcount36_n5a1(input [35:0] input_a, output [5:0] popcount36_n5a1_out);
  wire popcount36_n5a1_core_038;
  wire popcount36_n5a1_core_039;
  wire popcount36_n5a1_core_040;
  wire popcount36_n5a1_core_041;
  wire popcount36_n5a1_core_042;
  wire popcount36_n5a1_core_043;
  wire popcount36_n5a1_core_044;
  wire popcount36_n5a1_core_045;
  wire popcount36_n5a1_core_046;
  wire popcount36_n5a1_core_049;
  wire popcount36_n5a1_core_050;
  wire popcount36_n5a1_core_051;
  wire popcount36_n5a1_core_052;
  wire popcount36_n5a1_core_053;
  wire popcount36_n5a1_core_054;
  wire popcount36_n5a1_core_055;
  wire popcount36_n5a1_core_057;
  wire popcount36_n5a1_core_058;
  wire popcount36_n5a1_core_059;
  wire popcount36_n5a1_core_060;
  wire popcount36_n5a1_core_061;
  wire popcount36_n5a1_core_062;
  wire popcount36_n5a1_core_063;
  wire popcount36_n5a1_core_066;
  wire popcount36_n5a1_core_068;
  wire popcount36_n5a1_core_069;
  wire popcount36_n5a1_core_070;
  wire popcount36_n5a1_core_071;
  wire popcount36_n5a1_core_072;
  wire popcount36_n5a1_core_073;
  wire popcount36_n5a1_core_074;
  wire popcount36_n5a1_core_075;
  wire popcount36_n5a1_core_076;
  wire popcount36_n5a1_core_077;
  wire popcount36_n5a1_core_079;
  wire popcount36_n5a1_core_080;
  wire popcount36_n5a1_core_081;
  wire popcount36_n5a1_core_082;
  wire popcount36_n5a1_core_083;
  wire popcount36_n5a1_core_084;
  wire popcount36_n5a1_core_085;
  wire popcount36_n5a1_core_086;
  wire popcount36_n5a1_core_087;
  wire popcount36_n5a1_core_088;
  wire popcount36_n5a1_core_089;
  wire popcount36_n5a1_core_091;
  wire popcount36_n5a1_core_092;
  wire popcount36_n5a1_core_093;
  wire popcount36_n5a1_core_094;
  wire popcount36_n5a1_core_095;
  wire popcount36_n5a1_core_096;
  wire popcount36_n5a1_core_097;
  wire popcount36_n5a1_core_099;
  wire popcount36_n5a1_core_100;
  wire popcount36_n5a1_core_101;
  wire popcount36_n5a1_core_102;
  wire popcount36_n5a1_core_103;
  wire popcount36_n5a1_core_104;
  wire popcount36_n5a1_core_105;
  wire popcount36_n5a1_core_108;
  wire popcount36_n5a1_core_109;
  wire popcount36_n5a1_core_110;
  wire popcount36_n5a1_core_111;
  wire popcount36_n5a1_core_112;
  wire popcount36_n5a1_core_113;
  wire popcount36_n5a1_core_114;
  wire popcount36_n5a1_core_115;
  wire popcount36_n5a1_core_116;
  wire popcount36_n5a1_core_117;
  wire popcount36_n5a1_core_118;
  wire popcount36_n5a1_core_119;
  wire popcount36_n5a1_core_122;
  wire popcount36_n5a1_core_123;
  wire popcount36_n5a1_core_124;
  wire popcount36_n5a1_core_125;
  wire popcount36_n5a1_core_126;
  wire popcount36_n5a1_core_127;
  wire popcount36_n5a1_core_128;
  wire popcount36_n5a1_core_129;
  wire popcount36_n5a1_core_130;
  wire popcount36_n5a1_core_131;
  wire popcount36_n5a1_core_132;
  wire popcount36_n5a1_core_133;
  wire popcount36_n5a1_core_134;
  wire popcount36_n5a1_core_135;
  wire popcount36_n5a1_core_136;
  wire popcount36_n5a1_core_137;
  wire popcount36_n5a1_core_138;
  wire popcount36_n5a1_core_140;
  wire popcount36_n5a1_core_142;
  wire popcount36_n5a1_core_143;
  wire popcount36_n5a1_core_144;
  wire popcount36_n5a1_core_145;
  wire popcount36_n5a1_core_146;
  wire popcount36_n5a1_core_147;
  wire popcount36_n5a1_core_148;
  wire popcount36_n5a1_core_149;
  wire popcount36_n5a1_core_150;
  wire popcount36_n5a1_core_151;
  wire popcount36_n5a1_core_152;
  wire popcount36_n5a1_core_155;
  wire popcount36_n5a1_core_156;
  wire popcount36_n5a1_core_157;
  wire popcount36_n5a1_core_158;
  wire popcount36_n5a1_core_159;
  wire popcount36_n5a1_core_160;
  wire popcount36_n5a1_core_163;
  wire popcount36_n5a1_core_164;
  wire popcount36_n5a1_core_165;
  wire popcount36_n5a1_core_166;
  wire popcount36_n5a1_core_167;
  wire popcount36_n5a1_core_172;
  wire popcount36_n5a1_core_173;
  wire popcount36_n5a1_core_174;
  wire popcount36_n5a1_core_175;
  wire popcount36_n5a1_core_176;
  wire popcount36_n5a1_core_177;
  wire popcount36_n5a1_core_178;
  wire popcount36_n5a1_core_179;
  wire popcount36_n5a1_core_180;
  wire popcount36_n5a1_core_181;
  wire popcount36_n5a1_core_182;
  wire popcount36_n5a1_core_186;
  wire popcount36_n5a1_core_187;
  wire popcount36_n5a1_core_188;
  wire popcount36_n5a1_core_189;
  wire popcount36_n5a1_core_191;
  wire popcount36_n5a1_core_192;
  wire popcount36_n5a1_core_193;
  wire popcount36_n5a1_core_194;
  wire popcount36_n5a1_core_195;
  wire popcount36_n5a1_core_197;
  wire popcount36_n5a1_core_199;
  wire popcount36_n5a1_core_200;
  wire popcount36_n5a1_core_201;
  wire popcount36_n5a1_core_202;
  wire popcount36_n5a1_core_203;
  wire popcount36_n5a1_core_205;
  wire popcount36_n5a1_core_206;
  wire popcount36_n5a1_core_207;
  wire popcount36_n5a1_core_208;
  wire popcount36_n5a1_core_209;
  wire popcount36_n5a1_core_210;
  wire popcount36_n5a1_core_211;
  wire popcount36_n5a1_core_214;
  wire popcount36_n5a1_core_216;
  wire popcount36_n5a1_core_217;
  wire popcount36_n5a1_core_218;
  wire popcount36_n5a1_core_219;
  wire popcount36_n5a1_core_220;
  wire popcount36_n5a1_core_221;
  wire popcount36_n5a1_core_222;
  wire popcount36_n5a1_core_223;
  wire popcount36_n5a1_core_224;
  wire popcount36_n5a1_core_225;
  wire popcount36_n5a1_core_227;
  wire popcount36_n5a1_core_230;
  wire popcount36_n5a1_core_231;
  wire popcount36_n5a1_core_232;
  wire popcount36_n5a1_core_233;
  wire popcount36_n5a1_core_235;
  wire popcount36_n5a1_core_236;
  wire popcount36_n5a1_core_237;
  wire popcount36_n5a1_core_238;
  wire popcount36_n5a1_core_239;
  wire popcount36_n5a1_core_240;
  wire popcount36_n5a1_core_241;
  wire popcount36_n5a1_core_242;
  wire popcount36_n5a1_core_243;
  wire popcount36_n5a1_core_244;
  wire popcount36_n5a1_core_248;
  wire popcount36_n5a1_core_249;
  wire popcount36_n5a1_core_250;
  wire popcount36_n5a1_core_251;
  wire popcount36_n5a1_core_254;
  wire popcount36_n5a1_core_255;
  wire popcount36_n5a1_core_257;
  wire popcount36_n5a1_core_258;
  wire popcount36_n5a1_core_259;
  wire popcount36_n5a1_core_260;
  wire popcount36_n5a1_core_261;
  wire popcount36_n5a1_core_262;
  wire popcount36_n5a1_core_263;
  wire popcount36_n5a1_core_264;
  wire popcount36_n5a1_core_265;
  wire popcount36_n5a1_core_266;
  wire popcount36_n5a1_core_267;
  wire popcount36_n5a1_core_268;
  wire popcount36_n5a1_core_269;
  wire popcount36_n5a1_core_270;
  wire popcount36_n5a1_core_271;
  wire popcount36_n5a1_core_273;
  wire popcount36_n5a1_core_276;

  assign popcount36_n5a1_core_038 = input_a[0] ^ input_a[1];
  assign popcount36_n5a1_core_039 = input_a[0] & input_a[1];
  assign popcount36_n5a1_core_040 = input_a[2] ^ input_a[3];
  assign popcount36_n5a1_core_041 = input_a[2] & input_a[3];
  assign popcount36_n5a1_core_042 = popcount36_n5a1_core_038 ^ popcount36_n5a1_core_040;
  assign popcount36_n5a1_core_043 = popcount36_n5a1_core_038 & popcount36_n5a1_core_040;
  assign popcount36_n5a1_core_044 = popcount36_n5a1_core_039 ^ popcount36_n5a1_core_041;
  assign popcount36_n5a1_core_045 = popcount36_n5a1_core_039 & popcount36_n5a1_core_041;
  assign popcount36_n5a1_core_046 = popcount36_n5a1_core_044 | popcount36_n5a1_core_043;
  assign popcount36_n5a1_core_049 = ~(input_a[13] & input_a[9]);
  assign popcount36_n5a1_core_050 = input_a[4] & input_a[5];
  assign popcount36_n5a1_core_051 = input_a[7] ^ input_a[8];
  assign popcount36_n5a1_core_052 = input_a[7] & input_a[8];
  assign popcount36_n5a1_core_053 = input_a[6] ^ popcount36_n5a1_core_051;
  assign popcount36_n5a1_core_054 = input_a[6] & popcount36_n5a1_core_051;
  assign popcount36_n5a1_core_055 = popcount36_n5a1_core_052 | popcount36_n5a1_core_054;
  assign popcount36_n5a1_core_057 = ~(input_a[18] ^ input_a[5]);
  assign popcount36_n5a1_core_058 = input_a[32] & popcount36_n5a1_core_053;
  assign popcount36_n5a1_core_059 = popcount36_n5a1_core_050 ^ popcount36_n5a1_core_055;
  assign popcount36_n5a1_core_060 = popcount36_n5a1_core_050 & popcount36_n5a1_core_055;
  assign popcount36_n5a1_core_061 = popcount36_n5a1_core_059 ^ popcount36_n5a1_core_058;
  assign popcount36_n5a1_core_062 = popcount36_n5a1_core_059 & popcount36_n5a1_core_058;
  assign popcount36_n5a1_core_063 = popcount36_n5a1_core_060 | popcount36_n5a1_core_062;
  assign popcount36_n5a1_core_066 = ~popcount36_n5a1_core_042;
  assign popcount36_n5a1_core_068 = popcount36_n5a1_core_046 ^ popcount36_n5a1_core_061;
  assign popcount36_n5a1_core_069 = popcount36_n5a1_core_046 & popcount36_n5a1_core_061;
  assign popcount36_n5a1_core_070 = popcount36_n5a1_core_068 ^ popcount36_n5a1_core_042;
  assign popcount36_n5a1_core_071 = popcount36_n5a1_core_068 & popcount36_n5a1_core_042;
  assign popcount36_n5a1_core_072 = popcount36_n5a1_core_069 | popcount36_n5a1_core_071;
  assign popcount36_n5a1_core_073 = popcount36_n5a1_core_045 ^ popcount36_n5a1_core_063;
  assign popcount36_n5a1_core_074 = popcount36_n5a1_core_045 & popcount36_n5a1_core_063;
  assign popcount36_n5a1_core_075 = popcount36_n5a1_core_073 ^ popcount36_n5a1_core_072;
  assign popcount36_n5a1_core_076 = popcount36_n5a1_core_073 & popcount36_n5a1_core_072;
  assign popcount36_n5a1_core_077 = popcount36_n5a1_core_074 | popcount36_n5a1_core_076;
  assign popcount36_n5a1_core_079 = input_a[17] ^ input_a[5];
  assign popcount36_n5a1_core_080 = ~(input_a[9] & input_a[10]);
  assign popcount36_n5a1_core_081 = input_a[9] & input_a[10];
  assign popcount36_n5a1_core_082 = input_a[11] ^ input_a[12];
  assign popcount36_n5a1_core_083 = input_a[11] & input_a[12];
  assign popcount36_n5a1_core_084 = ~(popcount36_n5a1_core_080 & popcount36_n5a1_core_082);
  assign popcount36_n5a1_core_085 = popcount36_n5a1_core_080 & popcount36_n5a1_core_082;
  assign popcount36_n5a1_core_086 = popcount36_n5a1_core_081 ^ popcount36_n5a1_core_083;
  assign popcount36_n5a1_core_087 = popcount36_n5a1_core_081 & popcount36_n5a1_core_083;
  assign popcount36_n5a1_core_088 = popcount36_n5a1_core_086 | popcount36_n5a1_core_085;
  assign popcount36_n5a1_core_089 = ~input_a[29];
  assign popcount36_n5a1_core_091 = input_a[13] ^ input_a[14];
  assign popcount36_n5a1_core_092 = input_a[13] & input_a[14];
  assign popcount36_n5a1_core_093 = input_a[16] ^ input_a[17];
  assign popcount36_n5a1_core_094 = input_a[16] & input_a[17];
  assign popcount36_n5a1_core_095 = input_a[15] ^ popcount36_n5a1_core_093;
  assign popcount36_n5a1_core_096 = input_a[15] & popcount36_n5a1_core_093;
  assign popcount36_n5a1_core_097 = popcount36_n5a1_core_094 | popcount36_n5a1_core_096;
  assign popcount36_n5a1_core_099 = popcount36_n5a1_core_091 ^ popcount36_n5a1_core_095;
  assign popcount36_n5a1_core_100 = popcount36_n5a1_core_091 & popcount36_n5a1_core_095;
  assign popcount36_n5a1_core_101 = popcount36_n5a1_core_092 ^ popcount36_n5a1_core_097;
  assign popcount36_n5a1_core_102 = popcount36_n5a1_core_092 & popcount36_n5a1_core_097;
  assign popcount36_n5a1_core_103 = popcount36_n5a1_core_101 ^ popcount36_n5a1_core_100;
  assign popcount36_n5a1_core_104 = popcount36_n5a1_core_101 & popcount36_n5a1_core_100;
  assign popcount36_n5a1_core_105 = popcount36_n5a1_core_102 | popcount36_n5a1_core_104;
  assign popcount36_n5a1_core_108 = popcount36_n5a1_core_084 ^ popcount36_n5a1_core_099;
  assign popcount36_n5a1_core_109 = popcount36_n5a1_core_084 & popcount36_n5a1_core_099;
  assign popcount36_n5a1_core_110 = popcount36_n5a1_core_088 ^ popcount36_n5a1_core_103;
  assign popcount36_n5a1_core_111 = popcount36_n5a1_core_088 & popcount36_n5a1_core_103;
  assign popcount36_n5a1_core_112 = popcount36_n5a1_core_110 ^ popcount36_n5a1_core_109;
  assign popcount36_n5a1_core_113 = popcount36_n5a1_core_110 & popcount36_n5a1_core_109;
  assign popcount36_n5a1_core_114 = popcount36_n5a1_core_111 | popcount36_n5a1_core_113;
  assign popcount36_n5a1_core_115 = popcount36_n5a1_core_087 ^ popcount36_n5a1_core_105;
  assign popcount36_n5a1_core_116 = popcount36_n5a1_core_087 & popcount36_n5a1_core_105;
  assign popcount36_n5a1_core_117 = popcount36_n5a1_core_115 ^ popcount36_n5a1_core_114;
  assign popcount36_n5a1_core_118 = popcount36_n5a1_core_115 & popcount36_n5a1_core_114;
  assign popcount36_n5a1_core_119 = popcount36_n5a1_core_116 | popcount36_n5a1_core_118;
  assign popcount36_n5a1_core_122 = popcount36_n5a1_core_066 ^ popcount36_n5a1_core_108;
  assign popcount36_n5a1_core_123 = popcount36_n5a1_core_066 & popcount36_n5a1_core_108;
  assign popcount36_n5a1_core_124 = popcount36_n5a1_core_070 ^ popcount36_n5a1_core_112;
  assign popcount36_n5a1_core_125 = popcount36_n5a1_core_070 & popcount36_n5a1_core_112;
  assign popcount36_n5a1_core_126 = popcount36_n5a1_core_124 ^ popcount36_n5a1_core_123;
  assign popcount36_n5a1_core_127 = popcount36_n5a1_core_124 & popcount36_n5a1_core_123;
  assign popcount36_n5a1_core_128 = popcount36_n5a1_core_125 | popcount36_n5a1_core_127;
  assign popcount36_n5a1_core_129 = popcount36_n5a1_core_075 ^ popcount36_n5a1_core_117;
  assign popcount36_n5a1_core_130 = popcount36_n5a1_core_075 & popcount36_n5a1_core_117;
  assign popcount36_n5a1_core_131 = popcount36_n5a1_core_129 ^ popcount36_n5a1_core_128;
  assign popcount36_n5a1_core_132 = popcount36_n5a1_core_129 & popcount36_n5a1_core_128;
  assign popcount36_n5a1_core_133 = popcount36_n5a1_core_130 | popcount36_n5a1_core_132;
  assign popcount36_n5a1_core_134 = popcount36_n5a1_core_077 ^ popcount36_n5a1_core_119;
  assign popcount36_n5a1_core_135 = popcount36_n5a1_core_077 & popcount36_n5a1_core_119;
  assign popcount36_n5a1_core_136 = popcount36_n5a1_core_134 ^ popcount36_n5a1_core_133;
  assign popcount36_n5a1_core_137 = popcount36_n5a1_core_134 & popcount36_n5a1_core_133;
  assign popcount36_n5a1_core_138 = popcount36_n5a1_core_135 | popcount36_n5a1_core_137;
  assign popcount36_n5a1_core_140 = input_a[18] & input_a[7];
  assign popcount36_n5a1_core_142 = ~(input_a[31] | input_a[14]);
  assign popcount36_n5a1_core_143 = ~input_a[33];
  assign popcount36_n5a1_core_144 = input_a[18] ^ input_a[19];
  assign popcount36_n5a1_core_145 = input_a[18] & input_a[19];
  assign popcount36_n5a1_core_146 = input_a[20] ^ input_a[21];
  assign popcount36_n5a1_core_147 = input_a[20] & input_a[21];
  assign popcount36_n5a1_core_148 = popcount36_n5a1_core_144 ^ popcount36_n5a1_core_146;
  assign popcount36_n5a1_core_149 = popcount36_n5a1_core_144 & popcount36_n5a1_core_146;
  assign popcount36_n5a1_core_150 = popcount36_n5a1_core_145 ^ popcount36_n5a1_core_147;
  assign popcount36_n5a1_core_151 = popcount36_n5a1_core_145 & popcount36_n5a1_core_147;
  assign popcount36_n5a1_core_152 = popcount36_n5a1_core_150 | popcount36_n5a1_core_149;
  assign popcount36_n5a1_core_155 = input_a[22] ^ input_a[23];
  assign popcount36_n5a1_core_156 = input_a[22] & input_a[23];
  assign popcount36_n5a1_core_157 = ~(input_a[25] & input_a[26]);
  assign popcount36_n5a1_core_158 = input_a[25] & input_a[26];
  assign popcount36_n5a1_core_159 = input_a[24] & popcount36_n5a1_core_157;
  assign popcount36_n5a1_core_160 = input_a[21] ^ input_a[4];
  assign popcount36_n5a1_core_163 = popcount36_n5a1_core_155 ^ popcount36_n5a1_core_159;
  assign popcount36_n5a1_core_164 = popcount36_n5a1_core_155 & input_a[24];
  assign popcount36_n5a1_core_165 = popcount36_n5a1_core_156 ^ popcount36_n5a1_core_158;
  assign popcount36_n5a1_core_166 = popcount36_n5a1_core_156 & popcount36_n5a1_core_158;
  assign popcount36_n5a1_core_167 = popcount36_n5a1_core_165 | popcount36_n5a1_core_164;
  assign popcount36_n5a1_core_172 = popcount36_n5a1_core_148 ^ popcount36_n5a1_core_163;
  assign popcount36_n5a1_core_173 = popcount36_n5a1_core_148 & popcount36_n5a1_core_163;
  assign popcount36_n5a1_core_174 = popcount36_n5a1_core_152 ^ popcount36_n5a1_core_167;
  assign popcount36_n5a1_core_175 = popcount36_n5a1_core_152 & popcount36_n5a1_core_167;
  assign popcount36_n5a1_core_176 = popcount36_n5a1_core_174 ^ popcount36_n5a1_core_173;
  assign popcount36_n5a1_core_177 = popcount36_n5a1_core_174 & popcount36_n5a1_core_173;
  assign popcount36_n5a1_core_178 = popcount36_n5a1_core_175 | popcount36_n5a1_core_177;
  assign popcount36_n5a1_core_179 = popcount36_n5a1_core_151 ^ popcount36_n5a1_core_166;
  assign popcount36_n5a1_core_180 = popcount36_n5a1_core_151 & popcount36_n5a1_core_166;
  assign popcount36_n5a1_core_181 = popcount36_n5a1_core_179 | popcount36_n5a1_core_178;
  assign popcount36_n5a1_core_182 = ~(input_a[22] | input_a[7]);
  assign popcount36_n5a1_core_186 = input_a[27] ^ input_a[28];
  assign popcount36_n5a1_core_187 = input_a[27] & input_a[28];
  assign popcount36_n5a1_core_188 = input_a[29] | input_a[30];
  assign popcount36_n5a1_core_189 = input_a[29] & input_a[30];
  assign popcount36_n5a1_core_191 = popcount36_n5a1_core_186 & popcount36_n5a1_core_188;
  assign popcount36_n5a1_core_192 = popcount36_n5a1_core_187 ^ popcount36_n5a1_core_189;
  assign popcount36_n5a1_core_193 = popcount36_n5a1_core_187 & popcount36_n5a1_core_189;
  assign popcount36_n5a1_core_194 = popcount36_n5a1_core_192 | popcount36_n5a1_core_191;
  assign popcount36_n5a1_core_195 = ~(input_a[32] ^ input_a[20]);
  assign popcount36_n5a1_core_197 = ~input_a[31];
  assign popcount36_n5a1_core_199 = input_a[34] ^ input_a[35];
  assign popcount36_n5a1_core_200 = input_a[34] & input_a[35];
  assign popcount36_n5a1_core_201 = input_a[33] ^ popcount36_n5a1_core_199;
  assign popcount36_n5a1_core_202 = input_a[33] & popcount36_n5a1_core_199;
  assign popcount36_n5a1_core_203 = popcount36_n5a1_core_200 | popcount36_n5a1_core_202;
  assign popcount36_n5a1_core_205 = popcount36_n5a1_core_197 ^ popcount36_n5a1_core_201;
  assign popcount36_n5a1_core_206 = popcount36_n5a1_core_197 & popcount36_n5a1_core_201;
  assign popcount36_n5a1_core_207 = input_a[31] ^ popcount36_n5a1_core_203;
  assign popcount36_n5a1_core_208 = input_a[31] & popcount36_n5a1_core_203;
  assign popcount36_n5a1_core_209 = popcount36_n5a1_core_207 ^ popcount36_n5a1_core_206;
  assign popcount36_n5a1_core_210 = popcount36_n5a1_core_207 & popcount36_n5a1_core_206;
  assign popcount36_n5a1_core_211 = popcount36_n5a1_core_208 | popcount36_n5a1_core_210;
  assign popcount36_n5a1_core_214 = ~input_a[16];
  assign popcount36_n5a1_core_216 = popcount36_n5a1_core_194 ^ popcount36_n5a1_core_209;
  assign popcount36_n5a1_core_217 = popcount36_n5a1_core_194 & popcount36_n5a1_core_209;
  assign popcount36_n5a1_core_218 = popcount36_n5a1_core_216 ^ popcount36_n5a1_core_205;
  assign popcount36_n5a1_core_219 = popcount36_n5a1_core_216 & popcount36_n5a1_core_205;
  assign popcount36_n5a1_core_220 = popcount36_n5a1_core_217 | popcount36_n5a1_core_219;
  assign popcount36_n5a1_core_221 = popcount36_n5a1_core_193 ^ popcount36_n5a1_core_211;
  assign popcount36_n5a1_core_222 = popcount36_n5a1_core_193 & popcount36_n5a1_core_211;
  assign popcount36_n5a1_core_223 = popcount36_n5a1_core_221 ^ popcount36_n5a1_core_220;
  assign popcount36_n5a1_core_224 = popcount36_n5a1_core_221 & popcount36_n5a1_core_220;
  assign popcount36_n5a1_core_225 = popcount36_n5a1_core_222 | popcount36_n5a1_core_224;
  assign popcount36_n5a1_core_227 = input_a[18] & input_a[1];
  assign popcount36_n5a1_core_230 = input_a[20] & input_a[2];
  assign popcount36_n5a1_core_231 = popcount36_n5a1_core_176 & popcount36_n5a1_core_218;
  assign popcount36_n5a1_core_232 = input_a[17] ^ input_a[28];
  assign popcount36_n5a1_core_233 = ~(input_a[32] | input_a[23]);
  assign popcount36_n5a1_core_235 = popcount36_n5a1_core_181 ^ popcount36_n5a1_core_223;
  assign popcount36_n5a1_core_236 = popcount36_n5a1_core_181 & popcount36_n5a1_core_223;
  assign popcount36_n5a1_core_237 = popcount36_n5a1_core_235 ^ popcount36_n5a1_core_231;
  assign popcount36_n5a1_core_238 = popcount36_n5a1_core_235 & popcount36_n5a1_core_231;
  assign popcount36_n5a1_core_239 = popcount36_n5a1_core_236 | popcount36_n5a1_core_238;
  assign popcount36_n5a1_core_240 = popcount36_n5a1_core_180 ^ popcount36_n5a1_core_225;
  assign popcount36_n5a1_core_241 = popcount36_n5a1_core_180 & popcount36_n5a1_core_225;
  assign popcount36_n5a1_core_242 = popcount36_n5a1_core_240 ^ popcount36_n5a1_core_239;
  assign popcount36_n5a1_core_243 = popcount36_n5a1_core_240 & popcount36_n5a1_core_239;
  assign popcount36_n5a1_core_244 = popcount36_n5a1_core_241 | popcount36_n5a1_core_243;
  assign popcount36_n5a1_core_248 = input_a[4] & input_a[32];
  assign popcount36_n5a1_core_249 = input_a[27] & input_a[20];
  assign popcount36_n5a1_core_250 = popcount36_n5a1_core_122 ^ popcount36_n5a1_core_172;
  assign popcount36_n5a1_core_251 = popcount36_n5a1_core_122 & popcount36_n5a1_core_172;
  assign popcount36_n5a1_core_254 = popcount36_n5a1_core_126 ^ popcount36_n5a1_core_251;
  assign popcount36_n5a1_core_255 = popcount36_n5a1_core_126 & popcount36_n5a1_core_251;
  assign popcount36_n5a1_core_257 = popcount36_n5a1_core_131 ^ popcount36_n5a1_core_237;
  assign popcount36_n5a1_core_258 = popcount36_n5a1_core_131 & popcount36_n5a1_core_237;
  assign popcount36_n5a1_core_259 = popcount36_n5a1_core_257 ^ popcount36_n5a1_core_255;
  assign popcount36_n5a1_core_260 = popcount36_n5a1_core_257 & popcount36_n5a1_core_255;
  assign popcount36_n5a1_core_261 = popcount36_n5a1_core_258 | popcount36_n5a1_core_260;
  assign popcount36_n5a1_core_262 = popcount36_n5a1_core_136 ^ popcount36_n5a1_core_242;
  assign popcount36_n5a1_core_263 = popcount36_n5a1_core_136 & popcount36_n5a1_core_242;
  assign popcount36_n5a1_core_264 = popcount36_n5a1_core_262 ^ popcount36_n5a1_core_261;
  assign popcount36_n5a1_core_265 = popcount36_n5a1_core_262 & popcount36_n5a1_core_261;
  assign popcount36_n5a1_core_266 = popcount36_n5a1_core_263 | popcount36_n5a1_core_265;
  assign popcount36_n5a1_core_267 = popcount36_n5a1_core_138 ^ popcount36_n5a1_core_244;
  assign popcount36_n5a1_core_268 = popcount36_n5a1_core_138 & popcount36_n5a1_core_244;
  assign popcount36_n5a1_core_269 = popcount36_n5a1_core_267 ^ popcount36_n5a1_core_266;
  assign popcount36_n5a1_core_270 = popcount36_n5a1_core_267 & popcount36_n5a1_core_266;
  assign popcount36_n5a1_core_271 = popcount36_n5a1_core_268 | popcount36_n5a1_core_270;
  assign popcount36_n5a1_core_273 = input_a[32] | input_a[12];
  assign popcount36_n5a1_core_276 = ~(input_a[28] | input_a[8]);

  assign popcount36_n5a1_out[0] = popcount36_n5a1_core_250;
  assign popcount36_n5a1_out[1] = popcount36_n5a1_core_254;
  assign popcount36_n5a1_out[2] = popcount36_n5a1_core_259;
  assign popcount36_n5a1_out[3] = popcount36_n5a1_core_264;
  assign popcount36_n5a1_out[4] = popcount36_n5a1_core_269;
  assign popcount36_n5a1_out[5] = popcount36_n5a1_core_271;
endmodule