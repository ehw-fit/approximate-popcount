// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.84434
// WCE=19.0
// EP=0.890559%
// Printed PDK parameters:
//  Area=14922358.0
//  Delay=44415928.0
//  Power=526180.0

module popcount38_z7t9(input [37:0] input_a, output [5:0] popcount38_z7t9_out);
  wire popcount38_z7t9_core_041;
  wire popcount38_z7t9_core_042;
  wire popcount38_z7t9_core_045;
  wire popcount38_z7t9_core_046;
  wire popcount38_z7t9_core_047;
  wire popcount38_z7t9_core_048;
  wire popcount38_z7t9_core_049;
  wire popcount38_z7t9_core_050;
  wire popcount38_z7t9_core_051;
  wire popcount38_z7t9_core_052;
  wire popcount38_z7t9_core_056;
  wire popcount38_z7t9_core_057;
  wire popcount38_z7t9_core_058;
  wire popcount38_z7t9_core_059;
  wire popcount38_z7t9_core_060;
  wire popcount38_z7t9_core_061;
  wire popcount38_z7t9_core_064;
  wire popcount38_z7t9_core_067;
  wire popcount38_z7t9_core_068;
  wire popcount38_z7t9_core_069;
  wire popcount38_z7t9_core_070;
  wire popcount38_z7t9_core_071;
  wire popcount38_z7t9_core_072;
  wire popcount38_z7t9_core_074;
  wire popcount38_z7t9_core_076;
  wire popcount38_z7t9_core_078;
  wire popcount38_z7t9_core_079;
  wire popcount38_z7t9_core_080;
  wire popcount38_z7t9_core_081;
  wire popcount38_z7t9_core_082;
  wire popcount38_z7t9_core_083;
  wire popcount38_z7t9_core_084;
  wire popcount38_z7t9_core_085;
  wire popcount38_z7t9_core_086;
  wire popcount38_z7t9_core_087;
  wire popcount38_z7t9_core_088;
  wire popcount38_z7t9_core_091;
  wire popcount38_z7t9_core_092;
  wire popcount38_z7t9_core_093;
  wire popcount38_z7t9_core_094;
  wire popcount38_z7t9_core_095;
  wire popcount38_z7t9_core_096;
  wire popcount38_z7t9_core_097_not;
  wire popcount38_z7t9_core_098;
  wire popcount38_z7t9_core_099;
  wire popcount38_z7t9_core_100;
  wire popcount38_z7t9_core_101;
  wire popcount38_z7t9_core_104;
  wire popcount38_z7t9_core_107;
  wire popcount38_z7t9_core_110;
  wire popcount38_z7t9_core_111;
  wire popcount38_z7t9_core_112;
  wire popcount38_z7t9_core_113;
  wire popcount38_z7t9_core_114;
  wire popcount38_z7t9_core_117;
  wire popcount38_z7t9_core_118;
  wire popcount38_z7t9_core_121;
  wire popcount38_z7t9_core_122;
  wire popcount38_z7t9_core_124;
  wire popcount38_z7t9_core_125;
  wire popcount38_z7t9_core_126;
  wire popcount38_z7t9_core_127;
  wire popcount38_z7t9_core_130;
  wire popcount38_z7t9_core_131;
  wire popcount38_z7t9_core_133;
  wire popcount38_z7t9_core_134;
  wire popcount38_z7t9_core_135;
  wire popcount38_z7t9_core_137;
  wire popcount38_z7t9_core_138;
  wire popcount38_z7t9_core_139;
  wire popcount38_z7t9_core_142;
  wire popcount38_z7t9_core_143;
  wire popcount38_z7t9_core_145;
  wire popcount38_z7t9_core_147;
  wire popcount38_z7t9_core_148;
  wire popcount38_z7t9_core_153;
  wire popcount38_z7t9_core_154;
  wire popcount38_z7t9_core_156;
  wire popcount38_z7t9_core_157;
  wire popcount38_z7t9_core_159;
  wire popcount38_z7t9_core_160;
  wire popcount38_z7t9_core_161;
  wire popcount38_z7t9_core_164_not;
  wire popcount38_z7t9_core_165;
  wire popcount38_z7t9_core_167;
  wire popcount38_z7t9_core_168;
  wire popcount38_z7t9_core_171;
  wire popcount38_z7t9_core_172;
  wire popcount38_z7t9_core_173;
  wire popcount38_z7t9_core_174;
  wire popcount38_z7t9_core_175;
  wire popcount38_z7t9_core_177;
  wire popcount38_z7t9_core_178;
  wire popcount38_z7t9_core_179;
  wire popcount38_z7t9_core_181;
  wire popcount38_z7t9_core_182;
  wire popcount38_z7t9_core_186;
  wire popcount38_z7t9_core_187_not;
  wire popcount38_z7t9_core_189;
  wire popcount38_z7t9_core_190;
  wire popcount38_z7t9_core_195;
  wire popcount38_z7t9_core_199;
  wire popcount38_z7t9_core_200;
  wire popcount38_z7t9_core_201;
  wire popcount38_z7t9_core_204;
  wire popcount38_z7t9_core_205_not;
  wire popcount38_z7t9_core_210;
  wire popcount38_z7t9_core_211;
  wire popcount38_z7t9_core_212;
  wire popcount38_z7t9_core_215;
  wire popcount38_z7t9_core_218;
  wire popcount38_z7t9_core_219;
  wire popcount38_z7t9_core_221;
  wire popcount38_z7t9_core_222;
  wire popcount38_z7t9_core_223;
  wire popcount38_z7t9_core_224;
  wire popcount38_z7t9_core_225;
  wire popcount38_z7t9_core_226;
  wire popcount38_z7t9_core_228;
  wire popcount38_z7t9_core_229;
  wire popcount38_z7t9_core_230;
  wire popcount38_z7t9_core_231;
  wire popcount38_z7t9_core_234;
  wire popcount38_z7t9_core_236;
  wire popcount38_z7t9_core_240;
  wire popcount38_z7t9_core_241;
  wire popcount38_z7t9_core_242;
  wire popcount38_z7t9_core_243;
  wire popcount38_z7t9_core_244;
  wire popcount38_z7t9_core_245;
  wire popcount38_z7t9_core_246;
  wire popcount38_z7t9_core_248;
  wire popcount38_z7t9_core_249;
  wire popcount38_z7t9_core_250;
  wire popcount38_z7t9_core_252;
  wire popcount38_z7t9_core_255;
  wire popcount38_z7t9_core_258;
  wire popcount38_z7t9_core_260;
  wire popcount38_z7t9_core_261;
  wire popcount38_z7t9_core_263;
  wire popcount38_z7t9_core_264;
  wire popcount38_z7t9_core_267;
  wire popcount38_z7t9_core_269;
  wire popcount38_z7t9_core_270;
  wire popcount38_z7t9_core_273;
  wire popcount38_z7t9_core_274;
  wire popcount38_z7t9_core_275;
  wire popcount38_z7t9_core_276;
  wire popcount38_z7t9_core_277;
  wire popcount38_z7t9_core_279;
  wire popcount38_z7t9_core_280;
  wire popcount38_z7t9_core_281;
  wire popcount38_z7t9_core_284;
  wire popcount38_z7t9_core_285;
  wire popcount38_z7t9_core_289;
  wire popcount38_z7t9_core_291;
  wire popcount38_z7t9_core_292;
  wire popcount38_z7t9_core_293;
  wire popcount38_z7t9_core_294;

  assign popcount38_z7t9_core_041 = ~input_a[24];
  assign popcount38_z7t9_core_042 = ~(input_a[6] | input_a[28]);
  assign popcount38_z7t9_core_045 = ~(input_a[8] | input_a[18]);
  assign popcount38_z7t9_core_046 = input_a[27] ^ input_a[16];
  assign popcount38_z7t9_core_047 = ~input_a[34];
  assign popcount38_z7t9_core_048 = ~input_a[20];
  assign popcount38_z7t9_core_049 = ~(input_a[20] & input_a[18]);
  assign popcount38_z7t9_core_050 = input_a[15] & input_a[34];
  assign popcount38_z7t9_core_051 = ~(input_a[14] & input_a[34]);
  assign popcount38_z7t9_core_052 = ~(input_a[1] & input_a[37]);
  assign popcount38_z7t9_core_056 = input_a[27] ^ input_a[9];
  assign popcount38_z7t9_core_057 = input_a[31] ^ input_a[1];
  assign popcount38_z7t9_core_058 = input_a[0] | input_a[37];
  assign popcount38_z7t9_core_059 = input_a[13] | input_a[28];
  assign popcount38_z7t9_core_060 = input_a[6] ^ input_a[28];
  assign popcount38_z7t9_core_061 = input_a[7] ^ input_a[0];
  assign popcount38_z7t9_core_064 = ~input_a[3];
  assign popcount38_z7t9_core_067 = input_a[27] | input_a[20];
  assign popcount38_z7t9_core_068 = ~(input_a[10] ^ input_a[16]);
  assign popcount38_z7t9_core_069 = ~input_a[36];
  assign popcount38_z7t9_core_070 = input_a[37] ^ input_a[35];
  assign popcount38_z7t9_core_071 = ~input_a[20];
  assign popcount38_z7t9_core_072 = input_a[34] & input_a[12];
  assign popcount38_z7t9_core_074 = ~input_a[30];
  assign popcount38_z7t9_core_076 = ~input_a[16];
  assign popcount38_z7t9_core_078 = input_a[30] & input_a[22];
  assign popcount38_z7t9_core_079 = input_a[16] & input_a[17];
  assign popcount38_z7t9_core_080 = ~(input_a[27] & input_a[15]);
  assign popcount38_z7t9_core_081 = ~(input_a[27] & input_a[3]);
  assign popcount38_z7t9_core_082 = input_a[36] | input_a[21];
  assign popcount38_z7t9_core_083 = input_a[21] & input_a[20];
  assign popcount38_z7t9_core_084 = input_a[29] & input_a[8];
  assign popcount38_z7t9_core_085 = input_a[32] ^ input_a[22];
  assign popcount38_z7t9_core_086 = ~(input_a[26] ^ input_a[3]);
  assign popcount38_z7t9_core_087 = input_a[27] & input_a[11];
  assign popcount38_z7t9_core_088 = input_a[16] | input_a[29];
  assign popcount38_z7t9_core_091 = input_a[25] & input_a[5];
  assign popcount38_z7t9_core_092 = popcount38_z7t9_core_083 ^ popcount38_z7t9_core_088;
  assign popcount38_z7t9_core_093 = popcount38_z7t9_core_083 & popcount38_z7t9_core_088;
  assign popcount38_z7t9_core_094 = popcount38_z7t9_core_092 ^ popcount38_z7t9_core_091;
  assign popcount38_z7t9_core_095 = input_a[23] & popcount38_z7t9_core_091;
  assign popcount38_z7t9_core_096 = popcount38_z7t9_core_093 | popcount38_z7t9_core_095;
  assign popcount38_z7t9_core_097_not = ~popcount38_z7t9_core_096;
  assign popcount38_z7t9_core_098 = input_a[21] & input_a[20];
  assign popcount38_z7t9_core_099 = input_a[11] | input_a[5];
  assign popcount38_z7t9_core_100 = ~(input_a[8] ^ input_a[30]);
  assign popcount38_z7t9_core_101 = input_a[4] & input_a[27];
  assign popcount38_z7t9_core_104 = ~input_a[13];
  assign popcount38_z7t9_core_107 = ~(input_a[19] | input_a[24]);
  assign popcount38_z7t9_core_110 = ~(input_a[0] | input_a[12]);
  assign popcount38_z7t9_core_111 = ~(input_a[28] & input_a[2]);
  assign popcount38_z7t9_core_112 = input_a[11] & input_a[31];
  assign popcount38_z7t9_core_113 = ~(input_a[1] & input_a[14]);
  assign popcount38_z7t9_core_114 = ~(input_a[25] ^ input_a[26]);
  assign popcount38_z7t9_core_117 = input_a[31] ^ input_a[0];
  assign popcount38_z7t9_core_118 = ~(input_a[25] & input_a[25]);
  assign popcount38_z7t9_core_121 = input_a[11] & input_a[31];
  assign popcount38_z7t9_core_122 = popcount38_z7t9_core_094 | popcount38_z7t9_core_121;
  assign popcount38_z7t9_core_124 = ~(input_a[9] ^ input_a[19]);
  assign popcount38_z7t9_core_125 = popcount38_z7t9_core_097_not ^ popcount38_z7t9_core_122;
  assign popcount38_z7t9_core_126 = popcount38_z7t9_core_097_not & popcount38_z7t9_core_122;
  assign popcount38_z7t9_core_127 = input_a[29] | popcount38_z7t9_core_126;
  assign popcount38_z7t9_core_130 = popcount38_z7t9_core_098 | popcount38_z7t9_core_127;
  assign popcount38_z7t9_core_131 = ~(input_a[26] | input_a[30]);
  assign popcount38_z7t9_core_133 = input_a[27] & input_a[13];
  assign popcount38_z7t9_core_134 = input_a[35] | input_a[37];
  assign popcount38_z7t9_core_135 = ~(input_a[35] | input_a[33]);
  assign popcount38_z7t9_core_137 = input_a[21] | input_a[18];
  assign popcount38_z7t9_core_138 = ~(input_a[2] & input_a[31]);
  assign popcount38_z7t9_core_139 = ~input_a[2];
  assign popcount38_z7t9_core_142 = popcount38_z7t9_core_125 ^ input_a[23];
  assign popcount38_z7t9_core_143 = popcount38_z7t9_core_125 & input_a[23];
  assign popcount38_z7t9_core_145 = input_a[16] | popcount38_z7t9_core_130;
  assign popcount38_z7t9_core_147 = popcount38_z7t9_core_145 ^ popcount38_z7t9_core_143;
  assign popcount38_z7t9_core_148 = popcount38_z7t9_core_145 & input_a[23];
  assign popcount38_z7t9_core_153 = ~(input_a[27] & input_a[22]);
  assign popcount38_z7t9_core_154 = input_a[22] & input_a[17];
  assign popcount38_z7t9_core_156 = input_a[22] & input_a[21];
  assign popcount38_z7t9_core_157 = input_a[9] & input_a[37];
  assign popcount38_z7t9_core_159 = input_a[9] | input_a[17];
  assign popcount38_z7t9_core_160 = ~(input_a[30] ^ input_a[9]);
  assign popcount38_z7t9_core_161 = ~(input_a[21] ^ input_a[12]);
  assign popcount38_z7t9_core_164_not = ~input_a[10];
  assign popcount38_z7t9_core_165 = ~(input_a[14] & input_a[10]);
  assign popcount38_z7t9_core_167 = input_a[5] & input_a[29];
  assign popcount38_z7t9_core_168 = input_a[20] | input_a[17];
  assign popcount38_z7t9_core_171 = ~(input_a[25] & input_a[24]);
  assign popcount38_z7t9_core_172 = ~(input_a[35] & input_a[19]);
  assign popcount38_z7t9_core_173 = ~(input_a[8] & input_a[36]);
  assign popcount38_z7t9_core_174 = input_a[17] & input_a[16];
  assign popcount38_z7t9_core_175 = input_a[15] & input_a[11];
  assign popcount38_z7t9_core_177 = input_a[28] | input_a[19];
  assign popcount38_z7t9_core_178 = ~(input_a[35] ^ input_a[2]);
  assign popcount38_z7t9_core_179 = input_a[15] ^ input_a[1];
  assign popcount38_z7t9_core_181 = input_a[28] & input_a[12];
  assign popcount38_z7t9_core_182 = ~(input_a[3] | input_a[10]);
  assign popcount38_z7t9_core_186 = ~input_a[24];
  assign popcount38_z7t9_core_187_not = ~input_a[27];
  assign popcount38_z7t9_core_189 = ~(input_a[1] ^ input_a[20]);
  assign popcount38_z7t9_core_190 = ~(input_a[25] | input_a[0]);
  assign popcount38_z7t9_core_195 = input_a[36] ^ input_a[29];
  assign popcount38_z7t9_core_199 = input_a[30] ^ input_a[23];
  assign popcount38_z7t9_core_200 = ~(input_a[10] ^ input_a[25]);
  assign popcount38_z7t9_core_201 = ~(input_a[6] & input_a[27]);
  assign popcount38_z7t9_core_204 = ~(input_a[32] & input_a[22]);
  assign popcount38_z7t9_core_205_not = ~input_a[1];
  assign popcount38_z7t9_core_210 = ~input_a[7];
  assign popcount38_z7t9_core_211 = input_a[28] & input_a[2];
  assign popcount38_z7t9_core_212 = ~(input_a[28] | input_a[7]);
  assign popcount38_z7t9_core_215 = input_a[24] & input_a[20];
  assign popcount38_z7t9_core_218 = ~input_a[16];
  assign popcount38_z7t9_core_219 = ~(input_a[14] | input_a[37]);
  assign popcount38_z7t9_core_221 = input_a[13] & input_a[8];
  assign popcount38_z7t9_core_222 = ~(input_a[2] & input_a[3]);
  assign popcount38_z7t9_core_223 = input_a[1] ^ input_a[20];
  assign popcount38_z7t9_core_224 = ~(input_a[37] | input_a[19]);
  assign popcount38_z7t9_core_225 = ~(input_a[6] ^ input_a[26]);
  assign popcount38_z7t9_core_226 = input_a[5] ^ input_a[14];
  assign popcount38_z7t9_core_228 = ~(input_a[36] & input_a[2]);
  assign popcount38_z7t9_core_229 = ~(input_a[23] & input_a[17]);
  assign popcount38_z7t9_core_230 = ~(input_a[35] & input_a[20]);
  assign popcount38_z7t9_core_231 = ~(input_a[12] | input_a[8]);
  assign popcount38_z7t9_core_234 = input_a[35] | input_a[7];
  assign popcount38_z7t9_core_236 = ~input_a[13];
  assign popcount38_z7t9_core_240 = ~input_a[30];
  assign popcount38_z7t9_core_241 = ~input_a[26];
  assign popcount38_z7t9_core_242 = ~(input_a[24] & input_a[25]);
  assign popcount38_z7t9_core_243 = ~(input_a[15] | input_a[17]);
  assign popcount38_z7t9_core_244 = ~(input_a[14] & input_a[12]);
  assign popcount38_z7t9_core_245 = ~(input_a[13] ^ input_a[19]);
  assign popcount38_z7t9_core_246 = ~(input_a[22] & input_a[28]);
  assign popcount38_z7t9_core_248 = ~input_a[9];
  assign popcount38_z7t9_core_249 = input_a[18] & input_a[26];
  assign popcount38_z7t9_core_250 = ~(input_a[23] | input_a[22]);
  assign popcount38_z7t9_core_252 = ~(input_a[8] & input_a[16]);
  assign popcount38_z7t9_core_255 = ~input_a[1];
  assign popcount38_z7t9_core_258 = input_a[37] & input_a[33];
  assign popcount38_z7t9_core_260 = ~(input_a[18] | input_a[22]);
  assign popcount38_z7t9_core_261 = ~(input_a[28] ^ input_a[25]);
  assign popcount38_z7t9_core_263 = input_a[22] | input_a[4];
  assign popcount38_z7t9_core_264 = ~(input_a[12] | input_a[0]);
  assign popcount38_z7t9_core_267 = ~input_a[0];
  assign popcount38_z7t9_core_269 = ~(input_a[37] ^ input_a[9]);
  assign popcount38_z7t9_core_270 = input_a[20] | input_a[25];
  assign popcount38_z7t9_core_273 = input_a[11] | input_a[16];
  assign popcount38_z7t9_core_274 = input_a[17] & input_a[22];
  assign popcount38_z7t9_core_275 = ~(input_a[10] | input_a[6]);
  assign popcount38_z7t9_core_276 = input_a[35] | input_a[24];
  assign popcount38_z7t9_core_277 = ~popcount38_z7t9_core_142;
  assign popcount38_z7t9_core_279 = popcount38_z7t9_core_277 ^ popcount38_z7t9_core_276;
  assign popcount38_z7t9_core_280 = popcount38_z7t9_core_277 & popcount38_z7t9_core_276;
  assign popcount38_z7t9_core_281 = popcount38_z7t9_core_142 | popcount38_z7t9_core_280;
  assign popcount38_z7t9_core_284 = popcount38_z7t9_core_147 ^ popcount38_z7t9_core_281;
  assign popcount38_z7t9_core_285 = popcount38_z7t9_core_147 & popcount38_z7t9_core_281;
  assign popcount38_z7t9_core_289 = popcount38_z7t9_core_148 | popcount38_z7t9_core_285;
  assign popcount38_z7t9_core_291 = input_a[20] ^ input_a[4];
  assign popcount38_z7t9_core_292 = ~(input_a[15] ^ input_a[26]);
  assign popcount38_z7t9_core_293 = input_a[3] ^ input_a[4];
  assign popcount38_z7t9_core_294 = ~(input_a[15] ^ input_a[9]);

  assign popcount38_z7t9_out[0] = input_a[37];
  assign popcount38_z7t9_out[1] = 1'b1;
  assign popcount38_z7t9_out[2] = popcount38_z7t9_core_279;
  assign popcount38_z7t9_out[3] = popcount38_z7t9_core_284;
  assign popcount38_z7t9_out[4] = popcount38_z7t9_core_289;
  assign popcount38_z7t9_out[5] = 1'b0;
endmodule