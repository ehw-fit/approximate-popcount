// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.25293
// WCE=14.0
// EP=0.903075%
// Printed PDK parameters:
//  Area=15514901.0
//  Delay=39289576.0
//  Power=685370.0

module popcount28_ykzy(input [27:0] input_a, output [4:0] popcount28_ykzy_out);
  wire popcount28_ykzy_core_030;
  wire popcount28_ykzy_core_031;
  wire popcount28_ykzy_core_032;
  wire popcount28_ykzy_core_040;
  wire popcount28_ykzy_core_041;
  wire popcount28_ykzy_core_043;
  wire popcount28_ykzy_core_044;
  wire popcount28_ykzy_core_046;
  wire popcount28_ykzy_core_047;
  wire popcount28_ykzy_core_048;
  wire popcount28_ykzy_core_049;
  wire popcount28_ykzy_core_050;
  wire popcount28_ykzy_core_051;
  wire popcount28_ykzy_core_052;
  wire popcount28_ykzy_core_055;
  wire popcount28_ykzy_core_056;
  wire popcount28_ykzy_core_059;
  wire popcount28_ykzy_core_060;
  wire popcount28_ykzy_core_062;
  wire popcount28_ykzy_core_063;
  wire popcount28_ykzy_core_065;
  wire popcount28_ykzy_core_067;
  wire popcount28_ykzy_core_069;
  wire popcount28_ykzy_core_072;
  wire popcount28_ykzy_core_073;
  wire popcount28_ykzy_core_074;
  wire popcount28_ykzy_core_077;
  wire popcount28_ykzy_core_078;
  wire popcount28_ykzy_core_079;
  wire popcount28_ykzy_core_080;
  wire popcount28_ykzy_core_082;
  wire popcount28_ykzy_core_083;
  wire popcount28_ykzy_core_084;
  wire popcount28_ykzy_core_085;
  wire popcount28_ykzy_core_086_not;
  wire popcount28_ykzy_core_087;
  wire popcount28_ykzy_core_088;
  wire popcount28_ykzy_core_091;
  wire popcount28_ykzy_core_093;
  wire popcount28_ykzy_core_097;
  wire popcount28_ykzy_core_098;
  wire popcount28_ykzy_core_099;
  wire popcount28_ykzy_core_102;
  wire popcount28_ykzy_core_103;
  wire popcount28_ykzy_core_104;
  wire popcount28_ykzy_core_106;
  wire popcount28_ykzy_core_107;
  wire popcount28_ykzy_core_108;
  wire popcount28_ykzy_core_109;
  wire popcount28_ykzy_core_112;
  wire popcount28_ykzy_core_113;
  wire popcount28_ykzy_core_114;
  wire popcount28_ykzy_core_116;
  wire popcount28_ykzy_core_117;
  wire popcount28_ykzy_core_118;
  wire popcount28_ykzy_core_119;
  wire popcount28_ykzy_core_120;
  wire popcount28_ykzy_core_121;
  wire popcount28_ykzy_core_123;
  wire popcount28_ykzy_core_124;
  wire popcount28_ykzy_core_125;
  wire popcount28_ykzy_core_126;
  wire popcount28_ykzy_core_127;
  wire popcount28_ykzy_core_128;
  wire popcount28_ykzy_core_133;
  wire popcount28_ykzy_core_134;
  wire popcount28_ykzy_core_135;
  wire popcount28_ykzy_core_137;
  wire popcount28_ykzy_core_139;
  wire popcount28_ykzy_core_140;
  wire popcount28_ykzy_core_142;
  wire popcount28_ykzy_core_143;
  wire popcount28_ykzy_core_144;
  wire popcount28_ykzy_core_145;
  wire popcount28_ykzy_core_147;
  wire popcount28_ykzy_core_148;
  wire popcount28_ykzy_core_149;
  wire popcount28_ykzy_core_150;
  wire popcount28_ykzy_core_151;
  wire popcount28_ykzy_core_153;
  wire popcount28_ykzy_core_154;
  wire popcount28_ykzy_core_159;
  wire popcount28_ykzy_core_161;
  wire popcount28_ykzy_core_162;
  wire popcount28_ykzy_core_163;
  wire popcount28_ykzy_core_164;
  wire popcount28_ykzy_core_165;
  wire popcount28_ykzy_core_166;
  wire popcount28_ykzy_core_168;
  wire popcount28_ykzy_core_171;
  wire popcount28_ykzy_core_172;
  wire popcount28_ykzy_core_173;
  wire popcount28_ykzy_core_174;
  wire popcount28_ykzy_core_176;
  wire popcount28_ykzy_core_178;
  wire popcount28_ykzy_core_180;
  wire popcount28_ykzy_core_181;
  wire popcount28_ykzy_core_182_not;
  wire popcount28_ykzy_core_184;
  wire popcount28_ykzy_core_185;
  wire popcount28_ykzy_core_186;
  wire popcount28_ykzy_core_189_not;
  wire popcount28_ykzy_core_192;
  wire popcount28_ykzy_core_193;
  wire popcount28_ykzy_core_194;
  wire popcount28_ykzy_core_195;
  wire popcount28_ykzy_core_196;
  wire popcount28_ykzy_core_198;
  wire popcount28_ykzy_core_201;

  assign popcount28_ykzy_core_030 = input_a[24] | input_a[23];
  assign popcount28_ykzy_core_031 = ~(input_a[27] ^ input_a[2]);
  assign popcount28_ykzy_core_032 = ~(input_a[25] | input_a[9]);
  assign popcount28_ykzy_core_040 = ~input_a[3];
  assign popcount28_ykzy_core_041 = input_a[9] ^ input_a[23];
  assign popcount28_ykzy_core_043 = ~input_a[20];
  assign popcount28_ykzy_core_044 = input_a[5] & input_a[6];
  assign popcount28_ykzy_core_046 = ~(input_a[17] & input_a[24]);
  assign popcount28_ykzy_core_047 = input_a[24] | input_a[8];
  assign popcount28_ykzy_core_048 = ~(input_a[9] | input_a[16]);
  assign popcount28_ykzy_core_049 = input_a[4] ^ input_a[19];
  assign popcount28_ykzy_core_050 = ~input_a[27];
  assign popcount28_ykzy_core_051 = ~input_a[22];
  assign popcount28_ykzy_core_052 = ~(input_a[25] & input_a[17]);
  assign popcount28_ykzy_core_055 = input_a[3] ^ input_a[8];
  assign popcount28_ykzy_core_056 = ~(input_a[13] ^ input_a[26]);
  assign popcount28_ykzy_core_059 = ~(input_a[19] | input_a[21]);
  assign popcount28_ykzy_core_060 = ~(input_a[16] | input_a[18]);
  assign popcount28_ykzy_core_062 = ~(input_a[27] & input_a[25]);
  assign popcount28_ykzy_core_063 = ~(input_a[22] & input_a[4]);
  assign popcount28_ykzy_core_065 = ~(input_a[16] & input_a[10]);
  assign popcount28_ykzy_core_067 = input_a[2] ^ input_a[15];
  assign popcount28_ykzy_core_069 = ~input_a[22];
  assign popcount28_ykzy_core_072 = ~input_a[7];
  assign popcount28_ykzy_core_073 = input_a[22] ^ input_a[22];
  assign popcount28_ykzy_core_074 = ~(input_a[3] | input_a[5]);
  assign popcount28_ykzy_core_077 = input_a[5] & input_a[21];
  assign popcount28_ykzy_core_078 = ~(input_a[12] & input_a[5]);
  assign popcount28_ykzy_core_079 = ~(input_a[22] | input_a[15]);
  assign popcount28_ykzy_core_080 = ~(input_a[18] ^ input_a[5]);
  assign popcount28_ykzy_core_082 = ~(input_a[12] ^ input_a[19]);
  assign popcount28_ykzy_core_083 = ~(input_a[25] ^ input_a[16]);
  assign popcount28_ykzy_core_084 = ~(input_a[11] | input_a[16]);
  assign popcount28_ykzy_core_085 = input_a[23] & input_a[2];
  assign popcount28_ykzy_core_086_not = ~input_a[18];
  assign popcount28_ykzy_core_087 = input_a[8] ^ input_a[19];
  assign popcount28_ykzy_core_088 = input_a[23] | input_a[4];
  assign popcount28_ykzy_core_091 = ~(input_a[4] ^ input_a[17]);
  assign popcount28_ykzy_core_093 = ~input_a[14];
  assign popcount28_ykzy_core_097 = ~input_a[25];
  assign popcount28_ykzy_core_098 = ~(input_a[20] & input_a[22]);
  assign popcount28_ykzy_core_099 = ~input_a[22];
  assign popcount28_ykzy_core_102 = input_a[27] | input_a[5];
  assign popcount28_ykzy_core_103 = ~(input_a[25] & input_a[27]);
  assign popcount28_ykzy_core_104 = ~(input_a[24] ^ input_a[18]);
  assign popcount28_ykzy_core_106 = input_a[11] & input_a[3];
  assign popcount28_ykzy_core_107 = input_a[23] | input_a[2];
  assign popcount28_ykzy_core_108 = input_a[4] & input_a[20];
  assign popcount28_ykzy_core_109 = popcount28_ykzy_core_106 | popcount28_ykzy_core_108;
  assign popcount28_ykzy_core_112 = ~(input_a[20] ^ input_a[18]);
  assign popcount28_ykzy_core_113 = ~(input_a[10] ^ input_a[15]);
  assign popcount28_ykzy_core_114 = input_a[18] & input_a[12];
  assign popcount28_ykzy_core_116 = ~(input_a[0] & input_a[1]);
  assign popcount28_ykzy_core_117 = ~(input_a[21] | input_a[4]);
  assign popcount28_ykzy_core_118 = input_a[6] & input_a[17];
  assign popcount28_ykzy_core_119 = input_a[21] | input_a[17];
  assign popcount28_ykzy_core_120 = ~(input_a[15] & input_a[20]);
  assign popcount28_ykzy_core_121 = ~input_a[13];
  assign popcount28_ykzy_core_123 = input_a[2] & input_a[10];
  assign popcount28_ykzy_core_124 = popcount28_ykzy_core_109 ^ popcount28_ykzy_core_119;
  assign popcount28_ykzy_core_125 = popcount28_ykzy_core_109 & popcount28_ykzy_core_119;
  assign popcount28_ykzy_core_126 = popcount28_ykzy_core_124 ^ popcount28_ykzy_core_123;
  assign popcount28_ykzy_core_127 = popcount28_ykzy_core_124 & popcount28_ykzy_core_123;
  assign popcount28_ykzy_core_128 = popcount28_ykzy_core_125 | popcount28_ykzy_core_127;
  assign popcount28_ykzy_core_133 = input_a[11] ^ input_a[27];
  assign popcount28_ykzy_core_134 = ~input_a[8];
  assign popcount28_ykzy_core_135 = input_a[16] & input_a[9];
  assign popcount28_ykzy_core_137 = input_a[5] | input_a[14];
  assign popcount28_ykzy_core_139 = ~input_a[8];
  assign popcount28_ykzy_core_140 = input_a[4] ^ input_a[26];
  assign popcount28_ykzy_core_142 = input_a[6] & input_a[10];
  assign popcount28_ykzy_core_143 = input_a[7] & input_a[8];
  assign popcount28_ykzy_core_144 = ~(input_a[15] ^ input_a[8]);
  assign popcount28_ykzy_core_145 = input_a[18] & input_a[1];
  assign popcount28_ykzy_core_147 = input_a[1] | input_a[18];
  assign popcount28_ykzy_core_148 = popcount28_ykzy_core_143 | popcount28_ykzy_core_145;
  assign popcount28_ykzy_core_149 = ~(input_a[23] & input_a[2]);
  assign popcount28_ykzy_core_150 = ~(input_a[2] & input_a[17]);
  assign popcount28_ykzy_core_151 = ~(input_a[24] & input_a[2]);
  assign popcount28_ykzy_core_153 = popcount28_ykzy_core_135 ^ popcount28_ykzy_core_148;
  assign popcount28_ykzy_core_154 = popcount28_ykzy_core_135 & popcount28_ykzy_core_148;
  assign popcount28_ykzy_core_159 = ~(input_a[2] & input_a[12]);
  assign popcount28_ykzy_core_161 = ~(input_a[16] ^ input_a[27]);
  assign popcount28_ykzy_core_162 = input_a[3] | input_a[12];
  assign popcount28_ykzy_core_163 = ~(input_a[4] | input_a[22]);
  assign popcount28_ykzy_core_164 = ~input_a[24];
  assign popcount28_ykzy_core_165 = popcount28_ykzy_core_126 ^ popcount28_ykzy_core_153;
  assign popcount28_ykzy_core_166 = popcount28_ykzy_core_126 & popcount28_ykzy_core_153;
  assign popcount28_ykzy_core_168 = ~input_a[13];
  assign popcount28_ykzy_core_171 = popcount28_ykzy_core_128 & popcount28_ykzy_core_154;
  assign popcount28_ykzy_core_172 = ~(input_a[2] & input_a[8]);
  assign popcount28_ykzy_core_173 = popcount28_ykzy_core_128 & popcount28_ykzy_core_166;
  assign popcount28_ykzy_core_174 = popcount28_ykzy_core_171 | popcount28_ykzy_core_173;
  assign popcount28_ykzy_core_176 = ~(input_a[26] & input_a[22]);
  assign popcount28_ykzy_core_178 = ~input_a[9];
  assign popcount28_ykzy_core_180 = input_a[4] ^ input_a[2];
  assign popcount28_ykzy_core_181 = input_a[25] & input_a[24];
  assign popcount28_ykzy_core_182_not = ~popcount28_ykzy_core_165;
  assign popcount28_ykzy_core_184 = popcount28_ykzy_core_182_not ^ popcount28_ykzy_core_181;
  assign popcount28_ykzy_core_185 = input_a[24] & input_a[25];
  assign popcount28_ykzy_core_186 = popcount28_ykzy_core_165 | popcount28_ykzy_core_185;
  assign popcount28_ykzy_core_189_not = ~popcount28_ykzy_core_186;
  assign popcount28_ykzy_core_192 = popcount28_ykzy_core_102 ^ popcount28_ykzy_core_174;
  assign popcount28_ykzy_core_193 = popcount28_ykzy_core_102 & popcount28_ykzy_core_174;
  assign popcount28_ykzy_core_194 = popcount28_ykzy_core_192 ^ popcount28_ykzy_core_186;
  assign popcount28_ykzy_core_195 = popcount28_ykzy_core_192 & popcount28_ykzy_core_186;
  assign popcount28_ykzy_core_196 = popcount28_ykzy_core_193 | popcount28_ykzy_core_195;
  assign popcount28_ykzy_core_198 = ~(input_a[5] ^ input_a[18]);
  assign popcount28_ykzy_core_201 = ~(input_a[5] | input_a[8]);

  assign popcount28_ykzy_out[0] = input_a[12];
  assign popcount28_ykzy_out[1] = popcount28_ykzy_core_184;
  assign popcount28_ykzy_out[2] = popcount28_ykzy_core_189_not;
  assign popcount28_ykzy_out[3] = popcount28_ykzy_core_194;
  assign popcount28_ykzy_out[4] = popcount28_ykzy_core_196;
endmodule