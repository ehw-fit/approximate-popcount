// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.49708
// WCE=6.0
// EP=0.797477%
// Printed PDK parameters:
//  Area=51625074.0
//  Delay=69691200.0
//  Power=2557600.0

module popcount29_5oab(input [28:0] input_a, output [4:0] popcount29_5oab_out);
  wire popcount29_5oab_core_031;
  wire popcount29_5oab_core_032;
  wire popcount29_5oab_core_033;
  wire popcount29_5oab_core_034;
  wire popcount29_5oab_core_035;
  wire popcount29_5oab_core_037;
  wire popcount29_5oab_core_038;
  wire popcount29_5oab_core_039;
  wire popcount29_5oab_core_040;
  wire popcount29_5oab_core_041;
  wire popcount29_5oab_core_042;
  wire popcount29_5oab_core_043;
  wire popcount29_5oab_core_044;
  wire popcount29_5oab_core_045;
  wire popcount29_5oab_core_046;
  wire popcount29_5oab_core_048;
  wire popcount29_5oab_core_049;
  wire popcount29_5oab_core_050;
  wire popcount29_5oab_core_051;
  wire popcount29_5oab_core_052;
  wire popcount29_5oab_core_053;
  wire popcount29_5oab_core_054;
  wire popcount29_5oab_core_056;
  wire popcount29_5oab_core_057;
  wire popcount29_5oab_core_058;
  wire popcount29_5oab_core_061;
  wire popcount29_5oab_core_066;
  wire popcount29_5oab_core_067;
  wire popcount29_5oab_core_068;
  wire popcount29_5oab_core_069;
  wire popcount29_5oab_core_071;
  wire popcount29_5oab_core_072;
  wire popcount29_5oab_core_077;
  wire popcount29_5oab_core_079_not;
  wire popcount29_5oab_core_085;
  wire popcount29_5oab_core_089;
  wire popcount29_5oab_core_090;
  wire popcount29_5oab_core_091;
  wire popcount29_5oab_core_092;
  wire popcount29_5oab_core_094;
  wire popcount29_5oab_core_096;
  wire popcount29_5oab_core_097;
  wire popcount29_5oab_core_098;
  wire popcount29_5oab_core_099;
  wire popcount29_5oab_core_100;
  wire popcount29_5oab_core_102;
  wire popcount29_5oab_core_104;
  wire popcount29_5oab_core_107;
  wire popcount29_5oab_core_108;
  wire popcount29_5oab_core_109;
  wire popcount29_5oab_core_110;
  wire popcount29_5oab_core_112;
  wire popcount29_5oab_core_113;
  wire popcount29_5oab_core_114;
  wire popcount29_5oab_core_115;
  wire popcount29_5oab_core_116;
  wire popcount29_5oab_core_117;
  wire popcount29_5oab_core_118;
  wire popcount29_5oab_core_119;
  wire popcount29_5oab_core_120;
  wire popcount29_5oab_core_123;
  wire popcount29_5oab_core_124;
  wire popcount29_5oab_core_125;
  wire popcount29_5oab_core_126;
  wire popcount29_5oab_core_128;
  wire popcount29_5oab_core_131;
  wire popcount29_5oab_core_132;
  wire popcount29_5oab_core_135;
  wire popcount29_5oab_core_136;
  wire popcount29_5oab_core_137;
  wire popcount29_5oab_core_138;
  wire popcount29_5oab_core_139;
  wire popcount29_5oab_core_140;
  wire popcount29_5oab_core_141;
  wire popcount29_5oab_core_142;
  wire popcount29_5oab_core_143;
  wire popcount29_5oab_core_144;
  wire popcount29_5oab_core_146;
  wire popcount29_5oab_core_147;
  wire popcount29_5oab_core_148;
  wire popcount29_5oab_core_149;
  wire popcount29_5oab_core_150;
  wire popcount29_5oab_core_152;
  wire popcount29_5oab_core_153;
  wire popcount29_5oab_core_154;
  wire popcount29_5oab_core_155;
  wire popcount29_5oab_core_156;
  wire popcount29_5oab_core_158;
  wire popcount29_5oab_core_159;
  wire popcount29_5oab_core_160;
  wire popcount29_5oab_core_161;
  wire popcount29_5oab_core_162;
  wire popcount29_5oab_core_163;
  wire popcount29_5oab_core_164;
  wire popcount29_5oab_core_165;
  wire popcount29_5oab_core_166;
  wire popcount29_5oab_core_167;
  wire popcount29_5oab_core_168;
  wire popcount29_5oab_core_170;
  wire popcount29_5oab_core_171;
  wire popcount29_5oab_core_172;
  wire popcount29_5oab_core_174;
  wire popcount29_5oab_core_176;
  wire popcount29_5oab_core_177;
  wire popcount29_5oab_core_178;
  wire popcount29_5oab_core_179;
  wire popcount29_5oab_core_180;
  wire popcount29_5oab_core_183;
  wire popcount29_5oab_core_186;
  wire popcount29_5oab_core_188_not;
  wire popcount29_5oab_core_189;
  wire popcount29_5oab_core_190;
  wire popcount29_5oab_core_191;
  wire popcount29_5oab_core_193;
  wire popcount29_5oab_core_194;
  wire popcount29_5oab_core_195;
  wire popcount29_5oab_core_196;
  wire popcount29_5oab_core_197;
  wire popcount29_5oab_core_198;
  wire popcount29_5oab_core_199;
  wire popcount29_5oab_core_200;
  wire popcount29_5oab_core_201;
  wire popcount29_5oab_core_202;
  wire popcount29_5oab_core_207;

  assign popcount29_5oab_core_031 = input_a[10] & input_a[24];
  assign popcount29_5oab_core_032 = input_a[1] & input_a[2];
  assign popcount29_5oab_core_033 = ~(input_a[14] | input_a[11]);
  assign popcount29_5oab_core_034 = input_a[27] & input_a[0];
  assign popcount29_5oab_core_035 = popcount29_5oab_core_032 | popcount29_5oab_core_034;
  assign popcount29_5oab_core_037 = input_a[3] ^ input_a[4];
  assign popcount29_5oab_core_038 = input_a[3] & input_a[4];
  assign popcount29_5oab_core_039 = input_a[5] ^ input_a[6];
  assign popcount29_5oab_core_040 = input_a[5] & input_a[6];
  assign popcount29_5oab_core_041 = popcount29_5oab_core_037 ^ popcount29_5oab_core_039;
  assign popcount29_5oab_core_042 = popcount29_5oab_core_037 & popcount29_5oab_core_039;
  assign popcount29_5oab_core_043 = popcount29_5oab_core_038 ^ popcount29_5oab_core_040;
  assign popcount29_5oab_core_044 = popcount29_5oab_core_038 & popcount29_5oab_core_040;
  assign popcount29_5oab_core_045 = popcount29_5oab_core_043 | popcount29_5oab_core_042;
  assign popcount29_5oab_core_046 = ~input_a[10];
  assign popcount29_5oab_core_048 = input_a[23] ^ input_a[21];
  assign popcount29_5oab_core_049 = input_a[13] & popcount29_5oab_core_041;
  assign popcount29_5oab_core_050 = popcount29_5oab_core_035 ^ popcount29_5oab_core_045;
  assign popcount29_5oab_core_051 = popcount29_5oab_core_035 & popcount29_5oab_core_045;
  assign popcount29_5oab_core_052 = popcount29_5oab_core_050 ^ popcount29_5oab_core_049;
  assign popcount29_5oab_core_053 = popcount29_5oab_core_050 & popcount29_5oab_core_049;
  assign popcount29_5oab_core_054 = popcount29_5oab_core_051 | popcount29_5oab_core_053;
  assign popcount29_5oab_core_056 = ~(input_a[10] & input_a[0]);
  assign popcount29_5oab_core_057 = popcount29_5oab_core_044 | popcount29_5oab_core_054;
  assign popcount29_5oab_core_058 = input_a[28] ^ input_a[20];
  assign popcount29_5oab_core_061 = input_a[6] | input_a[15];
  assign popcount29_5oab_core_066 = input_a[4] & input_a[16];
  assign popcount29_5oab_core_067 = input_a[9] & input_a[11];
  assign popcount29_5oab_core_068 = input_a[20] ^ input_a[12];
  assign popcount29_5oab_core_069 = input_a[12] & input_a[8];
  assign popcount29_5oab_core_071 = ~(input_a[22] & input_a[19]);
  assign popcount29_5oab_core_072 = popcount29_5oab_core_067 | popcount29_5oab_core_069;
  assign popcount29_5oab_core_077 = input_a[1] & input_a[13];
  assign popcount29_5oab_core_079_not = ~popcount29_5oab_core_072;
  assign popcount29_5oab_core_085 = ~(input_a[5] | input_a[28]);
  assign popcount29_5oab_core_089 = input_a[9] & input_a[23];
  assign popcount29_5oab_core_090 = input_a[13] & input_a[6];
  assign popcount29_5oab_core_091 = popcount29_5oab_core_052 ^ popcount29_5oab_core_079_not;
  assign popcount29_5oab_core_092 = popcount29_5oab_core_052 & popcount29_5oab_core_079_not;
  assign popcount29_5oab_core_094 = input_a[10] | input_a[28];
  assign popcount29_5oab_core_096 = popcount29_5oab_core_057 ^ popcount29_5oab_core_072;
  assign popcount29_5oab_core_097 = popcount29_5oab_core_057 & popcount29_5oab_core_072;
  assign popcount29_5oab_core_098 = popcount29_5oab_core_096 ^ popcount29_5oab_core_092;
  assign popcount29_5oab_core_099 = popcount29_5oab_core_096 & popcount29_5oab_core_092;
  assign popcount29_5oab_core_100 = popcount29_5oab_core_097 | popcount29_5oab_core_099;
  assign popcount29_5oab_core_102 = input_a[28] | input_a[18];
  assign popcount29_5oab_core_104 = ~(input_a[28] ^ input_a[21]);
  assign popcount29_5oab_core_107 = input_a[15] & input_a[16];
  assign popcount29_5oab_core_108 = input_a[3] & input_a[5];
  assign popcount29_5oab_core_109 = input_a[14] & input_a[10];
  assign popcount29_5oab_core_110 = popcount29_5oab_core_107 | popcount29_5oab_core_109;
  assign popcount29_5oab_core_112 = input_a[17] | input_a[18];
  assign popcount29_5oab_core_113 = input_a[17] & input_a[18];
  assign popcount29_5oab_core_114 = input_a[19] ^ input_a[20];
  assign popcount29_5oab_core_115 = input_a[19] & input_a[20];
  assign popcount29_5oab_core_116 = ~input_a[19];
  assign popcount29_5oab_core_117 = popcount29_5oab_core_112 & popcount29_5oab_core_114;
  assign popcount29_5oab_core_118 = popcount29_5oab_core_113 ^ popcount29_5oab_core_115;
  assign popcount29_5oab_core_119 = popcount29_5oab_core_113 & popcount29_5oab_core_115;
  assign popcount29_5oab_core_120 = popcount29_5oab_core_118 | popcount29_5oab_core_117;
  assign popcount29_5oab_core_123 = ~(input_a[10] | input_a[22]);
  assign popcount29_5oab_core_124 = ~(input_a[0] | input_a[3]);
  assign popcount29_5oab_core_125 = popcount29_5oab_core_110 ^ popcount29_5oab_core_120;
  assign popcount29_5oab_core_126 = popcount29_5oab_core_110 & popcount29_5oab_core_120;
  assign popcount29_5oab_core_128 = ~(input_a[3] ^ input_a[24]);
  assign popcount29_5oab_core_131 = ~(input_a[8] ^ input_a[22]);
  assign popcount29_5oab_core_132 = popcount29_5oab_core_119 | popcount29_5oab_core_126;
  assign popcount29_5oab_core_135 = input_a[21] ^ input_a[22];
  assign popcount29_5oab_core_136 = input_a[21] & input_a[22];
  assign popcount29_5oab_core_137 = input_a[23] ^ input_a[24];
  assign popcount29_5oab_core_138 = input_a[23] & input_a[24];
  assign popcount29_5oab_core_139 = popcount29_5oab_core_135 ^ popcount29_5oab_core_137;
  assign popcount29_5oab_core_140 = popcount29_5oab_core_135 & popcount29_5oab_core_137;
  assign popcount29_5oab_core_141 = popcount29_5oab_core_136 ^ popcount29_5oab_core_138;
  assign popcount29_5oab_core_142 = popcount29_5oab_core_136 & popcount29_5oab_core_138;
  assign popcount29_5oab_core_143 = popcount29_5oab_core_141 | popcount29_5oab_core_140;
  assign popcount29_5oab_core_144 = input_a[2] ^ input_a[21];
  assign popcount29_5oab_core_146 = input_a[25] ^ input_a[26];
  assign popcount29_5oab_core_147 = input_a[25] & input_a[26];
  assign popcount29_5oab_core_148 = ~(input_a[20] | input_a[6]);
  assign popcount29_5oab_core_149 = input_a[7] & input_a[28];
  assign popcount29_5oab_core_150 = ~popcount29_5oab_core_146;
  assign popcount29_5oab_core_152 = popcount29_5oab_core_147 ^ popcount29_5oab_core_149;
  assign popcount29_5oab_core_153 = input_a[25] & popcount29_5oab_core_149;
  assign popcount29_5oab_core_154 = popcount29_5oab_core_152 ^ popcount29_5oab_core_146;
  assign popcount29_5oab_core_155 = popcount29_5oab_core_152 & popcount29_5oab_core_146;
  assign popcount29_5oab_core_156 = popcount29_5oab_core_153 | popcount29_5oab_core_155;
  assign popcount29_5oab_core_158 = popcount29_5oab_core_139 & popcount29_5oab_core_150;
  assign popcount29_5oab_core_159 = popcount29_5oab_core_143 ^ popcount29_5oab_core_154;
  assign popcount29_5oab_core_160 = popcount29_5oab_core_143 & popcount29_5oab_core_154;
  assign popcount29_5oab_core_161 = popcount29_5oab_core_159 ^ popcount29_5oab_core_158;
  assign popcount29_5oab_core_162 = popcount29_5oab_core_159 & popcount29_5oab_core_158;
  assign popcount29_5oab_core_163 = popcount29_5oab_core_160 | popcount29_5oab_core_162;
  assign popcount29_5oab_core_164 = popcount29_5oab_core_142 ^ popcount29_5oab_core_156;
  assign popcount29_5oab_core_165 = popcount29_5oab_core_142 & popcount29_5oab_core_156;
  assign popcount29_5oab_core_166 = popcount29_5oab_core_164 ^ popcount29_5oab_core_163;
  assign popcount29_5oab_core_167 = popcount29_5oab_core_164 & popcount29_5oab_core_163;
  assign popcount29_5oab_core_168 = popcount29_5oab_core_165 | popcount29_5oab_core_167;
  assign popcount29_5oab_core_170 = ~(input_a[16] | input_a[27]);
  assign popcount29_5oab_core_171 = popcount29_5oab_core_125 ^ popcount29_5oab_core_161;
  assign popcount29_5oab_core_172 = popcount29_5oab_core_125 & popcount29_5oab_core_161;
  assign popcount29_5oab_core_174 = ~input_a[10];
  assign popcount29_5oab_core_176 = popcount29_5oab_core_132 ^ popcount29_5oab_core_166;
  assign popcount29_5oab_core_177 = popcount29_5oab_core_132 & popcount29_5oab_core_166;
  assign popcount29_5oab_core_178 = popcount29_5oab_core_176 ^ popcount29_5oab_core_172;
  assign popcount29_5oab_core_179 = popcount29_5oab_core_176 & popcount29_5oab_core_172;
  assign popcount29_5oab_core_180 = popcount29_5oab_core_177 | popcount29_5oab_core_179;
  assign popcount29_5oab_core_183 = popcount29_5oab_core_168 | popcount29_5oab_core_180;
  assign popcount29_5oab_core_186 = ~(input_a[1] | input_a[5]);
  assign popcount29_5oab_core_188_not = ~input_a[15];
  assign popcount29_5oab_core_189 = popcount29_5oab_core_091 & popcount29_5oab_core_171;
  assign popcount29_5oab_core_190 = input_a[17] & input_a[21];
  assign popcount29_5oab_core_191 = input_a[0] ^ input_a[20];
  assign popcount29_5oab_core_193 = popcount29_5oab_core_098 ^ popcount29_5oab_core_178;
  assign popcount29_5oab_core_194 = popcount29_5oab_core_098 & popcount29_5oab_core_178;
  assign popcount29_5oab_core_195 = popcount29_5oab_core_193 ^ popcount29_5oab_core_189;
  assign popcount29_5oab_core_196 = popcount29_5oab_core_193 & popcount29_5oab_core_189;
  assign popcount29_5oab_core_197 = popcount29_5oab_core_194 | popcount29_5oab_core_196;
  assign popcount29_5oab_core_198 = popcount29_5oab_core_100 ^ popcount29_5oab_core_183;
  assign popcount29_5oab_core_199 = popcount29_5oab_core_100 & popcount29_5oab_core_183;
  assign popcount29_5oab_core_200 = popcount29_5oab_core_198 ^ popcount29_5oab_core_197;
  assign popcount29_5oab_core_201 = popcount29_5oab_core_198 & popcount29_5oab_core_197;
  assign popcount29_5oab_core_202 = popcount29_5oab_core_199 | popcount29_5oab_core_201;
  assign popcount29_5oab_core_207 = input_a[8] ^ input_a[19];

  assign popcount29_5oab_out[0] = 1'b1;
  assign popcount29_5oab_out[1] = 1'b1;
  assign popcount29_5oab_out[2] = popcount29_5oab_core_195;
  assign popcount29_5oab_out[3] = popcount29_5oab_core_200;
  assign popcount29_5oab_out[4] = popcount29_5oab_core_202;
endmodule