// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.65611
// WCE=20.0
// EP=0.922597%
// Printed PDK parameters:
//  Area=15567961.0
//  Delay=39393216.0
//  Power=666130.0

module popcount40_yc3h(input [39:0] input_a, output [5:0] popcount40_yc3h_out);
  wire popcount40_yc3h_core_042;
  wire popcount40_yc3h_core_043;
  wire popcount40_yc3h_core_044;
  wire popcount40_yc3h_core_045;
  wire popcount40_yc3h_core_046;
  wire popcount40_yc3h_core_047;
  wire popcount40_yc3h_core_049;
  wire popcount40_yc3h_core_050;
  wire popcount40_yc3h_core_051;
  wire popcount40_yc3h_core_052;
  wire popcount40_yc3h_core_053;
  wire popcount40_yc3h_core_056;
  wire popcount40_yc3h_core_057;
  wire popcount40_yc3h_core_058;
  wire popcount40_yc3h_core_059;
  wire popcount40_yc3h_core_061;
  wire popcount40_yc3h_core_063;
  wire popcount40_yc3h_core_064;
  wire popcount40_yc3h_core_066;
  wire popcount40_yc3h_core_067;
  wire popcount40_yc3h_core_069;
  wire popcount40_yc3h_core_071;
  wire popcount40_yc3h_core_072;
  wire popcount40_yc3h_core_073;
  wire popcount40_yc3h_core_076;
  wire popcount40_yc3h_core_077;
  wire popcount40_yc3h_core_080;
  wire popcount40_yc3h_core_081;
  wire popcount40_yc3h_core_084;
  wire popcount40_yc3h_core_087;
  wire popcount40_yc3h_core_088;
  wire popcount40_yc3h_core_089;
  wire popcount40_yc3h_core_090;
  wire popcount40_yc3h_core_094;
  wire popcount40_yc3h_core_095;
  wire popcount40_yc3h_core_096;
  wire popcount40_yc3h_core_097;
  wire popcount40_yc3h_core_098;
  wire popcount40_yc3h_core_099;
  wire popcount40_yc3h_core_101;
  wire popcount40_yc3h_core_105;
  wire popcount40_yc3h_core_106;
  wire popcount40_yc3h_core_107;
  wire popcount40_yc3h_core_109;
  wire popcount40_yc3h_core_110;
  wire popcount40_yc3h_core_114;
  wire popcount40_yc3h_core_116;
  wire popcount40_yc3h_core_118;
  wire popcount40_yc3h_core_120;
  wire popcount40_yc3h_core_121;
  wire popcount40_yc3h_core_123;
  wire popcount40_yc3h_core_124;
  wire popcount40_yc3h_core_125;
  wire popcount40_yc3h_core_127;
  wire popcount40_yc3h_core_128;
  wire popcount40_yc3h_core_132;
  wire popcount40_yc3h_core_133;
  wire popcount40_yc3h_core_134;
  wire popcount40_yc3h_core_135;
  wire popcount40_yc3h_core_137;
  wire popcount40_yc3h_core_139;
  wire popcount40_yc3h_core_142;
  wire popcount40_yc3h_core_144;
  wire popcount40_yc3h_core_145;
  wire popcount40_yc3h_core_146;
  wire popcount40_yc3h_core_147;
  wire popcount40_yc3h_core_148;
  wire popcount40_yc3h_core_149;
  wire popcount40_yc3h_core_151;
  wire popcount40_yc3h_core_153;
  wire popcount40_yc3h_core_154;
  wire popcount40_yc3h_core_155;
  wire popcount40_yc3h_core_156;
  wire popcount40_yc3h_core_157;
  wire popcount40_yc3h_core_158;
  wire popcount40_yc3h_core_159;
  wire popcount40_yc3h_core_160_not;
  wire popcount40_yc3h_core_164;
  wire popcount40_yc3h_core_167;
  wire popcount40_yc3h_core_168;
  wire popcount40_yc3h_core_169;
  wire popcount40_yc3h_core_170;
  wire popcount40_yc3h_core_171;
  wire popcount40_yc3h_core_172;
  wire popcount40_yc3h_core_173;
  wire popcount40_yc3h_core_174;
  wire popcount40_yc3h_core_175;
  wire popcount40_yc3h_core_176;
  wire popcount40_yc3h_core_177;
  wire popcount40_yc3h_core_178;
  wire popcount40_yc3h_core_179;
  wire popcount40_yc3h_core_181;
  wire popcount40_yc3h_core_185;
  wire popcount40_yc3h_core_186;
  wire popcount40_yc3h_core_187_not;
  wire popcount40_yc3h_core_190;
  wire popcount40_yc3h_core_194;
  wire popcount40_yc3h_core_195_not;
  wire popcount40_yc3h_core_196;
  wire popcount40_yc3h_core_197;
  wire popcount40_yc3h_core_198;
  wire popcount40_yc3h_core_201;
  wire popcount40_yc3h_core_202;
  wire popcount40_yc3h_core_204;
  wire popcount40_yc3h_core_205;
  wire popcount40_yc3h_core_206;
  wire popcount40_yc3h_core_209;
  wire popcount40_yc3h_core_210;
  wire popcount40_yc3h_core_219;
  wire popcount40_yc3h_core_220;
  wire popcount40_yc3h_core_221;
  wire popcount40_yc3h_core_223;
  wire popcount40_yc3h_core_224;
  wire popcount40_yc3h_core_225;
  wire popcount40_yc3h_core_226;
  wire popcount40_yc3h_core_227;
  wire popcount40_yc3h_core_230;
  wire popcount40_yc3h_core_231;
  wire popcount40_yc3h_core_232;
  wire popcount40_yc3h_core_233;
  wire popcount40_yc3h_core_234;
  wire popcount40_yc3h_core_237;
  wire popcount40_yc3h_core_238;
  wire popcount40_yc3h_core_239;
  wire popcount40_yc3h_core_240;
  wire popcount40_yc3h_core_242;
  wire popcount40_yc3h_core_243;
  wire popcount40_yc3h_core_244;
  wire popcount40_yc3h_core_246;
  wire popcount40_yc3h_core_247;
  wire popcount40_yc3h_core_248;
  wire popcount40_yc3h_core_249;
  wire popcount40_yc3h_core_250;
  wire popcount40_yc3h_core_251;
  wire popcount40_yc3h_core_252;
  wire popcount40_yc3h_core_253;
  wire popcount40_yc3h_core_254;
  wire popcount40_yc3h_core_255;
  wire popcount40_yc3h_core_260;
  wire popcount40_yc3h_core_261;
  wire popcount40_yc3h_core_264;
  wire popcount40_yc3h_core_267;
  wire popcount40_yc3h_core_268;
  wire popcount40_yc3h_core_269;
  wire popcount40_yc3h_core_271;
  wire popcount40_yc3h_core_272;
  wire popcount40_yc3h_core_275;
  wire popcount40_yc3h_core_276;
  wire popcount40_yc3h_core_277;
  wire popcount40_yc3h_core_278;
  wire popcount40_yc3h_core_279;
  wire popcount40_yc3h_core_280;
  wire popcount40_yc3h_core_281;
  wire popcount40_yc3h_core_282;
  wire popcount40_yc3h_core_283;
  wire popcount40_yc3h_core_284;
  wire popcount40_yc3h_core_289_not;
  wire popcount40_yc3h_core_291;
  wire popcount40_yc3h_core_292;
  wire popcount40_yc3h_core_294;
  wire popcount40_yc3h_core_295;
  wire popcount40_yc3h_core_297;
  wire popcount40_yc3h_core_298;
  wire popcount40_yc3h_core_299;
  wire popcount40_yc3h_core_300;
  wire popcount40_yc3h_core_301;
  wire popcount40_yc3h_core_302;
  wire popcount40_yc3h_core_303;
  wire popcount40_yc3h_core_304;
  wire popcount40_yc3h_core_305;
  wire popcount40_yc3h_core_306;
  wire popcount40_yc3h_core_309;
  wire popcount40_yc3h_core_310;
  wire popcount40_yc3h_core_312;
  wire popcount40_yc3h_core_314;
  wire popcount40_yc3h_core_316;

  assign popcount40_yc3h_core_042 = input_a[30] ^ input_a[33];
  assign popcount40_yc3h_core_043 = input_a[0] | input_a[10];
  assign popcount40_yc3h_core_044 = ~(input_a[15] | input_a[36]);
  assign popcount40_yc3h_core_045 = ~(input_a[11] | input_a[18]);
  assign popcount40_yc3h_core_046 = input_a[39] ^ input_a[17];
  assign popcount40_yc3h_core_047 = ~(input_a[34] | input_a[6]);
  assign popcount40_yc3h_core_049 = input_a[4] & input_a[8];
  assign popcount40_yc3h_core_050 = ~(input_a[5] | input_a[25]);
  assign popcount40_yc3h_core_051 = ~(input_a[32] ^ input_a[33]);
  assign popcount40_yc3h_core_052 = input_a[26] | input_a[26];
  assign popcount40_yc3h_core_053 = input_a[6] & input_a[4];
  assign popcount40_yc3h_core_056 = ~(input_a[26] & input_a[12]);
  assign popcount40_yc3h_core_057 = input_a[27] ^ input_a[35];
  assign popcount40_yc3h_core_058 = input_a[5] & input_a[15];
  assign popcount40_yc3h_core_059 = input_a[11] ^ input_a[30];
  assign popcount40_yc3h_core_061 = input_a[20] | input_a[32];
  assign popcount40_yc3h_core_063 = ~(input_a[24] & input_a[35]);
  assign popcount40_yc3h_core_064 = input_a[10] ^ input_a[37];
  assign popcount40_yc3h_core_066 = input_a[13] ^ input_a[1];
  assign popcount40_yc3h_core_067 = input_a[30] | input_a[32];
  assign popcount40_yc3h_core_069 = input_a[9] | input_a[32];
  assign popcount40_yc3h_core_071 = input_a[20] | input_a[10];
  assign popcount40_yc3h_core_072 = ~(input_a[0] ^ input_a[9]);
  assign popcount40_yc3h_core_073 = input_a[12] & input_a[28];
  assign popcount40_yc3h_core_076 = input_a[34] ^ input_a[1];
  assign popcount40_yc3h_core_077 = input_a[29] | input_a[39];
  assign popcount40_yc3h_core_080 = input_a[35] & input_a[14];
  assign popcount40_yc3h_core_081 = input_a[36] | input_a[38];
  assign popcount40_yc3h_core_084 = input_a[12] & input_a[6];
  assign popcount40_yc3h_core_087 = input_a[25] | input_a[34];
  assign popcount40_yc3h_core_088 = ~input_a[1];
  assign popcount40_yc3h_core_089 = input_a[2] ^ input_a[7];
  assign popcount40_yc3h_core_090 = input_a[30] ^ input_a[4];
  assign popcount40_yc3h_core_094 = ~(input_a[10] | input_a[30]);
  assign popcount40_yc3h_core_095 = ~(input_a[23] & input_a[2]);
  assign popcount40_yc3h_core_096 = ~(input_a[14] | input_a[11]);
  assign popcount40_yc3h_core_097 = input_a[28] | input_a[2];
  assign popcount40_yc3h_core_098 = ~input_a[2];
  assign popcount40_yc3h_core_099 = ~(input_a[2] ^ input_a[30]);
  assign popcount40_yc3h_core_101 = ~input_a[16];
  assign popcount40_yc3h_core_105 = input_a[18] ^ input_a[23];
  assign popcount40_yc3h_core_106 = input_a[36] | input_a[18];
  assign popcount40_yc3h_core_107 = ~input_a[9];
  assign popcount40_yc3h_core_109 = input_a[29] | input_a[12];
  assign popcount40_yc3h_core_110 = ~input_a[20];
  assign popcount40_yc3h_core_114 = input_a[31] & input_a[11];
  assign popcount40_yc3h_core_116 = input_a[7] | input_a[6];
  assign popcount40_yc3h_core_118 = ~(input_a[10] | input_a[36]);
  assign popcount40_yc3h_core_120 = ~(input_a[9] | input_a[6]);
  assign popcount40_yc3h_core_121 = ~(input_a[15] | input_a[15]);
  assign popcount40_yc3h_core_123 = input_a[11] | input_a[14];
  assign popcount40_yc3h_core_124 = ~(input_a[0] & input_a[3]);
  assign popcount40_yc3h_core_125 = input_a[16] ^ input_a[24];
  assign popcount40_yc3h_core_127 = ~(input_a[34] ^ input_a[28]);
  assign popcount40_yc3h_core_128 = ~(input_a[31] ^ input_a[24]);
  assign popcount40_yc3h_core_132 = input_a[0] ^ input_a[31];
  assign popcount40_yc3h_core_133 = ~input_a[23];
  assign popcount40_yc3h_core_134 = ~(input_a[31] & input_a[6]);
  assign popcount40_yc3h_core_135 = input_a[34] ^ input_a[10];
  assign popcount40_yc3h_core_137 = input_a[35] ^ input_a[38];
  assign popcount40_yc3h_core_139 = ~input_a[4];
  assign popcount40_yc3h_core_142 = ~(input_a[34] ^ input_a[23]);
  assign popcount40_yc3h_core_144 = ~(input_a[2] ^ input_a[16]);
  assign popcount40_yc3h_core_145 = ~input_a[10];
  assign popcount40_yc3h_core_146 = input_a[4] ^ input_a[9];
  assign popcount40_yc3h_core_147 = input_a[27] & input_a[10];
  assign popcount40_yc3h_core_148 = ~(input_a[14] & input_a[39]);
  assign popcount40_yc3h_core_149 = ~(input_a[36] | input_a[25]);
  assign popcount40_yc3h_core_151 = input_a[5] & input_a[3];
  assign popcount40_yc3h_core_153 = input_a[21] | input_a[8];
  assign popcount40_yc3h_core_154 = ~(input_a[37] & input_a[10]);
  assign popcount40_yc3h_core_155 = ~(input_a[15] ^ input_a[18]);
  assign popcount40_yc3h_core_156 = input_a[11] | input_a[30];
  assign popcount40_yc3h_core_157 = ~input_a[21];
  assign popcount40_yc3h_core_158 = input_a[39] | input_a[24];
  assign popcount40_yc3h_core_159 = input_a[18] ^ input_a[13];
  assign popcount40_yc3h_core_160_not = ~input_a[31];
  assign popcount40_yc3h_core_164 = input_a[25] ^ input_a[14];
  assign popcount40_yc3h_core_167 = input_a[20] & input_a[37];
  assign popcount40_yc3h_core_168 = ~(input_a[25] ^ input_a[24]);
  assign popcount40_yc3h_core_169 = input_a[32] & input_a[31];
  assign popcount40_yc3h_core_170 = input_a[27] ^ input_a[8];
  assign popcount40_yc3h_core_171 = input_a[2] & input_a[23];
  assign popcount40_yc3h_core_172 = popcount40_yc3h_core_169 | popcount40_yc3h_core_171;
  assign popcount40_yc3h_core_173 = popcount40_yc3h_core_169 & popcount40_yc3h_core_171;
  assign popcount40_yc3h_core_174 = input_a[6] ^ input_a[17];
  assign popcount40_yc3h_core_175 = input_a[19] ^ input_a[23];
  assign popcount40_yc3h_core_176 = input_a[29] & input_a[27];
  assign popcount40_yc3h_core_177 = popcount40_yc3h_core_167 & popcount40_yc3h_core_172;
  assign popcount40_yc3h_core_178 = input_a[28] & input_a[30];
  assign popcount40_yc3h_core_179 = ~(input_a[32] | input_a[24]);
  assign popcount40_yc3h_core_181 = popcount40_yc3h_core_173 | popcount40_yc3h_core_177;
  assign popcount40_yc3h_core_185 = input_a[28] | input_a[22];
  assign popcount40_yc3h_core_186 = ~(input_a[31] & input_a[1]);
  assign popcount40_yc3h_core_187_not = ~input_a[2];
  assign popcount40_yc3h_core_190 = ~(input_a[17] ^ input_a[29]);
  assign popcount40_yc3h_core_194 = ~(input_a[18] ^ input_a[28]);
  assign popcount40_yc3h_core_195_not = ~input_a[21];
  assign popcount40_yc3h_core_196 = input_a[10] | input_a[39];
  assign popcount40_yc3h_core_197 = ~(input_a[14] ^ input_a[30]);
  assign popcount40_yc3h_core_198 = input_a[31] | input_a[17];
  assign popcount40_yc3h_core_201 = input_a[0] & input_a[15];
  assign popcount40_yc3h_core_202 = ~popcount40_yc3h_core_178;
  assign popcount40_yc3h_core_204 = popcount40_yc3h_core_202 ^ popcount40_yc3h_core_201;
  assign popcount40_yc3h_core_205 = input_a[0] & input_a[15];
  assign popcount40_yc3h_core_206 = popcount40_yc3h_core_178 | popcount40_yc3h_core_205;
  assign popcount40_yc3h_core_209 = popcount40_yc3h_core_181 ^ popcount40_yc3h_core_206;
  assign popcount40_yc3h_core_210 = popcount40_yc3h_core_181 & popcount40_yc3h_core_206;
  assign popcount40_yc3h_core_219 = ~(input_a[29] & input_a[38]);
  assign popcount40_yc3h_core_220 = input_a[12] ^ input_a[27];
  assign popcount40_yc3h_core_221 = input_a[21] & input_a[28];
  assign popcount40_yc3h_core_223 = input_a[0] ^ input_a[1];
  assign popcount40_yc3h_core_224 = ~(input_a[26] & input_a[33]);
  assign popcount40_yc3h_core_225 = ~(input_a[25] & input_a[22]);
  assign popcount40_yc3h_core_226 = ~input_a[26];
  assign popcount40_yc3h_core_227 = ~(input_a[23] ^ input_a[8]);
  assign popcount40_yc3h_core_230 = ~input_a[26];
  assign popcount40_yc3h_core_231 = input_a[39] | input_a[19];
  assign popcount40_yc3h_core_232 = input_a[4] ^ input_a[34];
  assign popcount40_yc3h_core_233 = ~(input_a[25] ^ input_a[30]);
  assign popcount40_yc3h_core_234 = ~input_a[10];
  assign popcount40_yc3h_core_237 = ~input_a[15];
  assign popcount40_yc3h_core_238 = ~input_a[30];
  assign popcount40_yc3h_core_239 = ~(input_a[18] | input_a[14]);
  assign popcount40_yc3h_core_240 = input_a[13] & input_a[0];
  assign popcount40_yc3h_core_242 = ~(input_a[26] ^ input_a[20]);
  assign popcount40_yc3h_core_243 = ~(input_a[36] ^ input_a[24]);
  assign popcount40_yc3h_core_244 = ~(input_a[27] | input_a[8]);
  assign popcount40_yc3h_core_246 = ~(input_a[9] ^ input_a[31]);
  assign popcount40_yc3h_core_247 = ~input_a[33];
  assign popcount40_yc3h_core_248 = ~(input_a[11] | input_a[18]);
  assign popcount40_yc3h_core_249 = ~(input_a[1] | input_a[18]);
  assign popcount40_yc3h_core_250 = input_a[38] & input_a[20];
  assign popcount40_yc3h_core_251 = ~(input_a[24] & input_a[24]);
  assign popcount40_yc3h_core_252 = ~(input_a[23] | input_a[27]);
  assign popcount40_yc3h_core_253 = ~(input_a[29] & input_a[30]);
  assign popcount40_yc3h_core_254 = input_a[20] | input_a[19];
  assign popcount40_yc3h_core_255 = ~(input_a[4] & input_a[36]);
  assign popcount40_yc3h_core_260 = ~(input_a[4] & input_a[36]);
  assign popcount40_yc3h_core_261 = input_a[4] & input_a[36];
  assign popcount40_yc3h_core_264 = ~(input_a[39] | input_a[37]);
  assign popcount40_yc3h_core_267 = ~(input_a[20] ^ input_a[13]);
  assign popcount40_yc3h_core_268 = ~(input_a[14] ^ input_a[31]);
  assign popcount40_yc3h_core_269 = input_a[39] & input_a[17];
  assign popcount40_yc3h_core_271 = popcount40_yc3h_core_204 & popcount40_yc3h_core_255;
  assign popcount40_yc3h_core_272 = ~(input_a[21] & input_a[39]);
  assign popcount40_yc3h_core_275 = popcount40_yc3h_core_209 ^ popcount40_yc3h_core_260;
  assign popcount40_yc3h_core_276 = popcount40_yc3h_core_209 & popcount40_yc3h_core_260;
  assign popcount40_yc3h_core_277 = popcount40_yc3h_core_275 ^ popcount40_yc3h_core_271;
  assign popcount40_yc3h_core_278 = popcount40_yc3h_core_275 & popcount40_yc3h_core_271;
  assign popcount40_yc3h_core_279 = popcount40_yc3h_core_276 | popcount40_yc3h_core_278;
  assign popcount40_yc3h_core_280 = popcount40_yc3h_core_210 ^ popcount40_yc3h_core_261;
  assign popcount40_yc3h_core_281 = popcount40_yc3h_core_210 & popcount40_yc3h_core_261;
  assign popcount40_yc3h_core_282 = popcount40_yc3h_core_280 ^ popcount40_yc3h_core_279;
  assign popcount40_yc3h_core_283 = popcount40_yc3h_core_280 & popcount40_yc3h_core_279;
  assign popcount40_yc3h_core_284 = popcount40_yc3h_core_281 | popcount40_yc3h_core_283;
  assign popcount40_yc3h_core_289_not = ~input_a[20];
  assign popcount40_yc3h_core_291 = ~(input_a[31] | input_a[23]);
  assign popcount40_yc3h_core_292 = ~(input_a[17] | input_a[33]);
  assign popcount40_yc3h_core_294 = ~(input_a[33] & input_a[27]);
  assign popcount40_yc3h_core_295 = input_a[27] & input_a[33];
  assign popcount40_yc3h_core_297 = popcount40_yc3h_core_153 ^ popcount40_yc3h_core_277;
  assign popcount40_yc3h_core_298 = popcount40_yc3h_core_153 & popcount40_yc3h_core_277;
  assign popcount40_yc3h_core_299 = popcount40_yc3h_core_297 ^ popcount40_yc3h_core_295;
  assign popcount40_yc3h_core_300 = popcount40_yc3h_core_297 & popcount40_yc3h_core_295;
  assign popcount40_yc3h_core_301 = popcount40_yc3h_core_298 | popcount40_yc3h_core_300;
  assign popcount40_yc3h_core_302 = popcount40_yc3h_core_158 ^ popcount40_yc3h_core_282;
  assign popcount40_yc3h_core_303 = popcount40_yc3h_core_158 & popcount40_yc3h_core_282;
  assign popcount40_yc3h_core_304 = popcount40_yc3h_core_302 ^ popcount40_yc3h_core_301;
  assign popcount40_yc3h_core_305 = popcount40_yc3h_core_302 & popcount40_yc3h_core_301;
  assign popcount40_yc3h_core_306 = popcount40_yc3h_core_303 | popcount40_yc3h_core_305;
  assign popcount40_yc3h_core_309 = popcount40_yc3h_core_284 ^ popcount40_yc3h_core_306;
  assign popcount40_yc3h_core_310 = popcount40_yc3h_core_284 & popcount40_yc3h_core_306;
  assign popcount40_yc3h_core_312 = input_a[27] & input_a[7];
  assign popcount40_yc3h_core_314 = input_a[31] & input_a[27];
  assign popcount40_yc3h_core_316 = input_a[15] | input_a[21];

  assign popcount40_yc3h_out[0] = input_a[1];
  assign popcount40_yc3h_out[1] = popcount40_yc3h_core_294;
  assign popcount40_yc3h_out[2] = popcount40_yc3h_core_299;
  assign popcount40_yc3h_out[3] = popcount40_yc3h_core_304;
  assign popcount40_yc3h_out[4] = popcount40_yc3h_core_309;
  assign popcount40_yc3h_out[5] = popcount40_yc3h_core_310;
endmodule