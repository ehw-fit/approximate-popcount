// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.59882
// WCE=11.0
// EP=0.805995%
// Printed PDK parameters:
//  Area=38356024.0
//  Delay=60254912.0
//  Power=1727100.0

module popcount32_cdyi(input [31:0] input_a, output [5:0] popcount32_cdyi_out);
  wire popcount32_cdyi_core_034;
  wire popcount32_cdyi_core_035;
  wire popcount32_cdyi_core_037;
  wire popcount32_cdyi_core_039;
  wire popcount32_cdyi_core_040;
  wire popcount32_cdyi_core_041;
  wire popcount32_cdyi_core_042;
  wire popcount32_cdyi_core_043;
  wire popcount32_cdyi_core_045;
  wire popcount32_cdyi_core_049;
  wire popcount32_cdyi_core_050_not;
  wire popcount32_cdyi_core_053;
  wire popcount32_cdyi_core_054;
  wire popcount32_cdyi_core_056;
  wire popcount32_cdyi_core_058;
  wire popcount32_cdyi_core_060;
  wire popcount32_cdyi_core_061;
  wire popcount32_cdyi_core_064;
  wire popcount32_cdyi_core_065;
  wire popcount32_cdyi_core_067;
  wire popcount32_cdyi_core_068;
  wire popcount32_cdyi_core_069;
  wire popcount32_cdyi_core_071;
  wire popcount32_cdyi_core_073;
  wire popcount32_cdyi_core_074;
  wire popcount32_cdyi_core_075;
  wire popcount32_cdyi_core_077;
  wire popcount32_cdyi_core_079;
  wire popcount32_cdyi_core_081;
  wire popcount32_cdyi_core_082;
  wire popcount32_cdyi_core_084;
  wire popcount32_cdyi_core_085;
  wire popcount32_cdyi_core_087;
  wire popcount32_cdyi_core_089;
  wire popcount32_cdyi_core_092;
  wire popcount32_cdyi_core_093;
  wire popcount32_cdyi_core_098;
  wire popcount32_cdyi_core_099;
  wire popcount32_cdyi_core_102;
  wire popcount32_cdyi_core_103;
  wire popcount32_cdyi_core_104;
  wire popcount32_cdyi_core_105;
  wire popcount32_cdyi_core_106;
  wire popcount32_cdyi_core_107;
  wire popcount32_cdyi_core_108;
  wire popcount32_cdyi_core_109;
  wire popcount32_cdyi_core_110;
  wire popcount32_cdyi_core_111;
  wire popcount32_cdyi_core_112;
  wire popcount32_cdyi_core_113;
  wire popcount32_cdyi_core_117;
  wire popcount32_cdyi_core_120;
  wire popcount32_cdyi_core_122;
  wire popcount32_cdyi_core_123;
  wire popcount32_cdyi_core_124;
  wire popcount32_cdyi_core_125;
  wire popcount32_cdyi_core_127;
  wire popcount32_cdyi_core_128;
  wire popcount32_cdyi_core_129;
  wire popcount32_cdyi_core_131;
  wire popcount32_cdyi_core_132;
  wire popcount32_cdyi_core_134;
  wire popcount32_cdyi_core_137;
  wire popcount32_cdyi_core_139;
  wire popcount32_cdyi_core_141;
  wire popcount32_cdyi_core_143;
  wire popcount32_cdyi_core_144;
  wire popcount32_cdyi_core_146;
  wire popcount32_cdyi_core_149;
  wire popcount32_cdyi_core_151;
  wire popcount32_cdyi_core_152_not;
  wire popcount32_cdyi_core_154;
  wire popcount32_cdyi_core_155;
  wire popcount32_cdyi_core_156;
  wire popcount32_cdyi_core_157;
  wire popcount32_cdyi_core_158;
  wire popcount32_cdyi_core_159;
  wire popcount32_cdyi_core_160;
  wire popcount32_cdyi_core_161;
  wire popcount32_cdyi_core_163;
  wire popcount32_cdyi_core_164;
  wire popcount32_cdyi_core_165;
  wire popcount32_cdyi_core_166;
  wire popcount32_cdyi_core_167;
  wire popcount32_cdyi_core_169;
  wire popcount32_cdyi_core_170;
  wire popcount32_cdyi_core_171;
  wire popcount32_cdyi_core_172;
  wire popcount32_cdyi_core_173;
  wire popcount32_cdyi_core_174;
  wire popcount32_cdyi_core_175;
  wire popcount32_cdyi_core_176;
  wire popcount32_cdyi_core_177;
  wire popcount32_cdyi_core_178;
  wire popcount32_cdyi_core_179;
  wire popcount32_cdyi_core_180;
  wire popcount32_cdyi_core_181;
  wire popcount32_cdyi_core_183;
  wire popcount32_cdyi_core_185;
  wire popcount32_cdyi_core_186;
  wire popcount32_cdyi_core_187;
  wire popcount32_cdyi_core_189;
  wire popcount32_cdyi_core_191;
  wire popcount32_cdyi_core_193;
  wire popcount32_cdyi_core_194;
  wire popcount32_cdyi_core_195;
  wire popcount32_cdyi_core_196;
  wire popcount32_cdyi_core_197;
  wire popcount32_cdyi_core_198;
  wire popcount32_cdyi_core_200;
  wire popcount32_cdyi_core_203;
  wire popcount32_cdyi_core_204;
  wire popcount32_cdyi_core_206;
  wire popcount32_cdyi_core_208;
  wire popcount32_cdyi_core_210;
  wire popcount32_cdyi_core_211;
  wire popcount32_cdyi_core_212;
  wire popcount32_cdyi_core_213;
  wire popcount32_cdyi_core_214;
  wire popcount32_cdyi_core_215;
  wire popcount32_cdyi_core_216;
  wire popcount32_cdyi_core_217;
  wire popcount32_cdyi_core_218;
  wire popcount32_cdyi_core_219;
  wire popcount32_cdyi_core_220;
  wire popcount32_cdyi_core_222;
  wire popcount32_cdyi_core_224;

  assign popcount32_cdyi_core_034 = ~(input_a[31] & input_a[4]);
  assign popcount32_cdyi_core_035 = input_a[23] & input_a[14];
  assign popcount32_cdyi_core_037 = input_a[20] | input_a[14];
  assign popcount32_cdyi_core_039 = input_a[7] & input_a[9];
  assign popcount32_cdyi_core_040 = input_a[11] | input_a[27];
  assign popcount32_cdyi_core_041 = ~input_a[10];
  assign popcount32_cdyi_core_042 = popcount32_cdyi_core_040 | popcount32_cdyi_core_039;
  assign popcount32_cdyi_core_043 = ~input_a[16];
  assign popcount32_cdyi_core_045 = ~(input_a[12] | input_a[6]);
  assign popcount32_cdyi_core_049 = ~input_a[6];
  assign popcount32_cdyi_core_050_not = ~input_a[10];
  assign popcount32_cdyi_core_053 = ~(input_a[17] & input_a[21]);
  assign popcount32_cdyi_core_054 = ~input_a[11];
  assign popcount32_cdyi_core_056 = ~(input_a[11] & input_a[8]);
  assign popcount32_cdyi_core_058 = popcount32_cdyi_core_042 ^ input_a[6];
  assign popcount32_cdyi_core_060 = popcount32_cdyi_core_058 ^ popcount32_cdyi_core_049;
  assign popcount32_cdyi_core_061 = ~input_a[2];
  assign popcount32_cdyi_core_064 = input_a[21] & input_a[17];
  assign popcount32_cdyi_core_065 = input_a[11] | popcount32_cdyi_core_042;
  assign popcount32_cdyi_core_067 = input_a[16] ^ input_a[16];
  assign popcount32_cdyi_core_068 = input_a[2] & input_a[5];
  assign popcount32_cdyi_core_069 = input_a[19] & input_a[15];
  assign popcount32_cdyi_core_071 = input_a[24] & input_a[29];
  assign popcount32_cdyi_core_073 = input_a[14] & input_a[20];
  assign popcount32_cdyi_core_074 = popcount32_cdyi_core_069 ^ popcount32_cdyi_core_071;
  assign popcount32_cdyi_core_075 = popcount32_cdyi_core_069 & popcount32_cdyi_core_071;
  assign popcount32_cdyi_core_077 = input_a[4] ^ input_a[6];
  assign popcount32_cdyi_core_079 = ~(input_a[22] ^ input_a[29]);
  assign popcount32_cdyi_core_081 = input_a[8] & input_a[24];
  assign popcount32_cdyi_core_082 = input_a[0] | input_a[9];
  assign popcount32_cdyi_core_084 = input_a[29] ^ input_a[24];
  assign popcount32_cdyi_core_085 = input_a[17] ^ input_a[22];
  assign popcount32_cdyi_core_087 = input_a[26] | input_a[16];
  assign popcount32_cdyi_core_089 = input_a[27] ^ input_a[17];
  assign popcount32_cdyi_core_092 = popcount32_cdyi_core_074 ^ popcount32_cdyi_core_087;
  assign popcount32_cdyi_core_093 = popcount32_cdyi_core_074 & popcount32_cdyi_core_087;
  assign popcount32_cdyi_core_098 = input_a[1] ^ input_a[5];
  assign popcount32_cdyi_core_099 = popcount32_cdyi_core_075 | popcount32_cdyi_core_093;
  assign popcount32_cdyi_core_102 = input_a[12] & input_a[28];
  assign popcount32_cdyi_core_103 = input_a[8] & input_a[21];
  assign popcount32_cdyi_core_104 = popcount32_cdyi_core_060 ^ popcount32_cdyi_core_092;
  assign popcount32_cdyi_core_105 = popcount32_cdyi_core_060 & popcount32_cdyi_core_092;
  assign popcount32_cdyi_core_106 = popcount32_cdyi_core_104 ^ popcount32_cdyi_core_103;
  assign popcount32_cdyi_core_107 = popcount32_cdyi_core_104 & popcount32_cdyi_core_103;
  assign popcount32_cdyi_core_108 = popcount32_cdyi_core_105 | popcount32_cdyi_core_107;
  assign popcount32_cdyi_core_109 = popcount32_cdyi_core_065 ^ popcount32_cdyi_core_099;
  assign popcount32_cdyi_core_110 = popcount32_cdyi_core_065 & popcount32_cdyi_core_099;
  assign popcount32_cdyi_core_111 = popcount32_cdyi_core_109 ^ popcount32_cdyi_core_108;
  assign popcount32_cdyi_core_112 = popcount32_cdyi_core_109 & popcount32_cdyi_core_108;
  assign popcount32_cdyi_core_113 = popcount32_cdyi_core_110 | popcount32_cdyi_core_112;
  assign popcount32_cdyi_core_117 = input_a[6] | input_a[29];
  assign popcount32_cdyi_core_120 = input_a[8] ^ input_a[11];
  assign popcount32_cdyi_core_122 = ~(input_a[25] ^ input_a[19]);
  assign popcount32_cdyi_core_123 = input_a[21] ^ input_a[12];
  assign popcount32_cdyi_core_124 = ~input_a[2];
  assign popcount32_cdyi_core_125 = input_a[15] | input_a[21];
  assign popcount32_cdyi_core_127 = input_a[10] | input_a[6];
  assign popcount32_cdyi_core_128 = ~input_a[18];
  assign popcount32_cdyi_core_129 = input_a[12] & input_a[5];
  assign popcount32_cdyi_core_131 = input_a[12] & input_a[1];
  assign popcount32_cdyi_core_132 = ~(input_a[13] & input_a[3]);
  assign popcount32_cdyi_core_134 = ~(input_a[21] | input_a[4]);
  assign popcount32_cdyi_core_137 = ~(input_a[30] ^ input_a[18]);
  assign popcount32_cdyi_core_139 = input_a[14] | input_a[23];
  assign popcount32_cdyi_core_141 = input_a[31] ^ input_a[21];
  assign popcount32_cdyi_core_143 = popcount32_cdyi_core_127 ^ popcount32_cdyi_core_131;
  assign popcount32_cdyi_core_144 = popcount32_cdyi_core_127 & popcount32_cdyi_core_131;
  assign popcount32_cdyi_core_146 = input_a[21] & input_a[15];
  assign popcount32_cdyi_core_149 = ~(input_a[21] ^ input_a[27]);
  assign popcount32_cdyi_core_151 = ~input_a[19];
  assign popcount32_cdyi_core_152_not = ~input_a[4];
  assign popcount32_cdyi_core_154 = input_a[5] & input_a[0];
  assign popcount32_cdyi_core_155 = ~(input_a[3] | input_a[24]);
  assign popcount32_cdyi_core_156 = input_a[25] & input_a[9];
  assign popcount32_cdyi_core_157 = ~(input_a[3] ^ input_a[3]);
  assign popcount32_cdyi_core_158 = input_a[2] & input_a[28];
  assign popcount32_cdyi_core_159 = popcount32_cdyi_core_154 | popcount32_cdyi_core_156;
  assign popcount32_cdyi_core_160 = input_a[26] | input_a[1];
  assign popcount32_cdyi_core_161 = popcount32_cdyi_core_159 | popcount32_cdyi_core_158;
  assign popcount32_cdyi_core_163 = ~(input_a[3] & input_a[31]);
  assign popcount32_cdyi_core_164 = input_a[27] & input_a[25];
  assign popcount32_cdyi_core_165 = input_a[18] & input_a[20];
  assign popcount32_cdyi_core_166 = ~(input_a[6] ^ input_a[26]);
  assign popcount32_cdyi_core_167 = input_a[14] & input_a[17];
  assign popcount32_cdyi_core_169 = input_a[30] & input_a[22];
  assign popcount32_cdyi_core_170 = popcount32_cdyi_core_165 | popcount32_cdyi_core_167;
  assign popcount32_cdyi_core_171 = input_a[0] & input_a[30];
  assign popcount32_cdyi_core_172 = popcount32_cdyi_core_170 | popcount32_cdyi_core_169;
  assign popcount32_cdyi_core_173 = input_a[13] & input_a[2];
  assign popcount32_cdyi_core_174 = ~input_a[27];
  assign popcount32_cdyi_core_175 = ~(input_a[15] | input_a[21]);
  assign popcount32_cdyi_core_176 = input_a[4] & input_a[23];
  assign popcount32_cdyi_core_177 = popcount32_cdyi_core_161 ^ popcount32_cdyi_core_172;
  assign popcount32_cdyi_core_178 = popcount32_cdyi_core_161 & popcount32_cdyi_core_172;
  assign popcount32_cdyi_core_179 = popcount32_cdyi_core_177 ^ popcount32_cdyi_core_176;
  assign popcount32_cdyi_core_180 = popcount32_cdyi_core_177 & popcount32_cdyi_core_176;
  assign popcount32_cdyi_core_181 = popcount32_cdyi_core_178 | popcount32_cdyi_core_180;
  assign popcount32_cdyi_core_183 = ~(input_a[22] ^ input_a[21]);
  assign popcount32_cdyi_core_185 = ~(input_a[21] ^ input_a[31]);
  assign popcount32_cdyi_core_186 = ~input_a[13];
  assign popcount32_cdyi_core_187 = ~(input_a[4] ^ input_a[29]);
  assign popcount32_cdyi_core_189 = popcount32_cdyi_core_143 ^ popcount32_cdyi_core_179;
  assign popcount32_cdyi_core_191 = ~popcount32_cdyi_core_189;
  assign popcount32_cdyi_core_193 = popcount32_cdyi_core_143 | popcount32_cdyi_core_189;
  assign popcount32_cdyi_core_194 = popcount32_cdyi_core_144 ^ popcount32_cdyi_core_181;
  assign popcount32_cdyi_core_195 = popcount32_cdyi_core_144 & popcount32_cdyi_core_181;
  assign popcount32_cdyi_core_196 = popcount32_cdyi_core_194 ^ popcount32_cdyi_core_193;
  assign popcount32_cdyi_core_197 = popcount32_cdyi_core_194 & popcount32_cdyi_core_193;
  assign popcount32_cdyi_core_198 = popcount32_cdyi_core_195 | popcount32_cdyi_core_197;
  assign popcount32_cdyi_core_200 = input_a[12] | input_a[25];
  assign popcount32_cdyi_core_203 = input_a[10] ^ input_a[5];
  assign popcount32_cdyi_core_204 = ~input_a[6];
  assign popcount32_cdyi_core_206 = popcount32_cdyi_core_106 ^ popcount32_cdyi_core_191;
  assign popcount32_cdyi_core_208 = ~popcount32_cdyi_core_206;
  assign popcount32_cdyi_core_210 = popcount32_cdyi_core_106 | popcount32_cdyi_core_206;
  assign popcount32_cdyi_core_211 = popcount32_cdyi_core_111 ^ popcount32_cdyi_core_196;
  assign popcount32_cdyi_core_212 = popcount32_cdyi_core_111 & popcount32_cdyi_core_196;
  assign popcount32_cdyi_core_213 = popcount32_cdyi_core_211 ^ popcount32_cdyi_core_210;
  assign popcount32_cdyi_core_214 = popcount32_cdyi_core_211 & popcount32_cdyi_core_210;
  assign popcount32_cdyi_core_215 = popcount32_cdyi_core_212 | popcount32_cdyi_core_214;
  assign popcount32_cdyi_core_216 = popcount32_cdyi_core_113 ^ popcount32_cdyi_core_198;
  assign popcount32_cdyi_core_217 = popcount32_cdyi_core_113 & popcount32_cdyi_core_198;
  assign popcount32_cdyi_core_218 = popcount32_cdyi_core_216 ^ popcount32_cdyi_core_215;
  assign popcount32_cdyi_core_219 = popcount32_cdyi_core_216 & popcount32_cdyi_core_215;
  assign popcount32_cdyi_core_220 = popcount32_cdyi_core_217 | popcount32_cdyi_core_219;
  assign popcount32_cdyi_core_222 = input_a[22] & input_a[2];
  assign popcount32_cdyi_core_224 = ~input_a[30];

  assign popcount32_cdyi_out[0] = popcount32_cdyi_core_218;
  assign popcount32_cdyi_out[1] = popcount32_cdyi_core_208;
  assign popcount32_cdyi_out[2] = popcount32_cdyi_core_213;
  assign popcount32_cdyi_out[3] = popcount32_cdyi_core_218;
  assign popcount32_cdyi_out[4] = popcount32_cdyi_core_220;
  assign popcount32_cdyi_out[5] = 1'b0;
endmodule