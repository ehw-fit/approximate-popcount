// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.70029
// WCE=20.0
// EP=0.884273%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_d0i1(input [37:0] input_a, output [5:0] popcount38_d0i1_out);
  wire popcount38_d0i1_core_041;
  wire popcount38_d0i1_core_044_not;
  wire popcount38_d0i1_core_045;
  wire popcount38_d0i1_core_047;
  wire popcount38_d0i1_core_049;
  wire popcount38_d0i1_core_051;
  wire popcount38_d0i1_core_052;
  wire popcount38_d0i1_core_054;
  wire popcount38_d0i1_core_055;
  wire popcount38_d0i1_core_056;
  wire popcount38_d0i1_core_057;
  wire popcount38_d0i1_core_058;
  wire popcount38_d0i1_core_059;
  wire popcount38_d0i1_core_060;
  wire popcount38_d0i1_core_062;
  wire popcount38_d0i1_core_063;
  wire popcount38_d0i1_core_064;
  wire popcount38_d0i1_core_065;
  wire popcount38_d0i1_core_067;
  wire popcount38_d0i1_core_069;
  wire popcount38_d0i1_core_070;
  wire popcount38_d0i1_core_071;
  wire popcount38_d0i1_core_072;
  wire popcount38_d0i1_core_073;
  wire popcount38_d0i1_core_075;
  wire popcount38_d0i1_core_077;
  wire popcount38_d0i1_core_079;
  wire popcount38_d0i1_core_080;
  wire popcount38_d0i1_core_082;
  wire popcount38_d0i1_core_083;
  wire popcount38_d0i1_core_086;
  wire popcount38_d0i1_core_087;
  wire popcount38_d0i1_core_088;
  wire popcount38_d0i1_core_089;
  wire popcount38_d0i1_core_090;
  wire popcount38_d0i1_core_091;
  wire popcount38_d0i1_core_094;
  wire popcount38_d0i1_core_097;
  wire popcount38_d0i1_core_098;
  wire popcount38_d0i1_core_099;
  wire popcount38_d0i1_core_100;
  wire popcount38_d0i1_core_101;
  wire popcount38_d0i1_core_104;
  wire popcount38_d0i1_core_105;
  wire popcount38_d0i1_core_106;
  wire popcount38_d0i1_core_107;
  wire popcount38_d0i1_core_108;
  wire popcount38_d0i1_core_110;
  wire popcount38_d0i1_core_112;
  wire popcount38_d0i1_core_113;
  wire popcount38_d0i1_core_115;
  wire popcount38_d0i1_core_116;
  wire popcount38_d0i1_core_119;
  wire popcount38_d0i1_core_121;
  wire popcount38_d0i1_core_122;
  wire popcount38_d0i1_core_123;
  wire popcount38_d0i1_core_124;
  wire popcount38_d0i1_core_125;
  wire popcount38_d0i1_core_131_not;
  wire popcount38_d0i1_core_133;
  wire popcount38_d0i1_core_134;
  wire popcount38_d0i1_core_135;
  wire popcount38_d0i1_core_137;
  wire popcount38_d0i1_core_140;
  wire popcount38_d0i1_core_142;
  wire popcount38_d0i1_core_145;
  wire popcount38_d0i1_core_147;
  wire popcount38_d0i1_core_148;
  wire popcount38_d0i1_core_149;
  wire popcount38_d0i1_core_150;
  wire popcount38_d0i1_core_151;
  wire popcount38_d0i1_core_153;
  wire popcount38_d0i1_core_155;
  wire popcount38_d0i1_core_156;
  wire popcount38_d0i1_core_159;
  wire popcount38_d0i1_core_162;
  wire popcount38_d0i1_core_164;
  wire popcount38_d0i1_core_165;
  wire popcount38_d0i1_core_166;
  wire popcount38_d0i1_core_168;
  wire popcount38_d0i1_core_169;
  wire popcount38_d0i1_core_170;
  wire popcount38_d0i1_core_171;
  wire popcount38_d0i1_core_172;
  wire popcount38_d0i1_core_174;
  wire popcount38_d0i1_core_175;
  wire popcount38_d0i1_core_177;
  wire popcount38_d0i1_core_178;
  wire popcount38_d0i1_core_179;
  wire popcount38_d0i1_core_180;
  wire popcount38_d0i1_core_184;
  wire popcount38_d0i1_core_185;
  wire popcount38_d0i1_core_186;
  wire popcount38_d0i1_core_190;
  wire popcount38_d0i1_core_191;
  wire popcount38_d0i1_core_193;
  wire popcount38_d0i1_core_194_not;
  wire popcount38_d0i1_core_196;
  wire popcount38_d0i1_core_197;
  wire popcount38_d0i1_core_198;
  wire popcount38_d0i1_core_200;
  wire popcount38_d0i1_core_202;
  wire popcount38_d0i1_core_203;
  wire popcount38_d0i1_core_204;
  wire popcount38_d0i1_core_205;
  wire popcount38_d0i1_core_206_not;
  wire popcount38_d0i1_core_209;
  wire popcount38_d0i1_core_211;
  wire popcount38_d0i1_core_212;
  wire popcount38_d0i1_core_213;
  wire popcount38_d0i1_core_215;
  wire popcount38_d0i1_core_216;
  wire popcount38_d0i1_core_217;
  wire popcount38_d0i1_core_218;
  wire popcount38_d0i1_core_219;
  wire popcount38_d0i1_core_221;
  wire popcount38_d0i1_core_222;
  wire popcount38_d0i1_core_223;
  wire popcount38_d0i1_core_224;
  wire popcount38_d0i1_core_225;
  wire popcount38_d0i1_core_227;
  wire popcount38_d0i1_core_228;
  wire popcount38_d0i1_core_229;
  wire popcount38_d0i1_core_230;
  wire popcount38_d0i1_core_231;
  wire popcount38_d0i1_core_232;
  wire popcount38_d0i1_core_233;
  wire popcount38_d0i1_core_234;
  wire popcount38_d0i1_core_239;
  wire popcount38_d0i1_core_241;
  wire popcount38_d0i1_core_242;
  wire popcount38_d0i1_core_243;
  wire popcount38_d0i1_core_246;
  wire popcount38_d0i1_core_247;
  wire popcount38_d0i1_core_248_not;
  wire popcount38_d0i1_core_249;
  wire popcount38_d0i1_core_251;
  wire popcount38_d0i1_core_252;
  wire popcount38_d0i1_core_253;
  wire popcount38_d0i1_core_256;
  wire popcount38_d0i1_core_257;
  wire popcount38_d0i1_core_258;
  wire popcount38_d0i1_core_259;
  wire popcount38_d0i1_core_260;
  wire popcount38_d0i1_core_261;
  wire popcount38_d0i1_core_264;
  wire popcount38_d0i1_core_265;
  wire popcount38_d0i1_core_267;
  wire popcount38_d0i1_core_268;
  wire popcount38_d0i1_core_269;
  wire popcount38_d0i1_core_270;
  wire popcount38_d0i1_core_271;
  wire popcount38_d0i1_core_272;
  wire popcount38_d0i1_core_273;
  wire popcount38_d0i1_core_277;
  wire popcount38_d0i1_core_278;
  wire popcount38_d0i1_core_279;
  wire popcount38_d0i1_core_281;
  wire popcount38_d0i1_core_282;
  wire popcount38_d0i1_core_284;
  wire popcount38_d0i1_core_286;
  wire popcount38_d0i1_core_288_not;
  wire popcount38_d0i1_core_289;
  wire popcount38_d0i1_core_293;
  wire popcount38_d0i1_core_294;
  wire popcount38_d0i1_core_295;
  wire popcount38_d0i1_core_296;

  assign popcount38_d0i1_core_041 = input_a[33] & input_a[22];
  assign popcount38_d0i1_core_044_not = ~input_a[18];
  assign popcount38_d0i1_core_045 = input_a[30] & input_a[33];
  assign popcount38_d0i1_core_047 = ~input_a[12];
  assign popcount38_d0i1_core_049 = ~(input_a[8] & input_a[5]);
  assign popcount38_d0i1_core_051 = ~(input_a[16] | input_a[33]);
  assign popcount38_d0i1_core_052 = input_a[8] | input_a[3];
  assign popcount38_d0i1_core_054 = input_a[26] | input_a[37];
  assign popcount38_d0i1_core_055 = ~(input_a[29] | input_a[4]);
  assign popcount38_d0i1_core_056 = input_a[14] | input_a[17];
  assign popcount38_d0i1_core_057 = ~input_a[29];
  assign popcount38_d0i1_core_058 = input_a[7] & input_a[16];
  assign popcount38_d0i1_core_059 = ~input_a[9];
  assign popcount38_d0i1_core_060 = ~(input_a[16] & input_a[24]);
  assign popcount38_d0i1_core_062 = ~(input_a[31] | input_a[1]);
  assign popcount38_d0i1_core_063 = ~(input_a[21] & input_a[22]);
  assign popcount38_d0i1_core_064 = ~(input_a[11] ^ input_a[2]);
  assign popcount38_d0i1_core_065 = input_a[19] | input_a[12];
  assign popcount38_d0i1_core_067 = ~(input_a[5] | input_a[36]);
  assign popcount38_d0i1_core_069 = ~(input_a[30] & input_a[31]);
  assign popcount38_d0i1_core_070 = input_a[1] ^ input_a[36];
  assign popcount38_d0i1_core_071 = ~input_a[12];
  assign popcount38_d0i1_core_072 = ~input_a[28];
  assign popcount38_d0i1_core_073 = input_a[29] | input_a[29];
  assign popcount38_d0i1_core_075 = input_a[18] & input_a[4];
  assign popcount38_d0i1_core_077 = ~(input_a[1] ^ input_a[7]);
  assign popcount38_d0i1_core_079 = input_a[20] ^ input_a[32];
  assign popcount38_d0i1_core_080 = input_a[15] ^ input_a[15];
  assign popcount38_d0i1_core_082 = ~(input_a[11] | input_a[23]);
  assign popcount38_d0i1_core_083 = ~(input_a[6] & input_a[5]);
  assign popcount38_d0i1_core_086 = input_a[21] | input_a[37];
  assign popcount38_d0i1_core_087 = input_a[24] ^ input_a[9];
  assign popcount38_d0i1_core_088 = ~input_a[15];
  assign popcount38_d0i1_core_089 = ~(input_a[23] ^ input_a[10]);
  assign popcount38_d0i1_core_090 = ~(input_a[12] & input_a[19]);
  assign popcount38_d0i1_core_091 = input_a[14] & input_a[13];
  assign popcount38_d0i1_core_094 = ~(input_a[30] ^ input_a[7]);
  assign popcount38_d0i1_core_097 = input_a[16] ^ input_a[30];
  assign popcount38_d0i1_core_098 = input_a[3] | input_a[17];
  assign popcount38_d0i1_core_099 = input_a[20] | input_a[12];
  assign popcount38_d0i1_core_100 = ~input_a[30];
  assign popcount38_d0i1_core_101 = ~(input_a[12] | input_a[27]);
  assign popcount38_d0i1_core_104 = input_a[36] & input_a[21];
  assign popcount38_d0i1_core_105 = input_a[18] ^ input_a[23];
  assign popcount38_d0i1_core_106 = input_a[14] | input_a[31];
  assign popcount38_d0i1_core_107 = ~(input_a[34] | input_a[27]);
  assign popcount38_d0i1_core_108 = ~(input_a[35] & input_a[24]);
  assign popcount38_d0i1_core_110 = input_a[32] ^ input_a[16];
  assign popcount38_d0i1_core_112 = input_a[33] ^ input_a[33];
  assign popcount38_d0i1_core_113 = input_a[5] & input_a[1];
  assign popcount38_d0i1_core_115 = input_a[11] & input_a[19];
  assign popcount38_d0i1_core_116 = ~(input_a[34] ^ input_a[18]);
  assign popcount38_d0i1_core_119 = ~(input_a[13] | input_a[14]);
  assign popcount38_d0i1_core_121 = input_a[25] & input_a[32];
  assign popcount38_d0i1_core_122 = ~(input_a[16] & input_a[29]);
  assign popcount38_d0i1_core_123 = input_a[16] & input_a[16];
  assign popcount38_d0i1_core_124 = ~input_a[21];
  assign popcount38_d0i1_core_125 = input_a[2] ^ input_a[18];
  assign popcount38_d0i1_core_131_not = ~input_a[17];
  assign popcount38_d0i1_core_133 = ~(input_a[7] & input_a[23]);
  assign popcount38_d0i1_core_134 = input_a[34] & input_a[2];
  assign popcount38_d0i1_core_135 = ~(input_a[29] & input_a[26]);
  assign popcount38_d0i1_core_137 = ~(input_a[28] ^ input_a[37]);
  assign popcount38_d0i1_core_140 = input_a[14] | input_a[5];
  assign popcount38_d0i1_core_142 = ~input_a[25];
  assign popcount38_d0i1_core_145 = input_a[20] & input_a[21];
  assign popcount38_d0i1_core_147 = ~(input_a[1] | input_a[3]);
  assign popcount38_d0i1_core_148 = input_a[33] ^ input_a[29];
  assign popcount38_d0i1_core_149 = input_a[3] ^ input_a[13];
  assign popcount38_d0i1_core_150 = ~(input_a[21] ^ input_a[37]);
  assign popcount38_d0i1_core_151 = input_a[3] & input_a[17];
  assign popcount38_d0i1_core_153 = ~(input_a[34] ^ input_a[17]);
  assign popcount38_d0i1_core_155 = input_a[23] | input_a[18];
  assign popcount38_d0i1_core_156 = ~(input_a[4] | input_a[33]);
  assign popcount38_d0i1_core_159 = ~input_a[8];
  assign popcount38_d0i1_core_162 = ~(input_a[32] ^ input_a[9]);
  assign popcount38_d0i1_core_164 = ~input_a[16];
  assign popcount38_d0i1_core_165 = input_a[12] ^ input_a[11];
  assign popcount38_d0i1_core_166 = ~(input_a[22] & input_a[4]);
  assign popcount38_d0i1_core_168 = input_a[2] & input_a[26];
  assign popcount38_d0i1_core_169 = ~input_a[6];
  assign popcount38_d0i1_core_170 = input_a[32] ^ input_a[37];
  assign popcount38_d0i1_core_171 = ~input_a[11];
  assign popcount38_d0i1_core_172 = input_a[23] | input_a[5];
  assign popcount38_d0i1_core_174 = ~(input_a[33] & input_a[3]);
  assign popcount38_d0i1_core_175 = input_a[2] & input_a[13];
  assign popcount38_d0i1_core_177 = input_a[33] & input_a[23];
  assign popcount38_d0i1_core_178 = input_a[12] ^ input_a[19];
  assign popcount38_d0i1_core_179 = input_a[28] | input_a[30];
  assign popcount38_d0i1_core_180 = ~input_a[15];
  assign popcount38_d0i1_core_184 = input_a[5] & input_a[6];
  assign popcount38_d0i1_core_185 = input_a[30] ^ input_a[2];
  assign popcount38_d0i1_core_186 = input_a[5] ^ input_a[9];
  assign popcount38_d0i1_core_190 = input_a[0] | input_a[21];
  assign popcount38_d0i1_core_191 = input_a[30] | input_a[2];
  assign popcount38_d0i1_core_193 = ~(input_a[24] | input_a[6]);
  assign popcount38_d0i1_core_194_not = ~input_a[16];
  assign popcount38_d0i1_core_196 = input_a[8] | input_a[2];
  assign popcount38_d0i1_core_197 = input_a[8] ^ input_a[6];
  assign popcount38_d0i1_core_198 = ~input_a[9];
  assign popcount38_d0i1_core_200 = input_a[26] | input_a[10];
  assign popcount38_d0i1_core_202 = ~(input_a[2] & input_a[25]);
  assign popcount38_d0i1_core_203 = input_a[18] | input_a[34];
  assign popcount38_d0i1_core_204 = ~(input_a[18] & input_a[31]);
  assign popcount38_d0i1_core_205 = ~(input_a[26] & input_a[17]);
  assign popcount38_d0i1_core_206_not = ~input_a[37];
  assign popcount38_d0i1_core_209 = input_a[28] | input_a[8];
  assign popcount38_d0i1_core_211 = input_a[3] | input_a[27];
  assign popcount38_d0i1_core_212 = ~input_a[32];
  assign popcount38_d0i1_core_213 = input_a[17] ^ input_a[22];
  assign popcount38_d0i1_core_215 = ~(input_a[1] & input_a[22]);
  assign popcount38_d0i1_core_216 = input_a[10] ^ input_a[25];
  assign popcount38_d0i1_core_217 = ~input_a[27];
  assign popcount38_d0i1_core_218 = input_a[28] | input_a[18];
  assign popcount38_d0i1_core_219 = ~(input_a[31] | input_a[3]);
  assign popcount38_d0i1_core_221 = input_a[11] & input_a[11];
  assign popcount38_d0i1_core_222 = ~(input_a[21] & input_a[2]);
  assign popcount38_d0i1_core_223 = ~(input_a[17] ^ input_a[27]);
  assign popcount38_d0i1_core_224 = input_a[5] | input_a[19];
  assign popcount38_d0i1_core_225 = input_a[20] | input_a[26];
  assign popcount38_d0i1_core_227 = input_a[34] & input_a[34];
  assign popcount38_d0i1_core_228 = ~input_a[30];
  assign popcount38_d0i1_core_229 = ~input_a[21];
  assign popcount38_d0i1_core_230 = input_a[1] ^ input_a[7];
  assign popcount38_d0i1_core_231 = ~(input_a[0] & input_a[18]);
  assign popcount38_d0i1_core_232 = input_a[24] | input_a[19];
  assign popcount38_d0i1_core_233 = ~(input_a[20] | input_a[17]);
  assign popcount38_d0i1_core_234 = ~input_a[6];
  assign popcount38_d0i1_core_239 = ~input_a[17];
  assign popcount38_d0i1_core_241 = ~(input_a[17] & input_a[0]);
  assign popcount38_d0i1_core_242 = input_a[25] & input_a[37];
  assign popcount38_d0i1_core_243 = ~input_a[11];
  assign popcount38_d0i1_core_246 = input_a[31] & input_a[17];
  assign popcount38_d0i1_core_247 = ~(input_a[27] & input_a[30]);
  assign popcount38_d0i1_core_248_not = ~input_a[20];
  assign popcount38_d0i1_core_249 = input_a[13] & input_a[27];
  assign popcount38_d0i1_core_251 = input_a[33] ^ input_a[28];
  assign popcount38_d0i1_core_252 = ~(input_a[31] | input_a[32]);
  assign popcount38_d0i1_core_253 = input_a[24] | input_a[2];
  assign popcount38_d0i1_core_256 = input_a[3] | input_a[20];
  assign popcount38_d0i1_core_257 = ~(input_a[20] ^ input_a[25]);
  assign popcount38_d0i1_core_258 = ~input_a[31];
  assign popcount38_d0i1_core_259 = ~(input_a[26] & input_a[12]);
  assign popcount38_d0i1_core_260 = ~(input_a[14] ^ input_a[5]);
  assign popcount38_d0i1_core_261 = input_a[17] | input_a[27];
  assign popcount38_d0i1_core_264 = ~(input_a[37] & input_a[26]);
  assign popcount38_d0i1_core_265 = input_a[14] & input_a[13];
  assign popcount38_d0i1_core_267 = input_a[29] | input_a[16];
  assign popcount38_d0i1_core_268 = ~(input_a[3] | input_a[13]);
  assign popcount38_d0i1_core_269 = input_a[14] ^ input_a[17];
  assign popcount38_d0i1_core_270 = ~(input_a[16] ^ input_a[37]);
  assign popcount38_d0i1_core_271 = ~(input_a[27] | input_a[18]);
  assign popcount38_d0i1_core_272 = ~input_a[2];
  assign popcount38_d0i1_core_273 = ~(input_a[21] & input_a[30]);
  assign popcount38_d0i1_core_277 = input_a[32] ^ input_a[3];
  assign popcount38_d0i1_core_278 = ~(input_a[20] ^ input_a[2]);
  assign popcount38_d0i1_core_279 = input_a[24] ^ input_a[29];
  assign popcount38_d0i1_core_281 = input_a[36] & input_a[2];
  assign popcount38_d0i1_core_282 = input_a[21] ^ input_a[15];
  assign popcount38_d0i1_core_284 = input_a[3] | input_a[12];
  assign popcount38_d0i1_core_286 = ~input_a[22];
  assign popcount38_d0i1_core_288_not = ~input_a[24];
  assign popcount38_d0i1_core_289 = input_a[37] ^ input_a[35];
  assign popcount38_d0i1_core_293 = ~input_a[25];
  assign popcount38_d0i1_core_294 = input_a[3] | input_a[11];
  assign popcount38_d0i1_core_295 = ~(input_a[21] ^ input_a[13]);
  assign popcount38_d0i1_core_296 = ~(input_a[3] | input_a[26]);

  assign popcount38_d0i1_out[0] = input_a[8];
  assign popcount38_d0i1_out[1] = input_a[28];
  assign popcount38_d0i1_out[2] = input_a[4];
  assign popcount38_d0i1_out[3] = 1'b0;
  assign popcount38_d0i1_out[4] = 1'b1;
  assign popcount38_d0i1_out[5] = 1'b0;
endmodule