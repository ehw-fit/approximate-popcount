// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.39114
// WCE=15.0
// EP=0.87048%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_7cxv(input [27:0] input_a, output [4:0] popcount28_7cxv_out);
  wire popcount28_7cxv_core_030;
  wire popcount28_7cxv_core_033;
  wire popcount28_7cxv_core_034;
  wire popcount28_7cxv_core_035;
  wire popcount28_7cxv_core_036;
  wire popcount28_7cxv_core_038;
  wire popcount28_7cxv_core_039_not;
  wire popcount28_7cxv_core_040;
  wire popcount28_7cxv_core_041;
  wire popcount28_7cxv_core_042;
  wire popcount28_7cxv_core_044;
  wire popcount28_7cxv_core_045;
  wire popcount28_7cxv_core_047;
  wire popcount28_7cxv_core_052;
  wire popcount28_7cxv_core_054;
  wire popcount28_7cxv_core_056;
  wire popcount28_7cxv_core_058;
  wire popcount28_7cxv_core_059;
  wire popcount28_7cxv_core_061;
  wire popcount28_7cxv_core_062;
  wire popcount28_7cxv_core_063;
  wire popcount28_7cxv_core_064;
  wire popcount28_7cxv_core_065;
  wire popcount28_7cxv_core_066;
  wire popcount28_7cxv_core_067;
  wire popcount28_7cxv_core_069;
  wire popcount28_7cxv_core_071;
  wire popcount28_7cxv_core_073;
  wire popcount28_7cxv_core_074;
  wire popcount28_7cxv_core_075;
  wire popcount28_7cxv_core_076;
  wire popcount28_7cxv_core_078;
  wire popcount28_7cxv_core_080;
  wire popcount28_7cxv_core_081;
  wire popcount28_7cxv_core_084;
  wire popcount28_7cxv_core_085;
  wire popcount28_7cxv_core_086;
  wire popcount28_7cxv_core_087;
  wire popcount28_7cxv_core_088;
  wire popcount28_7cxv_core_089;
  wire popcount28_7cxv_core_090_not;
  wire popcount28_7cxv_core_091;
  wire popcount28_7cxv_core_092;
  wire popcount28_7cxv_core_094;
  wire popcount28_7cxv_core_095;
  wire popcount28_7cxv_core_096;
  wire popcount28_7cxv_core_098_not;
  wire popcount28_7cxv_core_099;
  wire popcount28_7cxv_core_100;
  wire popcount28_7cxv_core_102;
  wire popcount28_7cxv_core_104;
  wire popcount28_7cxv_core_105;
  wire popcount28_7cxv_core_106;
  wire popcount28_7cxv_core_107;
  wire popcount28_7cxv_core_111_not;
  wire popcount28_7cxv_core_112;
  wire popcount28_7cxv_core_113;
  wire popcount28_7cxv_core_114;
  wire popcount28_7cxv_core_115;
  wire popcount28_7cxv_core_116;
  wire popcount28_7cxv_core_117;
  wire popcount28_7cxv_core_118;
  wire popcount28_7cxv_core_120;
  wire popcount28_7cxv_core_121;
  wire popcount28_7cxv_core_123;
  wire popcount28_7cxv_core_125;
  wire popcount28_7cxv_core_126;
  wire popcount28_7cxv_core_128;
  wire popcount28_7cxv_core_130;
  wire popcount28_7cxv_core_134;
  wire popcount28_7cxv_core_135;
  wire popcount28_7cxv_core_137;
  wire popcount28_7cxv_core_138;
  wire popcount28_7cxv_core_139;
  wire popcount28_7cxv_core_140;
  wire popcount28_7cxv_core_141;
  wire popcount28_7cxv_core_142;
  wire popcount28_7cxv_core_143;
  wire popcount28_7cxv_core_144;
  wire popcount28_7cxv_core_145;
  wire popcount28_7cxv_core_146;
  wire popcount28_7cxv_core_151;
  wire popcount28_7cxv_core_152;
  wire popcount28_7cxv_core_154;
  wire popcount28_7cxv_core_155;
  wire popcount28_7cxv_core_156;
  wire popcount28_7cxv_core_157;
  wire popcount28_7cxv_core_158;
  wire popcount28_7cxv_core_159;
  wire popcount28_7cxv_core_160;
  wire popcount28_7cxv_core_162;
  wire popcount28_7cxv_core_164;
  wire popcount28_7cxv_core_169;
  wire popcount28_7cxv_core_170;
  wire popcount28_7cxv_core_171;
  wire popcount28_7cxv_core_172;
  wire popcount28_7cxv_core_173;
  wire popcount28_7cxv_core_174;
  wire popcount28_7cxv_core_176;
  wire popcount28_7cxv_core_177_not;
  wire popcount28_7cxv_core_178;
  wire popcount28_7cxv_core_179;
  wire popcount28_7cxv_core_180;
  wire popcount28_7cxv_core_182;
  wire popcount28_7cxv_core_185;
  wire popcount28_7cxv_core_186;
  wire popcount28_7cxv_core_188;
  wire popcount28_7cxv_core_189;
  wire popcount28_7cxv_core_190;
  wire popcount28_7cxv_core_191;
  wire popcount28_7cxv_core_193;
  wire popcount28_7cxv_core_195;
  wire popcount28_7cxv_core_197;
  wire popcount28_7cxv_core_198;

  assign popcount28_7cxv_core_030 = ~(input_a[7] | input_a[23]);
  assign popcount28_7cxv_core_033 = ~(input_a[20] | input_a[17]);
  assign popcount28_7cxv_core_034 = input_a[8] ^ input_a[8];
  assign popcount28_7cxv_core_035 = input_a[19] & input_a[6];
  assign popcount28_7cxv_core_036 = input_a[14] ^ input_a[26];
  assign popcount28_7cxv_core_038 = ~(input_a[24] & input_a[20]);
  assign popcount28_7cxv_core_039_not = ~input_a[12];
  assign popcount28_7cxv_core_040 = ~input_a[18];
  assign popcount28_7cxv_core_041 = ~(input_a[9] ^ input_a[25]);
  assign popcount28_7cxv_core_042 = ~(input_a[20] | input_a[18]);
  assign popcount28_7cxv_core_044 = input_a[6] | input_a[1];
  assign popcount28_7cxv_core_045 = input_a[27] & input_a[10];
  assign popcount28_7cxv_core_047 = ~input_a[8];
  assign popcount28_7cxv_core_052 = input_a[12] & input_a[22];
  assign popcount28_7cxv_core_054 = ~(input_a[7] | input_a[26]);
  assign popcount28_7cxv_core_056 = input_a[1] ^ input_a[20];
  assign popcount28_7cxv_core_058 = ~(input_a[20] | input_a[21]);
  assign popcount28_7cxv_core_059 = input_a[15] | input_a[9];
  assign popcount28_7cxv_core_061 = ~input_a[8];
  assign popcount28_7cxv_core_062 = input_a[20] & input_a[0];
  assign popcount28_7cxv_core_063 = input_a[22] | input_a[5];
  assign popcount28_7cxv_core_064 = input_a[18] | input_a[16];
  assign popcount28_7cxv_core_065 = ~(input_a[4] ^ input_a[17]);
  assign popcount28_7cxv_core_066 = input_a[26] | input_a[9];
  assign popcount28_7cxv_core_067 = input_a[25] & input_a[1];
  assign popcount28_7cxv_core_069 = ~(input_a[16] & input_a[7]);
  assign popcount28_7cxv_core_071 = input_a[0] | input_a[1];
  assign popcount28_7cxv_core_073 = ~(input_a[15] | input_a[24]);
  assign popcount28_7cxv_core_074 = ~input_a[22];
  assign popcount28_7cxv_core_075 = input_a[25] & input_a[9];
  assign popcount28_7cxv_core_076 = ~(input_a[15] | input_a[18]);
  assign popcount28_7cxv_core_078 = input_a[0] ^ input_a[13];
  assign popcount28_7cxv_core_080 = input_a[1] & input_a[22];
  assign popcount28_7cxv_core_081 = ~input_a[1];
  assign popcount28_7cxv_core_084 = input_a[17] ^ input_a[0];
  assign popcount28_7cxv_core_085 = input_a[1] & input_a[15];
  assign popcount28_7cxv_core_086 = ~(input_a[25] & input_a[0]);
  assign popcount28_7cxv_core_087 = input_a[6] ^ input_a[25];
  assign popcount28_7cxv_core_088 = ~input_a[23];
  assign popcount28_7cxv_core_089 = input_a[26] | input_a[15];
  assign popcount28_7cxv_core_090_not = ~input_a[11];
  assign popcount28_7cxv_core_091 = input_a[1] ^ input_a[14];
  assign popcount28_7cxv_core_092 = input_a[15] & input_a[22];
  assign popcount28_7cxv_core_094 = ~(input_a[1] ^ input_a[15]);
  assign popcount28_7cxv_core_095 = input_a[5] | input_a[25];
  assign popcount28_7cxv_core_096 = input_a[11] | input_a[23];
  assign popcount28_7cxv_core_098_not = ~input_a[6];
  assign popcount28_7cxv_core_099 = input_a[5] & input_a[25];
  assign popcount28_7cxv_core_100 = ~(input_a[23] | input_a[0]);
  assign popcount28_7cxv_core_102 = ~(input_a[9] & input_a[0]);
  assign popcount28_7cxv_core_104 = input_a[8] & input_a[17];
  assign popcount28_7cxv_core_105 = input_a[0] ^ input_a[24];
  assign popcount28_7cxv_core_106 = ~(input_a[11] | input_a[5]);
  assign popcount28_7cxv_core_107 = ~(input_a[16] | input_a[9]);
  assign popcount28_7cxv_core_111_not = ~input_a[8];
  assign popcount28_7cxv_core_112 = ~(input_a[26] ^ input_a[8]);
  assign popcount28_7cxv_core_113 = ~(input_a[27] & input_a[14]);
  assign popcount28_7cxv_core_114 = input_a[7] | input_a[26];
  assign popcount28_7cxv_core_115 = input_a[8] ^ input_a[0];
  assign popcount28_7cxv_core_116 = input_a[0] ^ input_a[13];
  assign popcount28_7cxv_core_117 = input_a[27] & input_a[21];
  assign popcount28_7cxv_core_118 = input_a[9] ^ input_a[23];
  assign popcount28_7cxv_core_120 = ~(input_a[14] | input_a[11]);
  assign popcount28_7cxv_core_121 = input_a[9] & input_a[13];
  assign popcount28_7cxv_core_123 = ~(input_a[9] ^ input_a[3]);
  assign popcount28_7cxv_core_125 = input_a[14] & input_a[20];
  assign popcount28_7cxv_core_126 = input_a[18] & input_a[22];
  assign popcount28_7cxv_core_128 = ~input_a[7];
  assign popcount28_7cxv_core_130 = input_a[8] | input_a[1];
  assign popcount28_7cxv_core_134 = ~(input_a[22] ^ input_a[9]);
  assign popcount28_7cxv_core_135 = input_a[3] & input_a[13];
  assign popcount28_7cxv_core_137 = ~(input_a[26] ^ input_a[12]);
  assign popcount28_7cxv_core_138 = input_a[9] | input_a[3];
  assign popcount28_7cxv_core_139 = ~(input_a[8] | input_a[0]);
  assign popcount28_7cxv_core_140 = input_a[0] ^ input_a[23];
  assign popcount28_7cxv_core_141 = ~input_a[11];
  assign popcount28_7cxv_core_142 = input_a[22] & input_a[8];
  assign popcount28_7cxv_core_143 = ~(input_a[4] | input_a[5]);
  assign popcount28_7cxv_core_144 = ~(input_a[3] & input_a[14]);
  assign popcount28_7cxv_core_145 = input_a[27] | input_a[9];
  assign popcount28_7cxv_core_146 = input_a[12] ^ input_a[25];
  assign popcount28_7cxv_core_151 = input_a[6] ^ input_a[14];
  assign popcount28_7cxv_core_152 = input_a[25] | input_a[13];
  assign popcount28_7cxv_core_154 = ~(input_a[1] & input_a[1]);
  assign popcount28_7cxv_core_155 = input_a[1] | input_a[17];
  assign popcount28_7cxv_core_156 = ~(input_a[17] | input_a[26]);
  assign popcount28_7cxv_core_157 = ~(input_a[25] ^ input_a[21]);
  assign popcount28_7cxv_core_158 = input_a[5] ^ input_a[19];
  assign popcount28_7cxv_core_159 = ~(input_a[15] | input_a[18]);
  assign popcount28_7cxv_core_160 = input_a[10] ^ input_a[9];
  assign popcount28_7cxv_core_162 = input_a[9] & input_a[17];
  assign popcount28_7cxv_core_164 = ~(input_a[12] ^ input_a[16]);
  assign popcount28_7cxv_core_169 = ~(input_a[2] & input_a[26]);
  assign popcount28_7cxv_core_170 = input_a[17] ^ input_a[24];
  assign popcount28_7cxv_core_171 = ~(input_a[7] | input_a[21]);
  assign popcount28_7cxv_core_172 = ~(input_a[15] & input_a[4]);
  assign popcount28_7cxv_core_173 = ~(input_a[18] & input_a[21]);
  assign popcount28_7cxv_core_174 = ~(input_a[10] | input_a[6]);
  assign popcount28_7cxv_core_176 = ~(input_a[13] & input_a[13]);
  assign popcount28_7cxv_core_177_not = ~input_a[5];
  assign popcount28_7cxv_core_178 = ~(input_a[12] | input_a[24]);
  assign popcount28_7cxv_core_179 = ~(input_a[25] & input_a[0]);
  assign popcount28_7cxv_core_180 = input_a[5] | input_a[8];
  assign popcount28_7cxv_core_182 = ~input_a[20];
  assign popcount28_7cxv_core_185 = input_a[10] & input_a[24];
  assign popcount28_7cxv_core_186 = ~input_a[13];
  assign popcount28_7cxv_core_188 = input_a[3] & input_a[14];
  assign popcount28_7cxv_core_189 = ~(input_a[25] & input_a[1]);
  assign popcount28_7cxv_core_190 = input_a[25] ^ input_a[2];
  assign popcount28_7cxv_core_191 = input_a[3] ^ input_a[10];
  assign popcount28_7cxv_core_193 = ~(input_a[21] | input_a[18]);
  assign popcount28_7cxv_core_195 = input_a[17] ^ input_a[27];
  assign popcount28_7cxv_core_197 = input_a[4] & input_a[12];
  assign popcount28_7cxv_core_198 = input_a[6] ^ input_a[25];

  assign popcount28_7cxv_out[0] = input_a[18];
  assign popcount28_7cxv_out[1] = 1'b0;
  assign popcount28_7cxv_out[2] = 1'b1;
  assign popcount28_7cxv_out[3] = 1'b1;
  assign popcount28_7cxv_out[4] = 1'b0;
endmodule