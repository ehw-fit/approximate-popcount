// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.07986
// WCE=29.0
// EP=0.949195%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_lhas(input [38:0] input_a, output [5:0] popcount39_lhas_out);
  wire popcount39_lhas_core_042;
  wire popcount39_lhas_core_043;
  wire popcount39_lhas_core_045;
  wire popcount39_lhas_core_046;
  wire popcount39_lhas_core_047;
  wire popcount39_lhas_core_048;
  wire popcount39_lhas_core_049;
  wire popcount39_lhas_core_051;
  wire popcount39_lhas_core_054;
  wire popcount39_lhas_core_056;
  wire popcount39_lhas_core_058;
  wire popcount39_lhas_core_059;
  wire popcount39_lhas_core_060;
  wire popcount39_lhas_core_061_not;
  wire popcount39_lhas_core_062;
  wire popcount39_lhas_core_063;
  wire popcount39_lhas_core_064;
  wire popcount39_lhas_core_065;
  wire popcount39_lhas_core_066_not;
  wire popcount39_lhas_core_067;
  wire popcount39_lhas_core_069;
  wire popcount39_lhas_core_070;
  wire popcount39_lhas_core_071;
  wire popcount39_lhas_core_072;
  wire popcount39_lhas_core_073;
  wire popcount39_lhas_core_074;
  wire popcount39_lhas_core_076;
  wire popcount39_lhas_core_077;
  wire popcount39_lhas_core_078;
  wire popcount39_lhas_core_079;
  wire popcount39_lhas_core_080;
  wire popcount39_lhas_core_082;
  wire popcount39_lhas_core_083;
  wire popcount39_lhas_core_085;
  wire popcount39_lhas_core_086;
  wire popcount39_lhas_core_089;
  wire popcount39_lhas_core_090;
  wire popcount39_lhas_core_092;
  wire popcount39_lhas_core_093;
  wire popcount39_lhas_core_094_not;
  wire popcount39_lhas_core_095;
  wire popcount39_lhas_core_099;
  wire popcount39_lhas_core_100;
  wire popcount39_lhas_core_101;
  wire popcount39_lhas_core_102;
  wire popcount39_lhas_core_105;
  wire popcount39_lhas_core_106;
  wire popcount39_lhas_core_107;
  wire popcount39_lhas_core_108;
  wire popcount39_lhas_core_109;
  wire popcount39_lhas_core_110;
  wire popcount39_lhas_core_111;
  wire popcount39_lhas_core_112;
  wire popcount39_lhas_core_114;
  wire popcount39_lhas_core_116;
  wire popcount39_lhas_core_117;
  wire popcount39_lhas_core_118;
  wire popcount39_lhas_core_119;
  wire popcount39_lhas_core_120;
  wire popcount39_lhas_core_121;
  wire popcount39_lhas_core_123;
  wire popcount39_lhas_core_124_not;
  wire popcount39_lhas_core_125;
  wire popcount39_lhas_core_126;
  wire popcount39_lhas_core_127;
  wire popcount39_lhas_core_129;
  wire popcount39_lhas_core_130;
  wire popcount39_lhas_core_131;
  wire popcount39_lhas_core_135;
  wire popcount39_lhas_core_136;
  wire popcount39_lhas_core_137;
  wire popcount39_lhas_core_138;
  wire popcount39_lhas_core_139;
  wire popcount39_lhas_core_140;
  wire popcount39_lhas_core_141;
  wire popcount39_lhas_core_144_not;
  wire popcount39_lhas_core_147;
  wire popcount39_lhas_core_150;
  wire popcount39_lhas_core_151;
  wire popcount39_lhas_core_152;
  wire popcount39_lhas_core_153;
  wire popcount39_lhas_core_156;
  wire popcount39_lhas_core_157;
  wire popcount39_lhas_core_158;
  wire popcount39_lhas_core_160;
  wire popcount39_lhas_core_162;
  wire popcount39_lhas_core_163;
  wire popcount39_lhas_core_166;
  wire popcount39_lhas_core_167;
  wire popcount39_lhas_core_168;
  wire popcount39_lhas_core_169;
  wire popcount39_lhas_core_172;
  wire popcount39_lhas_core_174;
  wire popcount39_lhas_core_177;
  wire popcount39_lhas_core_178;
  wire popcount39_lhas_core_179;
  wire popcount39_lhas_core_180;
  wire popcount39_lhas_core_181;
  wire popcount39_lhas_core_182;
  wire popcount39_lhas_core_183;
  wire popcount39_lhas_core_184;
  wire popcount39_lhas_core_185;
  wire popcount39_lhas_core_187;
  wire popcount39_lhas_core_188;
  wire popcount39_lhas_core_189_not;
  wire popcount39_lhas_core_190;
  wire popcount39_lhas_core_192;
  wire popcount39_lhas_core_194;
  wire popcount39_lhas_core_195;
  wire popcount39_lhas_core_196;
  wire popcount39_lhas_core_197;
  wire popcount39_lhas_core_198;
  wire popcount39_lhas_core_199;
  wire popcount39_lhas_core_200;
  wire popcount39_lhas_core_201;
  wire popcount39_lhas_core_202_not;
  wire popcount39_lhas_core_203;
  wire popcount39_lhas_core_205;
  wire popcount39_lhas_core_206;
  wire popcount39_lhas_core_207;
  wire popcount39_lhas_core_208;
  wire popcount39_lhas_core_210;
  wire popcount39_lhas_core_212;
  wire popcount39_lhas_core_213_not;
  wire popcount39_lhas_core_214;
  wire popcount39_lhas_core_215;
  wire popcount39_lhas_core_216;
  wire popcount39_lhas_core_217;
  wire popcount39_lhas_core_219;
  wire popcount39_lhas_core_221;
  wire popcount39_lhas_core_224;
  wire popcount39_lhas_core_225;
  wire popcount39_lhas_core_226;
  wire popcount39_lhas_core_227;
  wire popcount39_lhas_core_228;
  wire popcount39_lhas_core_229;
  wire popcount39_lhas_core_231;
  wire popcount39_lhas_core_233;
  wire popcount39_lhas_core_234;
  wire popcount39_lhas_core_235;
  wire popcount39_lhas_core_237;
  wire popcount39_lhas_core_238;
  wire popcount39_lhas_core_241;
  wire popcount39_lhas_core_242;
  wire popcount39_lhas_core_243;
  wire popcount39_lhas_core_244;
  wire popcount39_lhas_core_246;
  wire popcount39_lhas_core_249;
  wire popcount39_lhas_core_250;
  wire popcount39_lhas_core_251;
  wire popcount39_lhas_core_253;
  wire popcount39_lhas_core_256;
  wire popcount39_lhas_core_258;
  wire popcount39_lhas_core_260;
  wire popcount39_lhas_core_262;
  wire popcount39_lhas_core_264;
  wire popcount39_lhas_core_266;
  wire popcount39_lhas_core_271;
  wire popcount39_lhas_core_272;
  wire popcount39_lhas_core_273;
  wire popcount39_lhas_core_274;
  wire popcount39_lhas_core_276;
  wire popcount39_lhas_core_277;
  wire popcount39_lhas_core_278;
  wire popcount39_lhas_core_280;
  wire popcount39_lhas_core_281;
  wire popcount39_lhas_core_285;
  wire popcount39_lhas_core_286;
  wire popcount39_lhas_core_287;
  wire popcount39_lhas_core_289;
  wire popcount39_lhas_core_292;
  wire popcount39_lhas_core_294;
  wire popcount39_lhas_core_295;
  wire popcount39_lhas_core_299;
  wire popcount39_lhas_core_300;
  wire popcount39_lhas_core_301;
  wire popcount39_lhas_core_303;
  wire popcount39_lhas_core_304;
  wire popcount39_lhas_core_306;

  assign popcount39_lhas_core_042 = ~(input_a[31] & input_a[2]);
  assign popcount39_lhas_core_043 = ~(input_a[28] & input_a[11]);
  assign popcount39_lhas_core_045 = input_a[30] & input_a[34];
  assign popcount39_lhas_core_046 = input_a[12] | input_a[18];
  assign popcount39_lhas_core_047 = input_a[29] | input_a[34];
  assign popcount39_lhas_core_048 = ~(input_a[18] | input_a[3]);
  assign popcount39_lhas_core_049 = ~(input_a[29] ^ input_a[24]);
  assign popcount39_lhas_core_051 = ~(input_a[38] | input_a[25]);
  assign popcount39_lhas_core_054 = ~(input_a[6] ^ input_a[5]);
  assign popcount39_lhas_core_056 = ~(input_a[1] ^ input_a[13]);
  assign popcount39_lhas_core_058 = ~input_a[33];
  assign popcount39_lhas_core_059 = ~(input_a[32] ^ input_a[17]);
  assign popcount39_lhas_core_060 = input_a[17] ^ input_a[17];
  assign popcount39_lhas_core_061_not = ~input_a[35];
  assign popcount39_lhas_core_062 = input_a[15] | input_a[1];
  assign popcount39_lhas_core_063 = input_a[8] ^ input_a[2];
  assign popcount39_lhas_core_064 = input_a[0] | input_a[35];
  assign popcount39_lhas_core_065 = input_a[31] | input_a[16];
  assign popcount39_lhas_core_066_not = ~input_a[17];
  assign popcount39_lhas_core_067 = input_a[25] | input_a[37];
  assign popcount39_lhas_core_069 = ~(input_a[3] ^ input_a[11]);
  assign popcount39_lhas_core_070 = ~input_a[10];
  assign popcount39_lhas_core_071 = ~(input_a[25] ^ input_a[20]);
  assign popcount39_lhas_core_072 = ~(input_a[32] | input_a[12]);
  assign popcount39_lhas_core_073 = ~(input_a[0] ^ input_a[2]);
  assign popcount39_lhas_core_074 = input_a[32] & input_a[0];
  assign popcount39_lhas_core_076 = input_a[38] ^ input_a[37];
  assign popcount39_lhas_core_077 = ~(input_a[11] | input_a[2]);
  assign popcount39_lhas_core_078 = ~(input_a[29] ^ input_a[28]);
  assign popcount39_lhas_core_079 = ~input_a[15];
  assign popcount39_lhas_core_080 = ~(input_a[20] & input_a[11]);
  assign popcount39_lhas_core_082 = ~(input_a[8] ^ input_a[22]);
  assign popcount39_lhas_core_083 = ~(input_a[6] | input_a[24]);
  assign popcount39_lhas_core_085 = input_a[33] ^ input_a[20];
  assign popcount39_lhas_core_086 = input_a[22] | input_a[31];
  assign popcount39_lhas_core_089 = ~(input_a[14] & input_a[33]);
  assign popcount39_lhas_core_090 = input_a[2] & input_a[19];
  assign popcount39_lhas_core_092 = input_a[4] | input_a[20];
  assign popcount39_lhas_core_093 = input_a[18] ^ input_a[0];
  assign popcount39_lhas_core_094_not = ~input_a[6];
  assign popcount39_lhas_core_095 = ~input_a[6];
  assign popcount39_lhas_core_099 = input_a[27] & input_a[18];
  assign popcount39_lhas_core_100 = input_a[16] | input_a[35];
  assign popcount39_lhas_core_101 = ~(input_a[4] | input_a[33]);
  assign popcount39_lhas_core_102 = ~input_a[36];
  assign popcount39_lhas_core_105 = ~(input_a[6] ^ input_a[9]);
  assign popcount39_lhas_core_106 = input_a[3] & input_a[15];
  assign popcount39_lhas_core_107 = ~(input_a[37] ^ input_a[29]);
  assign popcount39_lhas_core_108 = ~(input_a[33] | input_a[6]);
  assign popcount39_lhas_core_109 = ~input_a[34];
  assign popcount39_lhas_core_110 = ~(input_a[0] & input_a[8]);
  assign popcount39_lhas_core_111 = ~(input_a[21] ^ input_a[15]);
  assign popcount39_lhas_core_112 = input_a[25] | input_a[3];
  assign popcount39_lhas_core_114 = ~input_a[9];
  assign popcount39_lhas_core_116 = ~(input_a[33] & input_a[5]);
  assign popcount39_lhas_core_117 = ~input_a[22];
  assign popcount39_lhas_core_118 = ~(input_a[25] ^ input_a[31]);
  assign popcount39_lhas_core_119 = input_a[33] ^ input_a[35];
  assign popcount39_lhas_core_120 = input_a[38] ^ input_a[0];
  assign popcount39_lhas_core_121 = input_a[23] ^ input_a[18];
  assign popcount39_lhas_core_123 = input_a[22] & input_a[36];
  assign popcount39_lhas_core_124_not = ~input_a[34];
  assign popcount39_lhas_core_125 = input_a[31] ^ input_a[24];
  assign popcount39_lhas_core_126 = ~(input_a[31] & input_a[0]);
  assign popcount39_lhas_core_127 = ~(input_a[6] & input_a[35]);
  assign popcount39_lhas_core_129 = input_a[19] | input_a[6];
  assign popcount39_lhas_core_130 = input_a[17] & input_a[19];
  assign popcount39_lhas_core_131 = ~input_a[27];
  assign popcount39_lhas_core_135 = ~(input_a[35] ^ input_a[31]);
  assign popcount39_lhas_core_136 = ~(input_a[14] | input_a[5]);
  assign popcount39_lhas_core_137 = ~(input_a[23] & input_a[16]);
  assign popcount39_lhas_core_138 = ~(input_a[18] | input_a[27]);
  assign popcount39_lhas_core_139 = input_a[24] & input_a[21];
  assign popcount39_lhas_core_140 = input_a[27] ^ input_a[4];
  assign popcount39_lhas_core_141 = input_a[6] | input_a[7];
  assign popcount39_lhas_core_144_not = ~input_a[16];
  assign popcount39_lhas_core_147 = ~(input_a[24] | input_a[37]);
  assign popcount39_lhas_core_150 = ~(input_a[16] | input_a[14]);
  assign popcount39_lhas_core_151 = ~(input_a[29] & input_a[35]);
  assign popcount39_lhas_core_152 = input_a[29] | input_a[30];
  assign popcount39_lhas_core_153 = input_a[10] | input_a[8];
  assign popcount39_lhas_core_156 = ~(input_a[19] & input_a[37]);
  assign popcount39_lhas_core_157 = input_a[37] ^ input_a[10];
  assign popcount39_lhas_core_158 = ~(input_a[1] | input_a[9]);
  assign popcount39_lhas_core_160 = input_a[37] | input_a[30];
  assign popcount39_lhas_core_162 = ~(input_a[15] | input_a[29]);
  assign popcount39_lhas_core_163 = ~(input_a[10] | input_a[36]);
  assign popcount39_lhas_core_166 = input_a[22] & input_a[18];
  assign popcount39_lhas_core_167 = ~(input_a[30] ^ input_a[22]);
  assign popcount39_lhas_core_168 = ~(input_a[2] ^ input_a[11]);
  assign popcount39_lhas_core_169 = ~(input_a[30] ^ input_a[20]);
  assign popcount39_lhas_core_172 = ~input_a[16];
  assign popcount39_lhas_core_174 = ~input_a[12];
  assign popcount39_lhas_core_177 = ~input_a[22];
  assign popcount39_lhas_core_178 = input_a[8] ^ input_a[20];
  assign popcount39_lhas_core_179 = input_a[25] | input_a[34];
  assign popcount39_lhas_core_180 = ~input_a[19];
  assign popcount39_lhas_core_181 = ~(input_a[16] ^ input_a[29]);
  assign popcount39_lhas_core_182 = input_a[35] | input_a[6];
  assign popcount39_lhas_core_183 = ~(input_a[33] & input_a[8]);
  assign popcount39_lhas_core_184 = ~(input_a[11] | input_a[3]);
  assign popcount39_lhas_core_185 = input_a[30] ^ input_a[8];
  assign popcount39_lhas_core_187 = ~input_a[1];
  assign popcount39_lhas_core_188 = input_a[0] | input_a[23];
  assign popcount39_lhas_core_189_not = ~input_a[5];
  assign popcount39_lhas_core_190 = ~(input_a[33] ^ input_a[14]);
  assign popcount39_lhas_core_192 = ~(input_a[26] & input_a[22]);
  assign popcount39_lhas_core_194 = ~(input_a[27] & input_a[25]);
  assign popcount39_lhas_core_195 = input_a[36] | input_a[17];
  assign popcount39_lhas_core_196 = ~input_a[11];
  assign popcount39_lhas_core_197 = ~input_a[3];
  assign popcount39_lhas_core_198 = input_a[26] ^ input_a[0];
  assign popcount39_lhas_core_199 = ~(input_a[5] | input_a[35]);
  assign popcount39_lhas_core_200 = ~input_a[24];
  assign popcount39_lhas_core_201 = input_a[22] & input_a[2];
  assign popcount39_lhas_core_202_not = ~input_a[16];
  assign popcount39_lhas_core_203 = input_a[36] & input_a[27];
  assign popcount39_lhas_core_205 = ~(input_a[21] | input_a[7]);
  assign popcount39_lhas_core_206 = ~(input_a[5] ^ input_a[23]);
  assign popcount39_lhas_core_207 = ~input_a[19];
  assign popcount39_lhas_core_208 = ~(input_a[18] | input_a[36]);
  assign popcount39_lhas_core_210 = ~(input_a[15] & input_a[26]);
  assign popcount39_lhas_core_212 = ~(input_a[16] | input_a[23]);
  assign popcount39_lhas_core_213_not = ~input_a[4];
  assign popcount39_lhas_core_214 = ~(input_a[22] ^ input_a[0]);
  assign popcount39_lhas_core_215 = ~input_a[37];
  assign popcount39_lhas_core_216 = input_a[13] | input_a[38];
  assign popcount39_lhas_core_217 = input_a[5] & input_a[14];
  assign popcount39_lhas_core_219 = input_a[3] & input_a[18];
  assign popcount39_lhas_core_221 = ~(input_a[19] | input_a[12]);
  assign popcount39_lhas_core_224 = ~(input_a[6] ^ input_a[2]);
  assign popcount39_lhas_core_225 = input_a[28] | input_a[17];
  assign popcount39_lhas_core_226 = ~(input_a[24] ^ input_a[7]);
  assign popcount39_lhas_core_227 = ~(input_a[5] & input_a[12]);
  assign popcount39_lhas_core_228 = ~(input_a[28] | input_a[0]);
  assign popcount39_lhas_core_229 = input_a[25] ^ input_a[13];
  assign popcount39_lhas_core_231 = ~(input_a[26] ^ input_a[4]);
  assign popcount39_lhas_core_233 = input_a[34] & input_a[2];
  assign popcount39_lhas_core_234 = input_a[5] ^ input_a[36];
  assign popcount39_lhas_core_235 = ~input_a[10];
  assign popcount39_lhas_core_237 = ~(input_a[12] ^ input_a[37]);
  assign popcount39_lhas_core_238 = ~input_a[31];
  assign popcount39_lhas_core_241 = ~(input_a[33] | input_a[16]);
  assign popcount39_lhas_core_242 = ~(input_a[38] & input_a[21]);
  assign popcount39_lhas_core_243 = ~input_a[9];
  assign popcount39_lhas_core_244 = input_a[32] | input_a[20];
  assign popcount39_lhas_core_246 = input_a[17] ^ input_a[34];
  assign popcount39_lhas_core_249 = ~(input_a[15] | input_a[19]);
  assign popcount39_lhas_core_250 = input_a[32] | input_a[15];
  assign popcount39_lhas_core_251 = ~(input_a[23] ^ input_a[3]);
  assign popcount39_lhas_core_253 = ~input_a[7];
  assign popcount39_lhas_core_256 = input_a[26] ^ input_a[19];
  assign popcount39_lhas_core_258 = input_a[37] ^ input_a[22];
  assign popcount39_lhas_core_260 = ~(input_a[30] & input_a[2]);
  assign popcount39_lhas_core_262 = ~input_a[12];
  assign popcount39_lhas_core_264 = input_a[14] ^ input_a[1];
  assign popcount39_lhas_core_266 = ~(input_a[12] & input_a[14]);
  assign popcount39_lhas_core_271 = input_a[19] | input_a[28];
  assign popcount39_lhas_core_272 = input_a[20] ^ input_a[6];
  assign popcount39_lhas_core_273 = ~(input_a[30] & input_a[37]);
  assign popcount39_lhas_core_274 = input_a[19] & input_a[32];
  assign popcount39_lhas_core_276 = ~input_a[38];
  assign popcount39_lhas_core_277 = input_a[5] & input_a[38];
  assign popcount39_lhas_core_278 = ~(input_a[28] ^ input_a[15]);
  assign popcount39_lhas_core_280 = input_a[13] & input_a[22];
  assign popcount39_lhas_core_281 = ~input_a[1];
  assign popcount39_lhas_core_285 = ~(input_a[38] & input_a[38]);
  assign popcount39_lhas_core_286 = ~input_a[8];
  assign popcount39_lhas_core_287 = ~(input_a[4] ^ input_a[2]);
  assign popcount39_lhas_core_289 = input_a[38] | input_a[22];
  assign popcount39_lhas_core_292 = input_a[2] & input_a[2];
  assign popcount39_lhas_core_294 = ~(input_a[19] | input_a[1]);
  assign popcount39_lhas_core_295 = input_a[32] | input_a[18];
  assign popcount39_lhas_core_299 = ~input_a[28];
  assign popcount39_lhas_core_300 = input_a[8] | input_a[11];
  assign popcount39_lhas_core_301 = ~(input_a[8] | input_a[1]);
  assign popcount39_lhas_core_303 = ~input_a[15];
  assign popcount39_lhas_core_304 = input_a[33] ^ input_a[19];
  assign popcount39_lhas_core_306 = ~input_a[36];

  assign popcount39_lhas_out[0] = 1'b1;
  assign popcount39_lhas_out[1] = 1'b1;
  assign popcount39_lhas_out[2] = input_a[12];
  assign popcount39_lhas_out[3] = input_a[0];
  assign popcount39_lhas_out[4] = 1'b1;
  assign popcount39_lhas_out[5] = 1'b0;
endmodule