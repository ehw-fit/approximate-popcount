// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.86888
// WCE=16.0
// EP=0.88674%
// Printed PDK parameters:
//  Area=17222368.0
//  Delay=49376748.0
//  Power=644080.0

module popcount31_asyy(input [30:0] input_a, output [4:0] popcount31_asyy_out);
  wire popcount31_asyy_core_033;
  wire popcount31_asyy_core_034;
  wire popcount31_asyy_core_036;
  wire popcount31_asyy_core_037;
  wire popcount31_asyy_core_040;
  wire popcount31_asyy_core_041;
  wire popcount31_asyy_core_042;
  wire popcount31_asyy_core_044;
  wire popcount31_asyy_core_045;
  wire popcount31_asyy_core_046;
  wire popcount31_asyy_core_047;
  wire popcount31_asyy_core_050;
  wire popcount31_asyy_core_051;
  wire popcount31_asyy_core_052;
  wire popcount31_asyy_core_054;
  wire popcount31_asyy_core_055;
  wire popcount31_asyy_core_056;
  wire popcount31_asyy_core_058;
  wire popcount31_asyy_core_060_not;
  wire popcount31_asyy_core_061;
  wire popcount31_asyy_core_062;
  wire popcount31_asyy_core_063;
  wire popcount31_asyy_core_065;
  wire popcount31_asyy_core_066;
  wire popcount31_asyy_core_067_not;
  wire popcount31_asyy_core_068;
  wire popcount31_asyy_core_069;
  wire popcount31_asyy_core_072;
  wire popcount31_asyy_core_073;
  wire popcount31_asyy_core_074;
  wire popcount31_asyy_core_075;
  wire popcount31_asyy_core_076;
  wire popcount31_asyy_core_080;
  wire popcount31_asyy_core_081;
  wire popcount31_asyy_core_082_not;
  wire popcount31_asyy_core_083;
  wire popcount31_asyy_core_084;
  wire popcount31_asyy_core_085;
  wire popcount31_asyy_core_086;
  wire popcount31_asyy_core_089;
  wire popcount31_asyy_core_092;
  wire popcount31_asyy_core_095;
  wire popcount31_asyy_core_096;
  wire popcount31_asyy_core_098;
  wire popcount31_asyy_core_101;
  wire popcount31_asyy_core_102;
  wire popcount31_asyy_core_103;
  wire popcount31_asyy_core_104;
  wire popcount31_asyy_core_106;
  wire popcount31_asyy_core_109;
  wire popcount31_asyy_core_111;
  wire popcount31_asyy_core_113;
  wire popcount31_asyy_core_114;
  wire popcount31_asyy_core_116;
  wire popcount31_asyy_core_117;
  wire popcount31_asyy_core_118;
  wire popcount31_asyy_core_119;
  wire popcount31_asyy_core_120;
  wire popcount31_asyy_core_122;
  wire popcount31_asyy_core_124;
  wire popcount31_asyy_core_125;
  wire popcount31_asyy_core_126;
  wire popcount31_asyy_core_127;
  wire popcount31_asyy_core_129;
  wire popcount31_asyy_core_130;
  wire popcount31_asyy_core_131;
  wire popcount31_asyy_core_132;
  wire popcount31_asyy_core_133;
  wire popcount31_asyy_core_134;
  wire popcount31_asyy_core_135;
  wire popcount31_asyy_core_136;
  wire popcount31_asyy_core_138;
  wire popcount31_asyy_core_140;
  wire popcount31_asyy_core_147;
  wire popcount31_asyy_core_148;
  wire popcount31_asyy_core_151_not;
  wire popcount31_asyy_core_152;
  wire popcount31_asyy_core_153;
  wire popcount31_asyy_core_156_not;
  wire popcount31_asyy_core_158;
  wire popcount31_asyy_core_159;
  wire popcount31_asyy_core_161;
  wire popcount31_asyy_core_162;
  wire popcount31_asyy_core_163;
  wire popcount31_asyy_core_164;
  wire popcount31_asyy_core_165;
  wire popcount31_asyy_core_166;
  wire popcount31_asyy_core_167;
  wire popcount31_asyy_core_169;
  wire popcount31_asyy_core_170;
  wire popcount31_asyy_core_171;
  wire popcount31_asyy_core_172;
  wire popcount31_asyy_core_173;
  wire popcount31_asyy_core_174;
  wire popcount31_asyy_core_175;
  wire popcount31_asyy_core_176;
  wire popcount31_asyy_core_177;
  wire popcount31_asyy_core_178;
  wire popcount31_asyy_core_179;
  wire popcount31_asyy_core_180;
  wire popcount31_asyy_core_181;
  wire popcount31_asyy_core_182;
  wire popcount31_asyy_core_183;
  wire popcount31_asyy_core_184;
  wire popcount31_asyy_core_186;
  wire popcount31_asyy_core_190;
  wire popcount31_asyy_core_191;
  wire popcount31_asyy_core_194;
  wire popcount31_asyy_core_195;
  wire popcount31_asyy_core_196;
  wire popcount31_asyy_core_198;
  wire popcount31_asyy_core_202;
  wire popcount31_asyy_core_208;
  wire popcount31_asyy_core_209;
  wire popcount31_asyy_core_210;
  wire popcount31_asyy_core_211;
  wire popcount31_asyy_core_212;
  wire popcount31_asyy_core_213;
  wire popcount31_asyy_core_214;
  wire popcount31_asyy_core_215;
  wire popcount31_asyy_core_218;

  assign popcount31_asyy_core_033 = ~(input_a[9] & input_a[14]);
  assign popcount31_asyy_core_034 = ~(input_a[29] & input_a[15]);
  assign popcount31_asyy_core_036 = ~(input_a[13] | input_a[3]);
  assign popcount31_asyy_core_037 = input_a[29] & input_a[12];
  assign popcount31_asyy_core_040 = input_a[28] & input_a[8];
  assign popcount31_asyy_core_041 = input_a[11] ^ input_a[4];
  assign popcount31_asyy_core_042 = input_a[21] & input_a[16];
  assign popcount31_asyy_core_044 = ~(input_a[27] & input_a[5]);
  assign popcount31_asyy_core_045 = ~(input_a[15] ^ input_a[5]);
  assign popcount31_asyy_core_046 = popcount31_asyy_core_040 & popcount31_asyy_core_042;
  assign popcount31_asyy_core_047 = ~(input_a[19] | input_a[5]);
  assign popcount31_asyy_core_050 = input_a[24] ^ input_a[16];
  assign popcount31_asyy_core_051 = input_a[6] ^ input_a[19];
  assign popcount31_asyy_core_052 = input_a[15] ^ input_a[16];
  assign popcount31_asyy_core_054 = ~(input_a[3] | input_a[28]);
  assign popcount31_asyy_core_055 = input_a[15] ^ input_a[10];
  assign popcount31_asyy_core_056 = ~input_a[28];
  assign popcount31_asyy_core_058 = ~(input_a[30] ^ input_a[4]);
  assign popcount31_asyy_core_060_not = ~input_a[11];
  assign popcount31_asyy_core_061 = ~input_a[16];
  assign popcount31_asyy_core_062 = input_a[19] ^ input_a[1];
  assign popcount31_asyy_core_063 = ~input_a[8];
  assign popcount31_asyy_core_065 = ~(input_a[19] ^ input_a[25]);
  assign popcount31_asyy_core_066 = ~input_a[25];
  assign popcount31_asyy_core_067_not = ~input_a[24];
  assign popcount31_asyy_core_068 = input_a[25] ^ input_a[15];
  assign popcount31_asyy_core_069 = input_a[26] ^ input_a[13];
  assign popcount31_asyy_core_072 = input_a[0] & input_a[27];
  assign popcount31_asyy_core_073 = ~input_a[8];
  assign popcount31_asyy_core_074 = ~input_a[21];
  assign popcount31_asyy_core_075 = ~(input_a[22] & input_a[8]);
  assign popcount31_asyy_core_076 = input_a[0] | input_a[29];
  assign popcount31_asyy_core_080 = input_a[1] ^ input_a[30];
  assign popcount31_asyy_core_081 = input_a[13] | input_a[22];
  assign popcount31_asyy_core_082_not = ~input_a[13];
  assign popcount31_asyy_core_083 = ~(input_a[20] & input_a[2]);
  assign popcount31_asyy_core_084 = input_a[7] & input_a[8];
  assign popcount31_asyy_core_085 = input_a[0] & input_a[23];
  assign popcount31_asyy_core_086 = ~(input_a[28] ^ input_a[3]);
  assign popcount31_asyy_core_089 = ~input_a[2];
  assign popcount31_asyy_core_092 = input_a[14] ^ input_a[18];
  assign popcount31_asyy_core_095 = ~(input_a[28] | input_a[18]);
  assign popcount31_asyy_core_096 = input_a[4] | input_a[6];
  assign popcount31_asyy_core_098 = ~(input_a[9] | input_a[28]);
  assign popcount31_asyy_core_101 = ~(input_a[28] | input_a[5]);
  assign popcount31_asyy_core_102 = ~(input_a[2] | input_a[8]);
  assign popcount31_asyy_core_103 = input_a[8] & input_a[16];
  assign popcount31_asyy_core_104 = popcount31_asyy_core_046 & input_a[12];
  assign popcount31_asyy_core_106 = input_a[8] & input_a[6];
  assign popcount31_asyy_core_109 = input_a[19] ^ input_a[20];
  assign popcount31_asyy_core_111 = ~(input_a[12] | input_a[0]);
  assign popcount31_asyy_core_113 = ~input_a[7];
  assign popcount31_asyy_core_114 = input_a[28] ^ input_a[17];
  assign popcount31_asyy_core_116 = input_a[6] ^ input_a[11];
  assign popcount31_asyy_core_117 = ~(input_a[26] ^ input_a[9]);
  assign popcount31_asyy_core_118 = ~(input_a[11] ^ input_a[25]);
  assign popcount31_asyy_core_119 = ~(input_a[2] & input_a[21]);
  assign popcount31_asyy_core_120 = ~input_a[11];
  assign popcount31_asyy_core_122 = ~(input_a[18] & input_a[22]);
  assign popcount31_asyy_core_124 = input_a[29] | input_a[9];
  assign popcount31_asyy_core_125 = input_a[3] & input_a[8];
  assign popcount31_asyy_core_126 = input_a[20] ^ input_a[1];
  assign popcount31_asyy_core_127 = input_a[10] ^ input_a[16];
  assign popcount31_asyy_core_129 = ~input_a[7];
  assign popcount31_asyy_core_130 = input_a[27] | input_a[10];
  assign popcount31_asyy_core_131 = ~(input_a[22] | input_a[9]);
  assign popcount31_asyy_core_132 = ~input_a[8];
  assign popcount31_asyy_core_133 = input_a[27] ^ input_a[25];
  assign popcount31_asyy_core_134 = ~(input_a[11] ^ input_a[27]);
  assign popcount31_asyy_core_135 = ~(input_a[10] ^ input_a[1]);
  assign popcount31_asyy_core_136 = input_a[26] ^ input_a[29];
  assign popcount31_asyy_core_138 = ~(input_a[24] | input_a[15]);
  assign popcount31_asyy_core_140 = input_a[21] & input_a[10];
  assign popcount31_asyy_core_147 = ~(input_a[9] | input_a[15]);
  assign popcount31_asyy_core_148 = input_a[20] & input_a[23];
  assign popcount31_asyy_core_151_not = ~input_a[6];
  assign popcount31_asyy_core_152 = ~(input_a[6] | input_a[15]);
  assign popcount31_asyy_core_153 = ~popcount31_asyy_core_148;
  assign popcount31_asyy_core_156_not = ~input_a[5];
  assign popcount31_asyy_core_158 = input_a[12] & input_a[6];
  assign popcount31_asyy_core_159 = input_a[26] & input_a[3];
  assign popcount31_asyy_core_161 = input_a[11] & input_a[0];
  assign popcount31_asyy_core_162 = input_a[30] | input_a[4];
  assign popcount31_asyy_core_163 = input_a[18] & input_a[27];
  assign popcount31_asyy_core_164 = popcount31_asyy_core_159 ^ popcount31_asyy_core_161;
  assign popcount31_asyy_core_165 = popcount31_asyy_core_159 & popcount31_asyy_core_161;
  assign popcount31_asyy_core_166 = popcount31_asyy_core_164 | popcount31_asyy_core_163;
  assign popcount31_asyy_core_167 = ~(input_a[22] | input_a[17]);
  assign popcount31_asyy_core_169 = ~(input_a[9] | input_a[27]);
  assign popcount31_asyy_core_170 = input_a[14] & input_a[29];
  assign popcount31_asyy_core_171 = popcount31_asyy_core_153 ^ popcount31_asyy_core_166;
  assign popcount31_asyy_core_172 = popcount31_asyy_core_153 & popcount31_asyy_core_166;
  assign popcount31_asyy_core_173 = popcount31_asyy_core_171 ^ popcount31_asyy_core_170;
  assign popcount31_asyy_core_174 = popcount31_asyy_core_171 & popcount31_asyy_core_170;
  assign popcount31_asyy_core_175 = popcount31_asyy_core_172 | popcount31_asyy_core_174;
  assign popcount31_asyy_core_176 = popcount31_asyy_core_148 ^ popcount31_asyy_core_165;
  assign popcount31_asyy_core_177 = popcount31_asyy_core_148 & popcount31_asyy_core_165;
  assign popcount31_asyy_core_178 = popcount31_asyy_core_176 ^ popcount31_asyy_core_175;
  assign popcount31_asyy_core_179 = popcount31_asyy_core_176 & popcount31_asyy_core_175;
  assign popcount31_asyy_core_180 = popcount31_asyy_core_177 | popcount31_asyy_core_179;
  assign popcount31_asyy_core_181 = ~(input_a[18] ^ input_a[27]);
  assign popcount31_asyy_core_182 = ~input_a[22];
  assign popcount31_asyy_core_183 = input_a[24] ^ input_a[23];
  assign popcount31_asyy_core_184 = input_a[10] & popcount31_asyy_core_173;
  assign popcount31_asyy_core_186 = ~(input_a[15] & input_a[12]);
  assign popcount31_asyy_core_190 = popcount31_asyy_core_178 ^ popcount31_asyy_core_184;
  assign popcount31_asyy_core_191 = popcount31_asyy_core_178 & popcount31_asyy_core_184;
  assign popcount31_asyy_core_194 = input_a[5] & input_a[15];
  assign popcount31_asyy_core_195 = popcount31_asyy_core_180 | popcount31_asyy_core_191;
  assign popcount31_asyy_core_196 = ~(input_a[6] ^ input_a[2]);
  assign popcount31_asyy_core_198 = ~(input_a[12] & input_a[17]);
  assign popcount31_asyy_core_202 = ~(input_a[4] & input_a[17]);
  assign popcount31_asyy_core_208 = input_a[17] & input_a[4];
  assign popcount31_asyy_core_209 = popcount31_asyy_core_190 | popcount31_asyy_core_208;
  assign popcount31_asyy_core_210 = popcount31_asyy_core_104 ^ popcount31_asyy_core_195;
  assign popcount31_asyy_core_211 = popcount31_asyy_core_104 & popcount31_asyy_core_195;
  assign popcount31_asyy_core_212 = popcount31_asyy_core_210 ^ popcount31_asyy_core_209;
  assign popcount31_asyy_core_213 = popcount31_asyy_core_210 & popcount31_asyy_core_209;
  assign popcount31_asyy_core_214 = popcount31_asyy_core_211 | popcount31_asyy_core_213;
  assign popcount31_asyy_core_215 = ~(input_a[9] ^ input_a[1]);
  assign popcount31_asyy_core_218 = ~(input_a[14] & input_a[6]);

  assign popcount31_asyy_out[0] = input_a[5];
  assign popcount31_asyy_out[1] = popcount31_asyy_core_202;
  assign popcount31_asyy_out[2] = 1'b1;
  assign popcount31_asyy_out[3] = popcount31_asyy_core_212;
  assign popcount31_asyy_out[4] = popcount31_asyy_core_214;
endmodule