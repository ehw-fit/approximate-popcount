// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.97801
// WCE=24.0
// EP=0.936686%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_8xzl(input [29:0] input_a, output [4:0] popcount30_8xzl_out);
  wire popcount30_8xzl_core_032;
  wire popcount30_8xzl_core_033;
  wire popcount30_8xzl_core_034;
  wire popcount30_8xzl_core_035;
  wire popcount30_8xzl_core_036;
  wire popcount30_8xzl_core_037;
  wire popcount30_8xzl_core_038;
  wire popcount30_8xzl_core_040;
  wire popcount30_8xzl_core_041;
  wire popcount30_8xzl_core_043_not;
  wire popcount30_8xzl_core_044;
  wire popcount30_8xzl_core_045;
  wire popcount30_8xzl_core_046;
  wire popcount30_8xzl_core_048;
  wire popcount30_8xzl_core_049;
  wire popcount30_8xzl_core_055;
  wire popcount30_8xzl_core_056;
  wire popcount30_8xzl_core_057;
  wire popcount30_8xzl_core_058;
  wire popcount30_8xzl_core_059;
  wire popcount30_8xzl_core_060;
  wire popcount30_8xzl_core_061;
  wire popcount30_8xzl_core_062;
  wire popcount30_8xzl_core_064;
  wire popcount30_8xzl_core_065;
  wire popcount30_8xzl_core_066;
  wire popcount30_8xzl_core_067;
  wire popcount30_8xzl_core_069;
  wire popcount30_8xzl_core_070;
  wire popcount30_8xzl_core_072;
  wire popcount30_8xzl_core_073;
  wire popcount30_8xzl_core_074;
  wire popcount30_8xzl_core_075;
  wire popcount30_8xzl_core_076;
  wire popcount30_8xzl_core_078;
  wire popcount30_8xzl_core_079;
  wire popcount30_8xzl_core_080;
  wire popcount30_8xzl_core_082;
  wire popcount30_8xzl_core_084;
  wire popcount30_8xzl_core_086;
  wire popcount30_8xzl_core_088;
  wire popcount30_8xzl_core_090;
  wire popcount30_8xzl_core_091;
  wire popcount30_8xzl_core_092;
  wire popcount30_8xzl_core_093;
  wire popcount30_8xzl_core_095;
  wire popcount30_8xzl_core_096;
  wire popcount30_8xzl_core_097;
  wire popcount30_8xzl_core_099;
  wire popcount30_8xzl_core_100;
  wire popcount30_8xzl_core_102;
  wire popcount30_8xzl_core_103;
  wire popcount30_8xzl_core_104;
  wire popcount30_8xzl_core_106;
  wire popcount30_8xzl_core_107;
  wire popcount30_8xzl_core_108;
  wire popcount30_8xzl_core_111;
  wire popcount30_8xzl_core_112;
  wire popcount30_8xzl_core_115;
  wire popcount30_8xzl_core_116_not;
  wire popcount30_8xzl_core_118;
  wire popcount30_8xzl_core_119;
  wire popcount30_8xzl_core_120;
  wire popcount30_8xzl_core_121;
  wire popcount30_8xzl_core_122;
  wire popcount30_8xzl_core_126;
  wire popcount30_8xzl_core_127;
  wire popcount30_8xzl_core_128;
  wire popcount30_8xzl_core_129;
  wire popcount30_8xzl_core_130;
  wire popcount30_8xzl_core_131;
  wire popcount30_8xzl_core_132;
  wire popcount30_8xzl_core_133;
  wire popcount30_8xzl_core_137;
  wire popcount30_8xzl_core_138;
  wire popcount30_8xzl_core_140;
  wire popcount30_8xzl_core_142;
  wire popcount30_8xzl_core_144;
  wire popcount30_8xzl_core_145_not;
  wire popcount30_8xzl_core_146;
  wire popcount30_8xzl_core_147;
  wire popcount30_8xzl_core_148;
  wire popcount30_8xzl_core_152;
  wire popcount30_8xzl_core_153;
  wire popcount30_8xzl_core_154;
  wire popcount30_8xzl_core_156;
  wire popcount30_8xzl_core_158;
  wire popcount30_8xzl_core_162;
  wire popcount30_8xzl_core_164_not;
  wire popcount30_8xzl_core_165;
  wire popcount30_8xzl_core_166;
  wire popcount30_8xzl_core_167;
  wire popcount30_8xzl_core_174;
  wire popcount30_8xzl_core_175;
  wire popcount30_8xzl_core_177;
  wire popcount30_8xzl_core_179;
  wire popcount30_8xzl_core_181;
  wire popcount30_8xzl_core_183;
  wire popcount30_8xzl_core_184;
  wire popcount30_8xzl_core_185;
  wire popcount30_8xzl_core_186;
  wire popcount30_8xzl_core_187;
  wire popcount30_8xzl_core_188;
  wire popcount30_8xzl_core_193;
  wire popcount30_8xzl_core_194;
  wire popcount30_8xzl_core_195;
  wire popcount30_8xzl_core_196;
  wire popcount30_8xzl_core_197;
  wire popcount30_8xzl_core_199;
  wire popcount30_8xzl_core_200;
  wire popcount30_8xzl_core_203;
  wire popcount30_8xzl_core_204;
  wire popcount30_8xzl_core_207;
  wire popcount30_8xzl_core_211;
  wire popcount30_8xzl_core_212;

  assign popcount30_8xzl_core_032 = input_a[19] ^ input_a[6];
  assign popcount30_8xzl_core_033 = ~(input_a[16] ^ input_a[25]);
  assign popcount30_8xzl_core_034 = ~(input_a[11] & input_a[19]);
  assign popcount30_8xzl_core_035 = input_a[11] ^ input_a[3];
  assign popcount30_8xzl_core_036 = input_a[10] ^ input_a[25];
  assign popcount30_8xzl_core_037 = input_a[24] | input_a[2];
  assign popcount30_8xzl_core_038 = input_a[2] & input_a[6];
  assign popcount30_8xzl_core_040 = input_a[7] | input_a[21];
  assign popcount30_8xzl_core_041 = input_a[27] & input_a[18];
  assign popcount30_8xzl_core_043_not = ~input_a[17];
  assign popcount30_8xzl_core_044 = ~(input_a[0] ^ input_a[11]);
  assign popcount30_8xzl_core_045 = ~(input_a[12] & input_a[21]);
  assign popcount30_8xzl_core_046 = input_a[11] & input_a[20];
  assign popcount30_8xzl_core_048 = input_a[18] ^ input_a[16];
  assign popcount30_8xzl_core_049 = input_a[29] | input_a[19];
  assign popcount30_8xzl_core_055 = ~(input_a[27] ^ input_a[2]);
  assign popcount30_8xzl_core_056 = ~input_a[1];
  assign popcount30_8xzl_core_057 = ~input_a[24];
  assign popcount30_8xzl_core_058 = input_a[7] & input_a[12];
  assign popcount30_8xzl_core_059 = ~(input_a[22] | input_a[4]);
  assign popcount30_8xzl_core_060 = ~(input_a[0] | input_a[1]);
  assign popcount30_8xzl_core_061 = ~input_a[0];
  assign popcount30_8xzl_core_062 = input_a[7] & input_a[8];
  assign popcount30_8xzl_core_064 = input_a[19] & input_a[11];
  assign popcount30_8xzl_core_065 = ~input_a[10];
  assign popcount30_8xzl_core_066 = ~input_a[10];
  assign popcount30_8xzl_core_067 = input_a[20] & input_a[22];
  assign popcount30_8xzl_core_069 = ~(input_a[21] ^ input_a[11]);
  assign popcount30_8xzl_core_070 = input_a[15] ^ input_a[25];
  assign popcount30_8xzl_core_072 = ~(input_a[9] & input_a[25]);
  assign popcount30_8xzl_core_073 = ~(input_a[18] ^ input_a[12]);
  assign popcount30_8xzl_core_074 = ~(input_a[24] | input_a[14]);
  assign popcount30_8xzl_core_075 = ~(input_a[26] & input_a[7]);
  assign popcount30_8xzl_core_076 = ~(input_a[15] ^ input_a[6]);
  assign popcount30_8xzl_core_078 = ~(input_a[19] | input_a[26]);
  assign popcount30_8xzl_core_079 = ~input_a[5];
  assign popcount30_8xzl_core_080 = ~(input_a[26] ^ input_a[24]);
  assign popcount30_8xzl_core_082 = ~input_a[24];
  assign popcount30_8xzl_core_084 = ~(input_a[7] ^ input_a[10]);
  assign popcount30_8xzl_core_086 = input_a[18] | input_a[3];
  assign popcount30_8xzl_core_088 = ~input_a[24];
  assign popcount30_8xzl_core_090 = ~input_a[9];
  assign popcount30_8xzl_core_091 = input_a[13] & input_a[6];
  assign popcount30_8xzl_core_092 = ~(input_a[18] ^ input_a[20]);
  assign popcount30_8xzl_core_093 = input_a[12] & input_a[26];
  assign popcount30_8xzl_core_095 = ~(input_a[7] | input_a[20]);
  assign popcount30_8xzl_core_096 = input_a[0] & input_a[15];
  assign popcount30_8xzl_core_097 = input_a[12] | input_a[20];
  assign popcount30_8xzl_core_099 = input_a[24] & input_a[11];
  assign popcount30_8xzl_core_100 = ~(input_a[7] ^ input_a[9]);
  assign popcount30_8xzl_core_102 = ~(input_a[1] | input_a[11]);
  assign popcount30_8xzl_core_103 = ~(input_a[1] & input_a[2]);
  assign popcount30_8xzl_core_104 = ~(input_a[16] | input_a[24]);
  assign popcount30_8xzl_core_106 = ~(input_a[0] & input_a[17]);
  assign popcount30_8xzl_core_107 = ~(input_a[11] & input_a[18]);
  assign popcount30_8xzl_core_108 = ~(input_a[25] & input_a[4]);
  assign popcount30_8xzl_core_111 = input_a[17] ^ input_a[17];
  assign popcount30_8xzl_core_112 = input_a[11] ^ input_a[13];
  assign popcount30_8xzl_core_115 = input_a[7] | input_a[9];
  assign popcount30_8xzl_core_116_not = ~input_a[17];
  assign popcount30_8xzl_core_118 = ~input_a[10];
  assign popcount30_8xzl_core_119 = ~(input_a[2] | input_a[0]);
  assign popcount30_8xzl_core_120 = ~(input_a[5] & input_a[5]);
  assign popcount30_8xzl_core_121 = ~(input_a[20] & input_a[2]);
  assign popcount30_8xzl_core_122 = input_a[14] ^ input_a[2];
  assign popcount30_8xzl_core_126 = ~(input_a[25] | input_a[11]);
  assign popcount30_8xzl_core_127 = input_a[14] & input_a[11];
  assign popcount30_8xzl_core_128 = ~input_a[11];
  assign popcount30_8xzl_core_129 = input_a[2] | input_a[28];
  assign popcount30_8xzl_core_130 = input_a[5] ^ input_a[19];
  assign popcount30_8xzl_core_131 = ~(input_a[12] | input_a[0]);
  assign popcount30_8xzl_core_132 = ~(input_a[7] & input_a[16]);
  assign popcount30_8xzl_core_133 = ~(input_a[26] | input_a[19]);
  assign popcount30_8xzl_core_137 = ~(input_a[3] | input_a[13]);
  assign popcount30_8xzl_core_138 = input_a[27] & input_a[27];
  assign popcount30_8xzl_core_140 = ~(input_a[2] & input_a[27]);
  assign popcount30_8xzl_core_142 = input_a[5] ^ input_a[28];
  assign popcount30_8xzl_core_144 = input_a[8] & input_a[23];
  assign popcount30_8xzl_core_145_not = ~input_a[25];
  assign popcount30_8xzl_core_146 = ~(input_a[0] & input_a[5]);
  assign popcount30_8xzl_core_147 = input_a[23] & input_a[8];
  assign popcount30_8xzl_core_148 = ~(input_a[27] | input_a[7]);
  assign popcount30_8xzl_core_152 = ~(input_a[24] & input_a[28]);
  assign popcount30_8xzl_core_153 = input_a[9] ^ input_a[19];
  assign popcount30_8xzl_core_154 = ~(input_a[17] | input_a[1]);
  assign popcount30_8xzl_core_156 = ~(input_a[23] | input_a[25]);
  assign popcount30_8xzl_core_158 = ~(input_a[6] | input_a[27]);
  assign popcount30_8xzl_core_162 = input_a[11] & input_a[6];
  assign popcount30_8xzl_core_164_not = ~input_a[22];
  assign popcount30_8xzl_core_165 = input_a[12] ^ input_a[11];
  assign popcount30_8xzl_core_166 = ~(input_a[9] ^ input_a[10]);
  assign popcount30_8xzl_core_167 = ~input_a[13];
  assign popcount30_8xzl_core_174 = ~(input_a[27] ^ input_a[7]);
  assign popcount30_8xzl_core_175 = input_a[21] ^ input_a[7];
  assign popcount30_8xzl_core_177 = input_a[20] ^ input_a[1];
  assign popcount30_8xzl_core_179 = ~(input_a[18] ^ input_a[3]);
  assign popcount30_8xzl_core_181 = input_a[17] | input_a[11];
  assign popcount30_8xzl_core_183 = ~(input_a[26] & input_a[2]);
  assign popcount30_8xzl_core_184 = ~input_a[17];
  assign popcount30_8xzl_core_185 = ~(input_a[17] & input_a[26]);
  assign popcount30_8xzl_core_186 = ~(input_a[22] | input_a[0]);
  assign popcount30_8xzl_core_187 = ~(input_a[21] | input_a[15]);
  assign popcount30_8xzl_core_188 = input_a[7] ^ input_a[25];
  assign popcount30_8xzl_core_193 = input_a[11] ^ input_a[11];
  assign popcount30_8xzl_core_194 = input_a[18] | input_a[2];
  assign popcount30_8xzl_core_195 = ~input_a[15];
  assign popcount30_8xzl_core_196 = input_a[4] & input_a[14];
  assign popcount30_8xzl_core_197 = input_a[4] & input_a[15];
  assign popcount30_8xzl_core_199 = ~(input_a[8] ^ input_a[25]);
  assign popcount30_8xzl_core_200 = input_a[14] ^ input_a[15];
  assign popcount30_8xzl_core_203 = input_a[23] ^ input_a[1];
  assign popcount30_8xzl_core_204 = input_a[15] ^ input_a[19];
  assign popcount30_8xzl_core_207 = ~input_a[29];
  assign popcount30_8xzl_core_211 = ~(input_a[6] | input_a[0]);
  assign popcount30_8xzl_core_212 = input_a[9] | input_a[23];

  assign popcount30_8xzl_out[0] = input_a[10];
  assign popcount30_8xzl_out[1] = input_a[25];
  assign popcount30_8xzl_out[2] = 1'b1;
  assign popcount30_8xzl_out[3] = 1'b1;
  assign popcount30_8xzl_out[4] = 1'b0;
endmodule