// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.01826
// WCE=12.0
// EP=0.845828%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_vqp7(input [21:0] input_a, output [4:0] popcount22_vqp7_out);
  wire popcount22_vqp7_core_024;
  wire popcount22_vqp7_core_025;
  wire popcount22_vqp7_core_026;
  wire popcount22_vqp7_core_028;
  wire popcount22_vqp7_core_030;
  wire popcount22_vqp7_core_031;
  wire popcount22_vqp7_core_032;
  wire popcount22_vqp7_core_033;
  wire popcount22_vqp7_core_034;
  wire popcount22_vqp7_core_036;
  wire popcount22_vqp7_core_037;
  wire popcount22_vqp7_core_038;
  wire popcount22_vqp7_core_039;
  wire popcount22_vqp7_core_040;
  wire popcount22_vqp7_core_041;
  wire popcount22_vqp7_core_042;
  wire popcount22_vqp7_core_044;
  wire popcount22_vqp7_core_046;
  wire popcount22_vqp7_core_047;
  wire popcount22_vqp7_core_049;
  wire popcount22_vqp7_core_052;
  wire popcount22_vqp7_core_053;
  wire popcount22_vqp7_core_054;
  wire popcount22_vqp7_core_058;
  wire popcount22_vqp7_core_059;
  wire popcount22_vqp7_core_060;
  wire popcount22_vqp7_core_061;
  wire popcount22_vqp7_core_062;
  wire popcount22_vqp7_core_063;
  wire popcount22_vqp7_core_064;
  wire popcount22_vqp7_core_067;
  wire popcount22_vqp7_core_070;
  wire popcount22_vqp7_core_075;
  wire popcount22_vqp7_core_076;
  wire popcount22_vqp7_core_078;
  wire popcount22_vqp7_core_079;
  wire popcount22_vqp7_core_080;
  wire popcount22_vqp7_core_081;
  wire popcount22_vqp7_core_082;
  wire popcount22_vqp7_core_083;
  wire popcount22_vqp7_core_084;
  wire popcount22_vqp7_core_085;
  wire popcount22_vqp7_core_086;
  wire popcount22_vqp7_core_087;
  wire popcount22_vqp7_core_088;
  wire popcount22_vqp7_core_089;
  wire popcount22_vqp7_core_090;
  wire popcount22_vqp7_core_091_not;
  wire popcount22_vqp7_core_092;
  wire popcount22_vqp7_core_095;
  wire popcount22_vqp7_core_098;
  wire popcount22_vqp7_core_100;
  wire popcount22_vqp7_core_103;
  wire popcount22_vqp7_core_104;
  wire popcount22_vqp7_core_108;
  wire popcount22_vqp7_core_109;
  wire popcount22_vqp7_core_112;
  wire popcount22_vqp7_core_119;
  wire popcount22_vqp7_core_120;
  wire popcount22_vqp7_core_121;
  wire popcount22_vqp7_core_123;
  wire popcount22_vqp7_core_124;
  wire popcount22_vqp7_core_125;
  wire popcount22_vqp7_core_127;
  wire popcount22_vqp7_core_128;
  wire popcount22_vqp7_core_130;
  wire popcount22_vqp7_core_133;
  wire popcount22_vqp7_core_135;
  wire popcount22_vqp7_core_136;
  wire popcount22_vqp7_core_137;
  wire popcount22_vqp7_core_139;
  wire popcount22_vqp7_core_140;
  wire popcount22_vqp7_core_141;
  wire popcount22_vqp7_core_142;
  wire popcount22_vqp7_core_144;
  wire popcount22_vqp7_core_146;
  wire popcount22_vqp7_core_147;
  wire popcount22_vqp7_core_149;
  wire popcount22_vqp7_core_152;
  wire popcount22_vqp7_core_155;
  wire popcount22_vqp7_core_157;
  wire popcount22_vqp7_core_160;
  wire popcount22_vqp7_core_161;

  assign popcount22_vqp7_core_024 = ~(input_a[8] | input_a[12]);
  assign popcount22_vqp7_core_025 = input_a[12] & input_a[13];
  assign popcount22_vqp7_core_026 = input_a[13] & input_a[15];
  assign popcount22_vqp7_core_028 = input_a[5] ^ input_a[1];
  assign popcount22_vqp7_core_030 = input_a[16] | input_a[0];
  assign popcount22_vqp7_core_031 = ~(input_a[12] & input_a[21]);
  assign popcount22_vqp7_core_032 = ~(input_a[1] | input_a[9]);
  assign popcount22_vqp7_core_033 = input_a[3] | input_a[2];
  assign popcount22_vqp7_core_034 = input_a[1] | input_a[16];
  assign popcount22_vqp7_core_036 = input_a[4] | input_a[12];
  assign popcount22_vqp7_core_037 = ~(input_a[12] | input_a[20]);
  assign popcount22_vqp7_core_038 = ~(input_a[5] | input_a[12]);
  assign popcount22_vqp7_core_039 = ~(input_a[2] | input_a[3]);
  assign popcount22_vqp7_core_040 = ~(input_a[16] & input_a[0]);
  assign popcount22_vqp7_core_041 = ~(input_a[8] & input_a[16]);
  assign popcount22_vqp7_core_042 = ~(input_a[13] ^ input_a[14]);
  assign popcount22_vqp7_core_044 = input_a[6] & input_a[4];
  assign popcount22_vqp7_core_046 = ~(input_a[0] | input_a[12]);
  assign popcount22_vqp7_core_047 = ~(input_a[15] | input_a[9]);
  assign popcount22_vqp7_core_049 = input_a[9] ^ input_a[9];
  assign popcount22_vqp7_core_052 = input_a[4] & input_a[2];
  assign popcount22_vqp7_core_053 = ~(input_a[16] & input_a[2]);
  assign popcount22_vqp7_core_054 = input_a[7] | input_a[3];
  assign popcount22_vqp7_core_058 = ~(input_a[6] & input_a[18]);
  assign popcount22_vqp7_core_059 = ~(input_a[14] & input_a[20]);
  assign popcount22_vqp7_core_060 = input_a[10] | input_a[18];
  assign popcount22_vqp7_core_061 = input_a[0] & input_a[9];
  assign popcount22_vqp7_core_062 = ~(input_a[10] | input_a[10]);
  assign popcount22_vqp7_core_063 = input_a[20] ^ input_a[1];
  assign popcount22_vqp7_core_064 = input_a[18] | input_a[15];
  assign popcount22_vqp7_core_067 = input_a[10] ^ input_a[0];
  assign popcount22_vqp7_core_070 = input_a[19] & input_a[18];
  assign popcount22_vqp7_core_075 = ~input_a[6];
  assign popcount22_vqp7_core_076 = input_a[15] & input_a[6];
  assign popcount22_vqp7_core_078 = input_a[1] & input_a[7];
  assign popcount22_vqp7_core_079 = input_a[1] | input_a[1];
  assign popcount22_vqp7_core_080 = input_a[14] ^ input_a[21];
  assign popcount22_vqp7_core_081 = ~(input_a[4] & input_a[10]);
  assign popcount22_vqp7_core_082 = input_a[6] | input_a[20];
  assign popcount22_vqp7_core_083 = ~input_a[21];
  assign popcount22_vqp7_core_084 = input_a[15] & input_a[0];
  assign popcount22_vqp7_core_085 = ~(input_a[19] | input_a[0]);
  assign popcount22_vqp7_core_086 = input_a[15] & input_a[2];
  assign popcount22_vqp7_core_087 = input_a[11] ^ input_a[19];
  assign popcount22_vqp7_core_088 = ~(input_a[21] | input_a[21]);
  assign popcount22_vqp7_core_089 = ~(input_a[12] ^ input_a[0]);
  assign popcount22_vqp7_core_090 = input_a[15] | input_a[15];
  assign popcount22_vqp7_core_091_not = ~input_a[6];
  assign popcount22_vqp7_core_092 = input_a[6] | input_a[6];
  assign popcount22_vqp7_core_095 = ~(input_a[19] ^ input_a[20]);
  assign popcount22_vqp7_core_098 = ~(input_a[14] & input_a[7]);
  assign popcount22_vqp7_core_100 = input_a[20] ^ input_a[0];
  assign popcount22_vqp7_core_103 = ~(input_a[19] ^ input_a[4]);
  assign popcount22_vqp7_core_104 = input_a[3] ^ input_a[5];
  assign popcount22_vqp7_core_108 = ~(input_a[18] ^ input_a[9]);
  assign popcount22_vqp7_core_109 = ~input_a[4];
  assign popcount22_vqp7_core_112 = ~(input_a[16] ^ input_a[11]);
  assign popcount22_vqp7_core_119 = input_a[17] | input_a[14];
  assign popcount22_vqp7_core_120 = input_a[6] ^ input_a[5];
  assign popcount22_vqp7_core_121 = ~(input_a[16] | input_a[1]);
  assign popcount22_vqp7_core_123 = input_a[12] ^ input_a[6];
  assign popcount22_vqp7_core_124 = input_a[21] ^ input_a[12];
  assign popcount22_vqp7_core_125 = ~(input_a[5] ^ input_a[2]);
  assign popcount22_vqp7_core_127 = input_a[2] ^ input_a[5];
  assign popcount22_vqp7_core_128 = ~(input_a[2] | input_a[21]);
  assign popcount22_vqp7_core_130 = input_a[14] & input_a[10];
  assign popcount22_vqp7_core_133 = ~(input_a[14] & input_a[0]);
  assign popcount22_vqp7_core_135 = ~(input_a[2] ^ input_a[9]);
  assign popcount22_vqp7_core_136 = ~(input_a[20] ^ input_a[20]);
  assign popcount22_vqp7_core_137 = ~(input_a[16] & input_a[16]);
  assign popcount22_vqp7_core_139 = ~(input_a[4] & input_a[9]);
  assign popcount22_vqp7_core_140 = ~(input_a[19] ^ input_a[19]);
  assign popcount22_vqp7_core_141 = ~(input_a[10] ^ input_a[12]);
  assign popcount22_vqp7_core_142 = ~(input_a[19] & input_a[2]);
  assign popcount22_vqp7_core_144 = input_a[17] & input_a[0];
  assign popcount22_vqp7_core_146 = ~(input_a[15] ^ input_a[7]);
  assign popcount22_vqp7_core_147 = ~(input_a[17] | input_a[20]);
  assign popcount22_vqp7_core_149 = ~(input_a[5] | input_a[19]);
  assign popcount22_vqp7_core_152 = input_a[19] ^ input_a[21];
  assign popcount22_vqp7_core_155 = ~input_a[6];
  assign popcount22_vqp7_core_157 = input_a[15] | input_a[21];
  assign popcount22_vqp7_core_160 = input_a[21] & input_a[21];
  assign popcount22_vqp7_core_161 = ~(input_a[17] & input_a[7]);

  assign popcount22_vqp7_out[0] = 1'b1;
  assign popcount22_vqp7_out[1] = input_a[11];
  assign popcount22_vqp7_out[2] = 1'b0;
  assign popcount22_vqp7_out[3] = 1'b1;
  assign popcount22_vqp7_out[4] = 1'b0;
endmodule