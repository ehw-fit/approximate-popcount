// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.70317
// WCE=26.0
// EP=0.968629%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_uhu8(input [26:0] input_a, output [4:0] popcount27_uhu8_out);
  wire popcount27_uhu8_core_030;
  wire popcount27_uhu8_core_031;
  wire popcount27_uhu8_core_032;
  wire popcount27_uhu8_core_034;
  wire popcount27_uhu8_core_038;
  wire popcount27_uhu8_core_040;
  wire popcount27_uhu8_core_044;
  wire popcount27_uhu8_core_045;
  wire popcount27_uhu8_core_046;
  wire popcount27_uhu8_core_048;
  wire popcount27_uhu8_core_049;
  wire popcount27_uhu8_core_051;
  wire popcount27_uhu8_core_056;
  wire popcount27_uhu8_core_057;
  wire popcount27_uhu8_core_058;
  wire popcount27_uhu8_core_061;
  wire popcount27_uhu8_core_063;
  wire popcount27_uhu8_core_066;
  wire popcount27_uhu8_core_069;
  wire popcount27_uhu8_core_071;
  wire popcount27_uhu8_core_073;
  wire popcount27_uhu8_core_076;
  wire popcount27_uhu8_core_077;
  wire popcount27_uhu8_core_078;
  wire popcount27_uhu8_core_080;
  wire popcount27_uhu8_core_081;
  wire popcount27_uhu8_core_082;
  wire popcount27_uhu8_core_083;
  wire popcount27_uhu8_core_084;
  wire popcount27_uhu8_core_085;
  wire popcount27_uhu8_core_087;
  wire popcount27_uhu8_core_088;
  wire popcount27_uhu8_core_092_not;
  wire popcount27_uhu8_core_097;
  wire popcount27_uhu8_core_101;
  wire popcount27_uhu8_core_102;
  wire popcount27_uhu8_core_103;
  wire popcount27_uhu8_core_104;
  wire popcount27_uhu8_core_105;
  wire popcount27_uhu8_core_106;
  wire popcount27_uhu8_core_107;
  wire popcount27_uhu8_core_108;
  wire popcount27_uhu8_core_109;
  wire popcount27_uhu8_core_111;
  wire popcount27_uhu8_core_112;
  wire popcount27_uhu8_core_113;
  wire popcount27_uhu8_core_115;
  wire popcount27_uhu8_core_116;
  wire popcount27_uhu8_core_117;
  wire popcount27_uhu8_core_118;
  wire popcount27_uhu8_core_120;
  wire popcount27_uhu8_core_121;
  wire popcount27_uhu8_core_122;
  wire popcount27_uhu8_core_125;
  wire popcount27_uhu8_core_126;
  wire popcount27_uhu8_core_129;
  wire popcount27_uhu8_core_131;
  wire popcount27_uhu8_core_132;
  wire popcount27_uhu8_core_133;
  wire popcount27_uhu8_core_135;
  wire popcount27_uhu8_core_137;
  wire popcount27_uhu8_core_138;
  wire popcount27_uhu8_core_139;
  wire popcount27_uhu8_core_141;
  wire popcount27_uhu8_core_142;
  wire popcount27_uhu8_core_143;
  wire popcount27_uhu8_core_148;
  wire popcount27_uhu8_core_149;
  wire popcount27_uhu8_core_150;
  wire popcount27_uhu8_core_151;
  wire popcount27_uhu8_core_152;
  wire popcount27_uhu8_core_153;
  wire popcount27_uhu8_core_155;
  wire popcount27_uhu8_core_158;
  wire popcount27_uhu8_core_159;
  wire popcount27_uhu8_core_162;
  wire popcount27_uhu8_core_163;
  wire popcount27_uhu8_core_164;
  wire popcount27_uhu8_core_168;
  wire popcount27_uhu8_core_169;
  wire popcount27_uhu8_core_174;
  wire popcount27_uhu8_core_176;
  wire popcount27_uhu8_core_177_not;
  wire popcount27_uhu8_core_179;
  wire popcount27_uhu8_core_180;
  wire popcount27_uhu8_core_181;
  wire popcount27_uhu8_core_183;
  wire popcount27_uhu8_core_184_not;
  wire popcount27_uhu8_core_185;
  wire popcount27_uhu8_core_188;
  wire popcount27_uhu8_core_189;
  wire popcount27_uhu8_core_190;
  wire popcount27_uhu8_core_192;
  wire popcount27_uhu8_core_193;
  wire popcount27_uhu8_core_194;
  wire popcount27_uhu8_core_195;

  assign popcount27_uhu8_core_030 = input_a[23] & input_a[12];
  assign popcount27_uhu8_core_031 = ~(input_a[8] & input_a[21]);
  assign popcount27_uhu8_core_032 = input_a[3] | input_a[6];
  assign popcount27_uhu8_core_034 = input_a[23] ^ input_a[6];
  assign popcount27_uhu8_core_038 = ~input_a[20];
  assign popcount27_uhu8_core_040 = input_a[2] & input_a[26];
  assign popcount27_uhu8_core_044 = input_a[11] & input_a[7];
  assign popcount27_uhu8_core_045 = ~input_a[1];
  assign popcount27_uhu8_core_046 = input_a[24] & input_a[21];
  assign popcount27_uhu8_core_048 = ~(input_a[20] ^ input_a[6]);
  assign popcount27_uhu8_core_049 = ~input_a[0];
  assign popcount27_uhu8_core_051 = ~input_a[2];
  assign popcount27_uhu8_core_056 = ~(input_a[11] & input_a[21]);
  assign popcount27_uhu8_core_057 = ~(input_a[3] ^ input_a[20]);
  assign popcount27_uhu8_core_058 = ~(input_a[9] & input_a[11]);
  assign popcount27_uhu8_core_061 = ~(input_a[6] ^ input_a[9]);
  assign popcount27_uhu8_core_063 = input_a[7] | input_a[23];
  assign popcount27_uhu8_core_066 = input_a[11] ^ input_a[0];
  assign popcount27_uhu8_core_069 = input_a[6] ^ input_a[20];
  assign popcount27_uhu8_core_071 = input_a[15] | input_a[11];
  assign popcount27_uhu8_core_073 = input_a[24] ^ input_a[14];
  assign popcount27_uhu8_core_076 = input_a[5] ^ input_a[9];
  assign popcount27_uhu8_core_077 = ~input_a[1];
  assign popcount27_uhu8_core_078 = ~(input_a[12] | input_a[5]);
  assign popcount27_uhu8_core_080 = input_a[18] ^ input_a[3];
  assign popcount27_uhu8_core_081 = ~input_a[1];
  assign popcount27_uhu8_core_082 = input_a[12] | input_a[18];
  assign popcount27_uhu8_core_083 = input_a[23] ^ input_a[2];
  assign popcount27_uhu8_core_084 = input_a[19] & input_a[19];
  assign popcount27_uhu8_core_085 = ~input_a[15];
  assign popcount27_uhu8_core_087 = ~input_a[7];
  assign popcount27_uhu8_core_088 = ~(input_a[3] ^ input_a[22]);
  assign popcount27_uhu8_core_092_not = ~input_a[22];
  assign popcount27_uhu8_core_097 = ~(input_a[23] & input_a[3]);
  assign popcount27_uhu8_core_101 = input_a[16] & input_a[7];
  assign popcount27_uhu8_core_102 = ~(input_a[17] | input_a[15]);
  assign popcount27_uhu8_core_103 = input_a[2] ^ input_a[2];
  assign popcount27_uhu8_core_104 = input_a[5] & input_a[4];
  assign popcount27_uhu8_core_105 = input_a[11] & input_a[4];
  assign popcount27_uhu8_core_106 = input_a[4] ^ input_a[6];
  assign popcount27_uhu8_core_107 = ~input_a[11];
  assign popcount27_uhu8_core_108 = input_a[5] ^ input_a[10];
  assign popcount27_uhu8_core_109 = ~(input_a[11] & input_a[25]);
  assign popcount27_uhu8_core_111 = ~(input_a[22] ^ input_a[13]);
  assign popcount27_uhu8_core_112 = ~(input_a[11] | input_a[17]);
  assign popcount27_uhu8_core_113 = input_a[6] ^ input_a[8];
  assign popcount27_uhu8_core_115 = ~(input_a[24] & input_a[23]);
  assign popcount27_uhu8_core_116 = ~(input_a[8] & input_a[7]);
  assign popcount27_uhu8_core_117 = input_a[24] & input_a[19];
  assign popcount27_uhu8_core_118 = ~(input_a[6] ^ input_a[10]);
  assign popcount27_uhu8_core_120 = ~(input_a[14] & input_a[15]);
  assign popcount27_uhu8_core_121 = ~(input_a[2] & input_a[7]);
  assign popcount27_uhu8_core_122 = ~(input_a[15] | input_a[16]);
  assign popcount27_uhu8_core_125 = input_a[13] ^ input_a[14];
  assign popcount27_uhu8_core_126 = ~(input_a[6] ^ input_a[26]);
  assign popcount27_uhu8_core_129 = input_a[24] & input_a[18];
  assign popcount27_uhu8_core_131 = input_a[19] | input_a[5];
  assign popcount27_uhu8_core_132 = ~(input_a[20] | input_a[6]);
  assign popcount27_uhu8_core_133 = input_a[18] & input_a[26];
  assign popcount27_uhu8_core_135 = input_a[6] ^ input_a[22];
  assign popcount27_uhu8_core_137 = ~(input_a[18] ^ input_a[5]);
  assign popcount27_uhu8_core_138 = ~(input_a[1] | input_a[4]);
  assign popcount27_uhu8_core_139 = input_a[10] & input_a[7];
  assign popcount27_uhu8_core_141 = ~(input_a[24] & input_a[5]);
  assign popcount27_uhu8_core_142 = input_a[9] & input_a[5];
  assign popcount27_uhu8_core_143 = input_a[3] | input_a[21];
  assign popcount27_uhu8_core_148 = input_a[16] | input_a[22];
  assign popcount27_uhu8_core_149 = input_a[16] | input_a[7];
  assign popcount27_uhu8_core_150 = ~(input_a[1] & input_a[23]);
  assign popcount27_uhu8_core_151 = input_a[8] ^ input_a[19];
  assign popcount27_uhu8_core_152 = ~(input_a[14] ^ input_a[13]);
  assign popcount27_uhu8_core_153 = input_a[11] | input_a[0];
  assign popcount27_uhu8_core_155 = ~(input_a[14] ^ input_a[8]);
  assign popcount27_uhu8_core_158 = input_a[20] & input_a[5];
  assign popcount27_uhu8_core_159 = input_a[9] ^ input_a[3];
  assign popcount27_uhu8_core_162 = input_a[1] ^ input_a[8];
  assign popcount27_uhu8_core_163 = input_a[21] | input_a[4];
  assign popcount27_uhu8_core_164 = input_a[17] & input_a[9];
  assign popcount27_uhu8_core_168 = ~input_a[25];
  assign popcount27_uhu8_core_169 = input_a[22] | input_a[19];
  assign popcount27_uhu8_core_174 = ~(input_a[8] | input_a[22]);
  assign popcount27_uhu8_core_176 = ~(input_a[2] ^ input_a[3]);
  assign popcount27_uhu8_core_177_not = ~input_a[24];
  assign popcount27_uhu8_core_179 = ~(input_a[14] & input_a[22]);
  assign popcount27_uhu8_core_180 = ~(input_a[4] ^ input_a[2]);
  assign popcount27_uhu8_core_181 = input_a[25] | input_a[3];
  assign popcount27_uhu8_core_183 = input_a[20] ^ input_a[3];
  assign popcount27_uhu8_core_184_not = ~input_a[17];
  assign popcount27_uhu8_core_185 = input_a[0] & input_a[16];
  assign popcount27_uhu8_core_188 = input_a[18] ^ input_a[24];
  assign popcount27_uhu8_core_189 = input_a[22] & input_a[5];
  assign popcount27_uhu8_core_190 = ~(input_a[8] ^ input_a[26]);
  assign popcount27_uhu8_core_192 = ~(input_a[8] | input_a[18]);
  assign popcount27_uhu8_core_193 = ~(input_a[10] & input_a[24]);
  assign popcount27_uhu8_core_194 = ~(input_a[13] | input_a[25]);
  assign popcount27_uhu8_core_195 = ~(input_a[9] ^ input_a[6]);

  assign popcount27_uhu8_out[0] = input_a[10];
  assign popcount27_uhu8_out[1] = input_a[1];
  assign popcount27_uhu8_out[2] = input_a[0];
  assign popcount27_uhu8_out[3] = input_a[16];
  assign popcount27_uhu8_out[4] = input_a[25];
endmodule