// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.63325
// WCE=27.0
// EP=0.971115%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_1j0h(input [30:0] input_a, output [4:0] popcount31_1j0h_out);
  wire popcount31_1j0h_core_033;
  wire popcount31_1j0h_core_037;
  wire popcount31_1j0h_core_040;
  wire popcount31_1j0h_core_041;
  wire popcount31_1j0h_core_043;
  wire popcount31_1j0h_core_044;
  wire popcount31_1j0h_core_045;
  wire popcount31_1j0h_core_047;
  wire popcount31_1j0h_core_049;
  wire popcount31_1j0h_core_052;
  wire popcount31_1j0h_core_053;
  wire popcount31_1j0h_core_056_not;
  wire popcount31_1j0h_core_059;
  wire popcount31_1j0h_core_060;
  wire popcount31_1j0h_core_062;
  wire popcount31_1j0h_core_064;
  wire popcount31_1j0h_core_065;
  wire popcount31_1j0h_core_066;
  wire popcount31_1j0h_core_067;
  wire popcount31_1j0h_core_068;
  wire popcount31_1j0h_core_071;
  wire popcount31_1j0h_core_072;
  wire popcount31_1j0h_core_074;
  wire popcount31_1j0h_core_077;
  wire popcount31_1j0h_core_078;
  wire popcount31_1j0h_core_079;
  wire popcount31_1j0h_core_081;
  wire popcount31_1j0h_core_082;
  wire popcount31_1j0h_core_084;
  wire popcount31_1j0h_core_085;
  wire popcount31_1j0h_core_089;
  wire popcount31_1j0h_core_092;
  wire popcount31_1j0h_core_093;
  wire popcount31_1j0h_core_094;
  wire popcount31_1j0h_core_096;
  wire popcount31_1j0h_core_097;
  wire popcount31_1j0h_core_098;
  wire popcount31_1j0h_core_101;
  wire popcount31_1j0h_core_107;
  wire popcount31_1j0h_core_109;
  wire popcount31_1j0h_core_111;
  wire popcount31_1j0h_core_112;
  wire popcount31_1j0h_core_113;
  wire popcount31_1j0h_core_114;
  wire popcount31_1j0h_core_115;
  wire popcount31_1j0h_core_117;
  wire popcount31_1j0h_core_118;
  wire popcount31_1j0h_core_119;
  wire popcount31_1j0h_core_120;
  wire popcount31_1j0h_core_122;
  wire popcount31_1j0h_core_123;
  wire popcount31_1j0h_core_125;
  wire popcount31_1j0h_core_127;
  wire popcount31_1j0h_core_128;
  wire popcount31_1j0h_core_129;
  wire popcount31_1j0h_core_130;
  wire popcount31_1j0h_core_132;
  wire popcount31_1j0h_core_133;
  wire popcount31_1j0h_core_134;
  wire popcount31_1j0h_core_135;
  wire popcount31_1j0h_core_136;
  wire popcount31_1j0h_core_137;
  wire popcount31_1j0h_core_139;
  wire popcount31_1j0h_core_140;
  wire popcount31_1j0h_core_141;
  wire popcount31_1j0h_core_143;
  wire popcount31_1j0h_core_144;
  wire popcount31_1j0h_core_145;
  wire popcount31_1j0h_core_147;
  wire popcount31_1j0h_core_148;
  wire popcount31_1j0h_core_149;
  wire popcount31_1j0h_core_150;
  wire popcount31_1j0h_core_151;
  wire popcount31_1j0h_core_152;
  wire popcount31_1j0h_core_153;
  wire popcount31_1j0h_core_154;
  wire popcount31_1j0h_core_156;
  wire popcount31_1j0h_core_157;
  wire popcount31_1j0h_core_160;
  wire popcount31_1j0h_core_161;
  wire popcount31_1j0h_core_162;
  wire popcount31_1j0h_core_163;
  wire popcount31_1j0h_core_164;
  wire popcount31_1j0h_core_165;
  wire popcount31_1j0h_core_167;
  wire popcount31_1j0h_core_169;
  wire popcount31_1j0h_core_170;
  wire popcount31_1j0h_core_171;
  wire popcount31_1j0h_core_172;
  wire popcount31_1j0h_core_173_not;
  wire popcount31_1j0h_core_175;
  wire popcount31_1j0h_core_176;
  wire popcount31_1j0h_core_177;
  wire popcount31_1j0h_core_178;
  wire popcount31_1j0h_core_182;
  wire popcount31_1j0h_core_184;
  wire popcount31_1j0h_core_185;
  wire popcount31_1j0h_core_186;
  wire popcount31_1j0h_core_188;
  wire popcount31_1j0h_core_189;
  wire popcount31_1j0h_core_190;
  wire popcount31_1j0h_core_191;
  wire popcount31_1j0h_core_192;
  wire popcount31_1j0h_core_194;
  wire popcount31_1j0h_core_195;
  wire popcount31_1j0h_core_196;
  wire popcount31_1j0h_core_198;
  wire popcount31_1j0h_core_199;
  wire popcount31_1j0h_core_200;
  wire popcount31_1j0h_core_201;
  wire popcount31_1j0h_core_202;
  wire popcount31_1j0h_core_203;
  wire popcount31_1j0h_core_209;
  wire popcount31_1j0h_core_210;
  wire popcount31_1j0h_core_211;
  wire popcount31_1j0h_core_215_not;
  wire popcount31_1j0h_core_216;
  wire popcount31_1j0h_core_217;
  wire popcount31_1j0h_core_218;
  wire popcount31_1j0h_core_219;

  assign popcount31_1j0h_core_033 = ~(input_a[25] & input_a[8]);
  assign popcount31_1j0h_core_037 = ~(input_a[2] ^ input_a[12]);
  assign popcount31_1j0h_core_040 = ~(input_a[20] | input_a[6]);
  assign popcount31_1j0h_core_041 = ~(input_a[22] ^ input_a[16]);
  assign popcount31_1j0h_core_043 = ~(input_a[24] | input_a[9]);
  assign popcount31_1j0h_core_044 = input_a[17] & input_a[1];
  assign popcount31_1j0h_core_045 = input_a[28] ^ input_a[2];
  assign popcount31_1j0h_core_047 = input_a[4] | input_a[22];
  assign popcount31_1j0h_core_049 = ~(input_a[19] & input_a[7]);
  assign popcount31_1j0h_core_052 = ~(input_a[12] ^ input_a[8]);
  assign popcount31_1j0h_core_053 = ~input_a[14];
  assign popcount31_1j0h_core_056_not = ~input_a[25];
  assign popcount31_1j0h_core_059 = input_a[7] & input_a[24];
  assign popcount31_1j0h_core_060 = ~(input_a[14] ^ input_a[1]);
  assign popcount31_1j0h_core_062 = ~(input_a[11] ^ input_a[5]);
  assign popcount31_1j0h_core_064 = ~input_a[8];
  assign popcount31_1j0h_core_065 = ~(input_a[5] | input_a[22]);
  assign popcount31_1j0h_core_066 = ~(input_a[6] | input_a[10]);
  assign popcount31_1j0h_core_067 = ~(input_a[0] | input_a[21]);
  assign popcount31_1j0h_core_068 = input_a[30] ^ input_a[28];
  assign popcount31_1j0h_core_071 = ~(input_a[26] | input_a[8]);
  assign popcount31_1j0h_core_072 = input_a[14] | input_a[26];
  assign popcount31_1j0h_core_074 = input_a[5] & input_a[28];
  assign popcount31_1j0h_core_077 = ~(input_a[26] | input_a[18]);
  assign popcount31_1j0h_core_078 = input_a[22] & input_a[27];
  assign popcount31_1j0h_core_079 = ~input_a[9];
  assign popcount31_1j0h_core_081 = input_a[27] | input_a[9];
  assign popcount31_1j0h_core_082 = ~(input_a[2] & input_a[30]);
  assign popcount31_1j0h_core_084 = input_a[18] ^ input_a[2];
  assign popcount31_1j0h_core_085 = input_a[20] & input_a[14];
  assign popcount31_1j0h_core_089 = ~input_a[0];
  assign popcount31_1j0h_core_092 = ~(input_a[26] | input_a[8]);
  assign popcount31_1j0h_core_093 = input_a[14] ^ input_a[22];
  assign popcount31_1j0h_core_094 = input_a[3] | input_a[2];
  assign popcount31_1j0h_core_096 = ~(input_a[30] & input_a[10]);
  assign popcount31_1j0h_core_097 = ~input_a[19];
  assign popcount31_1j0h_core_098 = input_a[5] & input_a[0];
  assign popcount31_1j0h_core_101 = input_a[19] ^ input_a[17];
  assign popcount31_1j0h_core_107 = input_a[18] | input_a[8];
  assign popcount31_1j0h_core_109 = ~(input_a[24] | input_a[9]);
  assign popcount31_1j0h_core_111 = input_a[23] & input_a[21];
  assign popcount31_1j0h_core_112 = input_a[26] ^ input_a[20];
  assign popcount31_1j0h_core_113 = input_a[15] | input_a[30];
  assign popcount31_1j0h_core_114 = ~(input_a[9] | input_a[13]);
  assign popcount31_1j0h_core_115 = ~(input_a[19] & input_a[20]);
  assign popcount31_1j0h_core_117 = ~(input_a[19] & input_a[30]);
  assign popcount31_1j0h_core_118 = ~(input_a[7] | input_a[13]);
  assign popcount31_1j0h_core_119 = ~(input_a[8] ^ input_a[23]);
  assign popcount31_1j0h_core_120 = input_a[12] & input_a[1];
  assign popcount31_1j0h_core_122 = input_a[16] & input_a[11];
  assign popcount31_1j0h_core_123 = ~(input_a[5] | input_a[25]);
  assign popcount31_1j0h_core_125 = input_a[30] & input_a[4];
  assign popcount31_1j0h_core_127 = input_a[20] ^ input_a[20];
  assign popcount31_1j0h_core_128 = ~(input_a[2] | input_a[2]);
  assign popcount31_1j0h_core_129 = ~(input_a[10] & input_a[16]);
  assign popcount31_1j0h_core_130 = ~(input_a[3] | input_a[13]);
  assign popcount31_1j0h_core_132 = input_a[5] ^ input_a[2];
  assign popcount31_1j0h_core_133 = input_a[14] | input_a[20];
  assign popcount31_1j0h_core_134 = ~(input_a[19] ^ input_a[11]);
  assign popcount31_1j0h_core_135 = input_a[1] | input_a[18];
  assign popcount31_1j0h_core_136 = ~input_a[7];
  assign popcount31_1j0h_core_137 = input_a[1] | input_a[4];
  assign popcount31_1j0h_core_139 = ~(input_a[4] | input_a[26]);
  assign popcount31_1j0h_core_140 = ~(input_a[19] & input_a[17]);
  assign popcount31_1j0h_core_141 = ~(input_a[7] | input_a[10]);
  assign popcount31_1j0h_core_143 = input_a[19] ^ input_a[23];
  assign popcount31_1j0h_core_144 = input_a[16] | input_a[11];
  assign popcount31_1j0h_core_145 = ~(input_a[21] | input_a[18]);
  assign popcount31_1j0h_core_147 = ~(input_a[29] & input_a[25]);
  assign popcount31_1j0h_core_148 = ~(input_a[6] ^ input_a[20]);
  assign popcount31_1j0h_core_149 = ~input_a[28];
  assign popcount31_1j0h_core_150 = ~input_a[22];
  assign popcount31_1j0h_core_151 = ~input_a[5];
  assign popcount31_1j0h_core_152 = input_a[8] & input_a[8];
  assign popcount31_1j0h_core_153 = ~(input_a[24] ^ input_a[2]);
  assign popcount31_1j0h_core_154 = ~(input_a[20] & input_a[10]);
  assign popcount31_1j0h_core_156 = ~input_a[21];
  assign popcount31_1j0h_core_157 = ~(input_a[18] | input_a[26]);
  assign popcount31_1j0h_core_160 = ~(input_a[4] & input_a[26]);
  assign popcount31_1j0h_core_161 = input_a[26] ^ input_a[23];
  assign popcount31_1j0h_core_162 = input_a[26] & input_a[8];
  assign popcount31_1j0h_core_163 = ~input_a[2];
  assign popcount31_1j0h_core_164 = ~input_a[7];
  assign popcount31_1j0h_core_165 = ~(input_a[0] ^ input_a[0]);
  assign popcount31_1j0h_core_167 = ~(input_a[23] | input_a[9]);
  assign popcount31_1j0h_core_169 = ~(input_a[5] | input_a[7]);
  assign popcount31_1j0h_core_170 = input_a[1] | input_a[7];
  assign popcount31_1j0h_core_171 = input_a[11] | input_a[12];
  assign popcount31_1j0h_core_172 = ~(input_a[11] & input_a[30]);
  assign popcount31_1j0h_core_173_not = ~input_a[19];
  assign popcount31_1j0h_core_175 = ~(input_a[29] ^ input_a[14]);
  assign popcount31_1j0h_core_176 = ~input_a[16];
  assign popcount31_1j0h_core_177 = ~(input_a[2] & input_a[26]);
  assign popcount31_1j0h_core_178 = input_a[1] | input_a[9];
  assign popcount31_1j0h_core_182 = input_a[16] | input_a[12];
  assign popcount31_1j0h_core_184 = ~(input_a[3] | input_a[20]);
  assign popcount31_1j0h_core_185 = ~(input_a[3] | input_a[28]);
  assign popcount31_1j0h_core_186 = ~(input_a[30] | input_a[4]);
  assign popcount31_1j0h_core_188 = ~(input_a[24] | input_a[21]);
  assign popcount31_1j0h_core_189 = input_a[16] | input_a[1];
  assign popcount31_1j0h_core_190 = input_a[1] | input_a[6];
  assign popcount31_1j0h_core_191 = input_a[5] | input_a[12];
  assign popcount31_1j0h_core_192 = ~(input_a[22] | input_a[10]);
  assign popcount31_1j0h_core_194 = ~(input_a[13] & input_a[8]);
  assign popcount31_1j0h_core_195 = ~(input_a[30] | input_a[20]);
  assign popcount31_1j0h_core_196 = input_a[8] ^ input_a[25];
  assign popcount31_1j0h_core_198 = ~(input_a[1] ^ input_a[19]);
  assign popcount31_1j0h_core_199 = ~(input_a[13] | input_a[28]);
  assign popcount31_1j0h_core_200 = input_a[12] | input_a[12];
  assign popcount31_1j0h_core_201 = ~(input_a[23] | input_a[19]);
  assign popcount31_1j0h_core_202 = ~(input_a[8] ^ input_a[27]);
  assign popcount31_1j0h_core_203 = ~(input_a[15] & input_a[19]);
  assign popcount31_1j0h_core_209 = ~(input_a[13] | input_a[25]);
  assign popcount31_1j0h_core_210 = input_a[4] | input_a[1];
  assign popcount31_1j0h_core_211 = ~(input_a[1] | input_a[8]);
  assign popcount31_1j0h_core_215_not = ~input_a[23];
  assign popcount31_1j0h_core_216 = input_a[24] | input_a[22];
  assign popcount31_1j0h_core_217 = input_a[0] ^ input_a[22];
  assign popcount31_1j0h_core_218 = ~(input_a[5] | input_a[20]);
  assign popcount31_1j0h_core_219 = ~(input_a[28] & input_a[18]);

  assign popcount31_1j0h_out[0] = 1'b0;
  assign popcount31_1j0h_out[1] = input_a[8];
  assign popcount31_1j0h_out[2] = input_a[27];
  assign popcount31_1j0h_out[3] = input_a[0];
  assign popcount31_1j0h_out[4] = 1'b1;
endmodule