// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.89695
// WCE=21.0
// EP=0.835582%
// Printed PDK parameters:
//  Area=52216272.0
//  Delay=70459976.0
//  Power=2494900.0

module popcount38_debw(input [37:0] input_a, output [5:0] popcount38_debw_out);
  wire popcount38_debw_core_041;
  wire popcount38_debw_core_042;
  wire popcount38_debw_core_043;
  wire popcount38_debw_core_045;
  wire popcount38_debw_core_046;
  wire popcount38_debw_core_047;
  wire popcount38_debw_core_049;
  wire popcount38_debw_core_051;
  wire popcount38_debw_core_054;
  wire popcount38_debw_core_055;
  wire popcount38_debw_core_059;
  wire popcount38_debw_core_060;
  wire popcount38_debw_core_061;
  wire popcount38_debw_core_062;
  wire popcount38_debw_core_063;
  wire popcount38_debw_core_064;
  wire popcount38_debw_core_065;
  wire popcount38_debw_core_069;
  wire popcount38_debw_core_070;
  wire popcount38_debw_core_071;
  wire popcount38_debw_core_073;
  wire popcount38_debw_core_075;
  wire popcount38_debw_core_077;
  wire popcount38_debw_core_081;
  wire popcount38_debw_core_082;
  wire popcount38_debw_core_083;
  wire popcount38_debw_core_085;
  wire popcount38_debw_core_086;
  wire popcount38_debw_core_087;
  wire popcount38_debw_core_088;
  wire popcount38_debw_core_092;
  wire popcount38_debw_core_093;
  wire popcount38_debw_core_094;
  wire popcount38_debw_core_095;
  wire popcount38_debw_core_096;
  wire popcount38_debw_core_098;
  wire popcount38_debw_core_099;
  wire popcount38_debw_core_100;
  wire popcount38_debw_core_101;
  wire popcount38_debw_core_102;
  wire popcount38_debw_core_104;
  wire popcount38_debw_core_105;
  wire popcount38_debw_core_106;
  wire popcount38_debw_core_107;
  wire popcount38_debw_core_109;
  wire popcount38_debw_core_110;
  wire popcount38_debw_core_111;
  wire popcount38_debw_core_112;
  wire popcount38_debw_core_113;
  wire popcount38_debw_core_114;
  wire popcount38_debw_core_115;
  wire popcount38_debw_core_116;
  wire popcount38_debw_core_117;
  wire popcount38_debw_core_118;
  wire popcount38_debw_core_119;
  wire popcount38_debw_core_120;
  wire popcount38_debw_core_121;
  wire popcount38_debw_core_122;
  wire popcount38_debw_core_123;
  wire popcount38_debw_core_124;
  wire popcount38_debw_core_125;
  wire popcount38_debw_core_126;
  wire popcount38_debw_core_127;
  wire popcount38_debw_core_129;
  wire popcount38_debw_core_132;
  wire popcount38_debw_core_133;
  wire popcount38_debw_core_134;
  wire popcount38_debw_core_135_not;
  wire popcount38_debw_core_138;
  wire popcount38_debw_core_140;
  wire popcount38_debw_core_141;
  wire popcount38_debw_core_142;
  wire popcount38_debw_core_143;
  wire popcount38_debw_core_144;
  wire popcount38_debw_core_147;
  wire popcount38_debw_core_151;
  wire popcount38_debw_core_154;
  wire popcount38_debw_core_155;
  wire popcount38_debw_core_156;
  wire popcount38_debw_core_157;
  wire popcount38_debw_core_159;
  wire popcount38_debw_core_161;
  wire popcount38_debw_core_162;
  wire popcount38_debw_core_163_not;
  wire popcount38_debw_core_164;
  wire popcount38_debw_core_165;
  wire popcount38_debw_core_166;
  wire popcount38_debw_core_167;
  wire popcount38_debw_core_168;
  wire popcount38_debw_core_170;
  wire popcount38_debw_core_171;
  wire popcount38_debw_core_173;
  wire popcount38_debw_core_174;
  wire popcount38_debw_core_175;
  wire popcount38_debw_core_176;
  wire popcount38_debw_core_177;
  wire popcount38_debw_core_178;
  wire popcount38_debw_core_179;
  wire popcount38_debw_core_184;
  wire popcount38_debw_core_185;
  wire popcount38_debw_core_186;
  wire popcount38_debw_core_188;
  wire popcount38_debw_core_189;
  wire popcount38_debw_core_190;
  wire popcount38_debw_core_191;
  wire popcount38_debw_core_193;
  wire popcount38_debw_core_194;
  wire popcount38_debw_core_197;
  wire popcount38_debw_core_198;
  wire popcount38_debw_core_200;
  wire popcount38_debw_core_201;
  wire popcount38_debw_core_202;
  wire popcount38_debw_core_203;
  wire popcount38_debw_core_205;
  wire popcount38_debw_core_209;
  wire popcount38_debw_core_210;
  wire popcount38_debw_core_214;
  wire popcount38_debw_core_215;
  wire popcount38_debw_core_216;
  wire popcount38_debw_core_217;
  wire popcount38_debw_core_218;
  wire popcount38_debw_core_219;
  wire popcount38_debw_core_220;
  wire popcount38_debw_core_222;
  wire popcount38_debw_core_223;
  wire popcount38_debw_core_224;
  wire popcount38_debw_core_225;
  wire popcount38_debw_core_226;
  wire popcount38_debw_core_227;
  wire popcount38_debw_core_228;
  wire popcount38_debw_core_230;
  wire popcount38_debw_core_232;
  wire popcount38_debw_core_233;
  wire popcount38_debw_core_234;
  wire popcount38_debw_core_235;
  wire popcount38_debw_core_236;
  wire popcount38_debw_core_237;
  wire popcount38_debw_core_238;
  wire popcount38_debw_core_239;
  wire popcount38_debw_core_240;
  wire popcount38_debw_core_242;
  wire popcount38_debw_core_244;
  wire popcount38_debw_core_247;
  wire popcount38_debw_core_248;
  wire popcount38_debw_core_249;
  wire popcount38_debw_core_251;
  wire popcount38_debw_core_253;
  wire popcount38_debw_core_254;
  wire popcount38_debw_core_255_not;
  wire popcount38_debw_core_258;
  wire popcount38_debw_core_262;
  wire popcount38_debw_core_263_not;
  wire popcount38_debw_core_264;
  wire popcount38_debw_core_265;
  wire popcount38_debw_core_266;
  wire popcount38_debw_core_268;
  wire popcount38_debw_core_269;
  wire popcount38_debw_core_270;
  wire popcount38_debw_core_271;
  wire popcount38_debw_core_272;
  wire popcount38_debw_core_273;
  wire popcount38_debw_core_274;
  wire popcount38_debw_core_275;
  wire popcount38_debw_core_276;
  wire popcount38_debw_core_277;
  wire popcount38_debw_core_278;
  wire popcount38_debw_core_279;
  wire popcount38_debw_core_280;
  wire popcount38_debw_core_281;
  wire popcount38_debw_core_282;
  wire popcount38_debw_core_283;
  wire popcount38_debw_core_284;
  wire popcount38_debw_core_285;
  wire popcount38_debw_core_286;
  wire popcount38_debw_core_288;
  wire popcount38_debw_core_289;
  wire popcount38_debw_core_291;
  wire popcount38_debw_core_293;
  wire popcount38_debw_core_294;
  wire popcount38_debw_core_295;

  assign popcount38_debw_core_041 = input_a[11] & input_a[3];
  assign popcount38_debw_core_042 = ~(input_a[12] | input_a[20]);
  assign popcount38_debw_core_043 = input_a[20] & input_a[23];
  assign popcount38_debw_core_045 = ~(input_a[30] ^ input_a[37]);
  assign popcount38_debw_core_046 = popcount38_debw_core_041 | popcount38_debw_core_043;
  assign popcount38_debw_core_047 = popcount38_debw_core_041 & input_a[12];
  assign popcount38_debw_core_049 = ~input_a[33];
  assign popcount38_debw_core_051 = input_a[20] | input_a[27];
  assign popcount38_debw_core_054 = ~(input_a[23] | input_a[28]);
  assign popcount38_debw_core_055 = input_a[0] | input_a[6];
  assign popcount38_debw_core_059 = input_a[35] | input_a[3];
  assign popcount38_debw_core_060 = input_a[37] & input_a[18];
  assign popcount38_debw_core_061 = ~(input_a[28] | input_a[36]);
  assign popcount38_debw_core_062 = input_a[7] & input_a[21];
  assign popcount38_debw_core_063 = ~(input_a[15] | input_a[32]);
  assign popcount38_debw_core_064 = input_a[22] & input_a[5];
  assign popcount38_debw_core_065 = popcount38_debw_core_062 | popcount38_debw_core_064;
  assign popcount38_debw_core_069 = ~(input_a[30] | input_a[11]);
  assign popcount38_debw_core_070 = ~input_a[2];
  assign popcount38_debw_core_071 = popcount38_debw_core_046 & input_a[1];
  assign popcount38_debw_core_073 = input_a[32] ^ input_a[4];
  assign popcount38_debw_core_075 = popcount38_debw_core_047 | popcount38_debw_core_065;
  assign popcount38_debw_core_077 = popcount38_debw_core_075 | popcount38_debw_core_071;
  assign popcount38_debw_core_081 = ~(input_a[12] & input_a[18]);
  assign popcount38_debw_core_082 = input_a[9] ^ input_a[10];
  assign popcount38_debw_core_083 = input_a[9] & input_a[10];
  assign popcount38_debw_core_085 = input_a[6] & input_a[26];
  assign popcount38_debw_core_086 = ~(input_a[1] | input_a[35]);
  assign popcount38_debw_core_087 = input_a[4] & input_a[25];
  assign popcount38_debw_core_088 = popcount38_debw_core_085 | popcount38_debw_core_087;
  assign popcount38_debw_core_092 = popcount38_debw_core_083 ^ popcount38_debw_core_088;
  assign popcount38_debw_core_093 = input_a[10] & popcount38_debw_core_088;
  assign popcount38_debw_core_094 = popcount38_debw_core_092 ^ popcount38_debw_core_082;
  assign popcount38_debw_core_095 = popcount38_debw_core_092 & popcount38_debw_core_082;
  assign popcount38_debw_core_096 = popcount38_debw_core_093 | popcount38_debw_core_095;
  assign popcount38_debw_core_098 = input_a[36] | input_a[18];
  assign popcount38_debw_core_099 = input_a[14] ^ input_a[15];
  assign popcount38_debw_core_100 = input_a[14] & input_a[15];
  assign popcount38_debw_core_101 = input_a[32] & input_a[18];
  assign popcount38_debw_core_102 = input_a[29] & input_a[13];
  assign popcount38_debw_core_104 = input_a[16] & popcount38_debw_core_101;
  assign popcount38_debw_core_105 = popcount38_debw_core_102 | popcount38_debw_core_104;
  assign popcount38_debw_core_106 = popcount38_debw_core_102 & popcount38_debw_core_104;
  assign popcount38_debw_core_107 = ~popcount38_debw_core_099;
  assign popcount38_debw_core_109 = popcount38_debw_core_100 ^ popcount38_debw_core_105;
  assign popcount38_debw_core_110 = input_a[15] & popcount38_debw_core_105;
  assign popcount38_debw_core_111 = popcount38_debw_core_109 ^ popcount38_debw_core_099;
  assign popcount38_debw_core_112 = popcount38_debw_core_109 & popcount38_debw_core_099;
  assign popcount38_debw_core_113 = popcount38_debw_core_110 | popcount38_debw_core_112;
  assign popcount38_debw_core_114 = popcount38_debw_core_106 | popcount38_debw_core_113;
  assign popcount38_debw_core_115 = input_a[29] & input_a[19];
  assign popcount38_debw_core_116 = ~(input_a[13] | input_a[7]);
  assign popcount38_debw_core_117 = input_a[30] & popcount38_debw_core_107;
  assign popcount38_debw_core_118 = popcount38_debw_core_094 ^ popcount38_debw_core_111;
  assign popcount38_debw_core_119 = popcount38_debw_core_094 & popcount38_debw_core_111;
  assign popcount38_debw_core_120 = popcount38_debw_core_118 ^ popcount38_debw_core_117;
  assign popcount38_debw_core_121 = popcount38_debw_core_118 & popcount38_debw_core_117;
  assign popcount38_debw_core_122 = popcount38_debw_core_119 | popcount38_debw_core_121;
  assign popcount38_debw_core_123 = popcount38_debw_core_096 ^ popcount38_debw_core_114;
  assign popcount38_debw_core_124 = popcount38_debw_core_096 & popcount38_debw_core_114;
  assign popcount38_debw_core_125 = popcount38_debw_core_123 ^ popcount38_debw_core_122;
  assign popcount38_debw_core_126 = popcount38_debw_core_123 & popcount38_debw_core_122;
  assign popcount38_debw_core_127 = popcount38_debw_core_124 | popcount38_debw_core_126;
  assign popcount38_debw_core_129 = input_a[24] & input_a[1];
  assign popcount38_debw_core_132 = input_a[35] ^ input_a[19];
  assign popcount38_debw_core_133 = ~input_a[33];
  assign popcount38_debw_core_134 = ~input_a[9];
  assign popcount38_debw_core_135_not = ~popcount38_debw_core_120;
  assign popcount38_debw_core_138 = ~(input_a[25] ^ input_a[17]);
  assign popcount38_debw_core_140 = popcount38_debw_core_077 ^ popcount38_debw_core_125;
  assign popcount38_debw_core_141 = popcount38_debw_core_077 & popcount38_debw_core_125;
  assign popcount38_debw_core_142 = popcount38_debw_core_140 ^ popcount38_debw_core_120;
  assign popcount38_debw_core_143 = popcount38_debw_core_140 & popcount38_debw_core_120;
  assign popcount38_debw_core_144 = popcount38_debw_core_141 | popcount38_debw_core_143;
  assign popcount38_debw_core_147 = popcount38_debw_core_127 ^ popcount38_debw_core_144;
  assign popcount38_debw_core_151 = ~(input_a[37] & input_a[12]);
  assign popcount38_debw_core_154 = ~(input_a[17] ^ input_a[15]);
  assign popcount38_debw_core_155 = ~(input_a[25] | input_a[36]);
  assign popcount38_debw_core_156 = input_a[0] | input_a[28];
  assign popcount38_debw_core_157 = ~(input_a[30] | input_a[13]);
  assign popcount38_debw_core_159 = input_a[6] & input_a[0];
  assign popcount38_debw_core_161 = ~(input_a[32] ^ input_a[23]);
  assign popcount38_debw_core_162 = ~input_a[35];
  assign popcount38_debw_core_163_not = ~input_a[19];
  assign popcount38_debw_core_164 = ~(input_a[16] & input_a[31]);
  assign popcount38_debw_core_165 = input_a[24] ^ input_a[15];
  assign popcount38_debw_core_166 = ~(input_a[18] ^ input_a[5]);
  assign popcount38_debw_core_167 = input_a[28] & input_a[25];
  assign popcount38_debw_core_168 = ~(input_a[27] | input_a[17]);
  assign popcount38_debw_core_170 = ~(input_a[35] ^ input_a[2]);
  assign popcount38_debw_core_171 = ~(input_a[22] & input_a[16]);
  assign popcount38_debw_core_173 = input_a[17] ^ input_a[33];
  assign popcount38_debw_core_174 = input_a[3] ^ input_a[6];
  assign popcount38_debw_core_175 = input_a[3] | input_a[27];
  assign popcount38_debw_core_176 = ~input_a[11];
  assign popcount38_debw_core_177 = input_a[34] & input_a[32];
  assign popcount38_debw_core_178 = ~(input_a[30] | input_a[5]);
  assign popcount38_debw_core_179 = ~input_a[15];
  assign popcount38_debw_core_184 = ~input_a[5];
  assign popcount38_debw_core_185 = ~(input_a[11] ^ input_a[5]);
  assign popcount38_debw_core_186 = input_a[36] | input_a[36];
  assign popcount38_debw_core_188 = ~(input_a[30] ^ input_a[18]);
  assign popcount38_debw_core_189 = ~(input_a[5] ^ input_a[34]);
  assign popcount38_debw_core_190 = input_a[13] & input_a[10];
  assign popcount38_debw_core_191 = ~(input_a[3] ^ input_a[13]);
  assign popcount38_debw_core_193 = input_a[25] & input_a[24];
  assign popcount38_debw_core_194 = input_a[9] & input_a[20];
  assign popcount38_debw_core_197 = ~(input_a[12] & input_a[23]);
  assign popcount38_debw_core_198 = ~(input_a[7] & input_a[11]);
  assign popcount38_debw_core_200 = ~(input_a[34] | input_a[26]);
  assign popcount38_debw_core_201 = ~(input_a[13] & input_a[18]);
  assign popcount38_debw_core_202 = ~(input_a[31] | input_a[2]);
  assign popcount38_debw_core_203 = input_a[1] | input_a[30];
  assign popcount38_debw_core_205 = ~(input_a[24] | input_a[14]);
  assign popcount38_debw_core_209 = ~(input_a[31] & input_a[0]);
  assign popcount38_debw_core_210 = input_a[31] & input_a[0];
  assign popcount38_debw_core_214 = input_a[33] ^ input_a[34];
  assign popcount38_debw_core_215 = input_a[33] & input_a[34];
  assign popcount38_debw_core_216 = input_a[36] ^ input_a[37];
  assign popcount38_debw_core_217 = input_a[36] & input_a[37];
  assign popcount38_debw_core_218 = input_a[35] ^ popcount38_debw_core_216;
  assign popcount38_debw_core_219 = input_a[35] & popcount38_debw_core_216;
  assign popcount38_debw_core_220 = popcount38_debw_core_217 | popcount38_debw_core_219;
  assign popcount38_debw_core_222 = input_a[36] | popcount38_debw_core_218;
  assign popcount38_debw_core_223 = popcount38_debw_core_214 & popcount38_debw_core_218;
  assign popcount38_debw_core_224 = popcount38_debw_core_215 ^ popcount38_debw_core_220;
  assign popcount38_debw_core_225 = popcount38_debw_core_215 & popcount38_debw_core_220;
  assign popcount38_debw_core_226 = popcount38_debw_core_224 ^ popcount38_debw_core_223;
  assign popcount38_debw_core_227 = popcount38_debw_core_224 & popcount38_debw_core_223;
  assign popcount38_debw_core_228 = popcount38_debw_core_225 | popcount38_debw_core_227;
  assign popcount38_debw_core_230 = input_a[20] ^ input_a[22];
  assign popcount38_debw_core_232 = input_a[19] & input_a[28];
  assign popcount38_debw_core_233 = popcount38_debw_core_209 ^ popcount38_debw_core_226;
  assign popcount38_debw_core_234 = popcount38_debw_core_209 & popcount38_debw_core_226;
  assign popcount38_debw_core_235 = popcount38_debw_core_233 ^ popcount38_debw_core_232;
  assign popcount38_debw_core_236 = popcount38_debw_core_233 & popcount38_debw_core_232;
  assign popcount38_debw_core_237 = popcount38_debw_core_234 | popcount38_debw_core_236;
  assign popcount38_debw_core_238 = popcount38_debw_core_210 ^ popcount38_debw_core_228;
  assign popcount38_debw_core_239 = input_a[31] & input_a[0];
  assign popcount38_debw_core_240 = popcount38_debw_core_238 ^ popcount38_debw_core_237;
  assign popcount38_debw_core_242 = popcount38_debw_core_239 | popcount38_debw_core_238;
  assign popcount38_debw_core_244 = ~(input_a[0] & input_a[8]);
  assign popcount38_debw_core_247 = ~input_a[27];
  assign popcount38_debw_core_248 = ~input_a[21];
  assign popcount38_debw_core_249 = ~input_a[34];
  assign popcount38_debw_core_251 = input_a[0] | input_a[22];
  assign popcount38_debw_core_253 = ~(input_a[5] & input_a[6]);
  assign popcount38_debw_core_254 = input_a[28] & input_a[5];
  assign popcount38_debw_core_255_not = ~popcount38_debw_core_240;
  assign popcount38_debw_core_258 = ~(input_a[20] ^ input_a[14]);
  assign popcount38_debw_core_262 = popcount38_debw_core_242 | popcount38_debw_core_240;
  assign popcount38_debw_core_263_not = ~input_a[34];
  assign popcount38_debw_core_264 = input_a[19] ^ input_a[5];
  assign popcount38_debw_core_265 = input_a[35] ^ input_a[9];
  assign popcount38_debw_core_266 = ~input_a[22];
  assign popcount38_debw_core_268 = input_a[24] ^ input_a[3];
  assign popcount38_debw_core_269 = ~(input_a[0] | input_a[37]);
  assign popcount38_debw_core_270 = ~(input_a[5] & input_a[8]);
  assign popcount38_debw_core_271 = input_a[8] & input_a[24];
  assign popcount38_debw_core_272 = popcount38_debw_core_135_not ^ popcount38_debw_core_235;
  assign popcount38_debw_core_273 = popcount38_debw_core_135_not & popcount38_debw_core_235;
  assign popcount38_debw_core_274 = popcount38_debw_core_272 ^ popcount38_debw_core_271;
  assign popcount38_debw_core_275 = popcount38_debw_core_272 & popcount38_debw_core_271;
  assign popcount38_debw_core_276 = popcount38_debw_core_273 | popcount38_debw_core_275;
  assign popcount38_debw_core_277 = popcount38_debw_core_142 ^ popcount38_debw_core_255_not;
  assign popcount38_debw_core_278 = popcount38_debw_core_142 & popcount38_debw_core_255_not;
  assign popcount38_debw_core_279 = popcount38_debw_core_277 ^ popcount38_debw_core_276;
  assign popcount38_debw_core_280 = popcount38_debw_core_277 & popcount38_debw_core_276;
  assign popcount38_debw_core_281 = popcount38_debw_core_278 | popcount38_debw_core_280;
  assign popcount38_debw_core_282 = popcount38_debw_core_147 ^ popcount38_debw_core_262;
  assign popcount38_debw_core_283 = popcount38_debw_core_147 & popcount38_debw_core_262;
  assign popcount38_debw_core_284 = popcount38_debw_core_282 ^ popcount38_debw_core_281;
  assign popcount38_debw_core_285 = popcount38_debw_core_282 & popcount38_debw_core_281;
  assign popcount38_debw_core_286 = popcount38_debw_core_283 | popcount38_debw_core_285;
  assign popcount38_debw_core_288 = ~(input_a[13] & input_a[15]);
  assign popcount38_debw_core_289 = popcount38_debw_core_127 | popcount38_debw_core_286;
  assign popcount38_debw_core_291 = ~(input_a[27] ^ input_a[9]);
  assign popcount38_debw_core_293 = input_a[36] & input_a[2];
  assign popcount38_debw_core_294 = ~(input_a[26] | input_a[15]);
  assign popcount38_debw_core_295 = input_a[2] ^ input_a[24];

  assign popcount38_debw_out[0] = popcount38_debw_core_282;
  assign popcount38_debw_out[1] = popcount38_debw_core_274;
  assign popcount38_debw_out[2] = popcount38_debw_core_279;
  assign popcount38_debw_out[3] = popcount38_debw_core_284;
  assign popcount38_debw_out[4] = popcount38_debw_core_289;
  assign popcount38_debw_out[5] = 1'b0;
endmodule