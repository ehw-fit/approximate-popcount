// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.59907
// WCE=13.0
// EP=0.806548%
// Printed PDK parameters:
//  Area=53426718.0
//  Delay=72147680.0
//  Power=2534600.0

module popcount32_iick(input [31:0] input_a, output [5:0] popcount32_iick_out);
  wire popcount32_iick_core_035;
  wire popcount32_iick_core_036;
  wire popcount32_iick_core_038;
  wire popcount32_iick_core_040;
  wire popcount32_iick_core_041;
  wire popcount32_iick_core_042;
  wire popcount32_iick_core_043;
  wire popcount32_iick_core_045;
  wire popcount32_iick_core_046;
  wire popcount32_iick_core_049;
  wire popcount32_iick_core_051;
  wire popcount32_iick_core_052;
  wire popcount32_iick_core_053;
  wire popcount32_iick_core_056;
  wire popcount32_iick_core_058;
  wire popcount32_iick_core_059;
  wire popcount32_iick_core_061;
  wire popcount32_iick_core_064;
  wire popcount32_iick_core_065;
  wire popcount32_iick_core_066;
  wire popcount32_iick_core_068;
  wire popcount32_iick_core_069;
  wire popcount32_iick_core_070;
  wire popcount32_iick_core_072;
  wire popcount32_iick_core_074;
  wire popcount32_iick_core_075;
  wire popcount32_iick_core_076;
  wire popcount32_iick_core_077;
  wire popcount32_iick_core_078;
  wire popcount32_iick_core_079;
  wire popcount32_iick_core_080;
  wire popcount32_iick_core_081;
  wire popcount32_iick_core_082;
  wire popcount32_iick_core_083;
  wire popcount32_iick_core_084;
  wire popcount32_iick_core_085;
  wire popcount32_iick_core_086;
  wire popcount32_iick_core_087;
  wire popcount32_iick_core_088;
  wire popcount32_iick_core_089;
  wire popcount32_iick_core_091;
  wire popcount32_iick_core_092;
  wire popcount32_iick_core_093;
  wire popcount32_iick_core_094;
  wire popcount32_iick_core_095;
  wire popcount32_iick_core_096;
  wire popcount32_iick_core_097;
  wire popcount32_iick_core_098;
  wire popcount32_iick_core_099;
  wire popcount32_iick_core_100;
  wire popcount32_iick_core_101;
  wire popcount32_iick_core_103;
  wire popcount32_iick_core_104;
  wire popcount32_iick_core_105;
  wire popcount32_iick_core_106;
  wire popcount32_iick_core_109;
  wire popcount32_iick_core_110;
  wire popcount32_iick_core_111;
  wire popcount32_iick_core_112;
  wire popcount32_iick_core_113;
  wire popcount32_iick_core_115_not;
  wire popcount32_iick_core_116;
  wire popcount32_iick_core_118;
  wire popcount32_iick_core_119;
  wire popcount32_iick_core_120;
  wire popcount32_iick_core_121;
  wire popcount32_iick_core_122;
  wire popcount32_iick_core_123;
  wire popcount32_iick_core_125;
  wire popcount32_iick_core_126;
  wire popcount32_iick_core_127;
  wire popcount32_iick_core_130;
  wire popcount32_iick_core_131;
  wire popcount32_iick_core_132;
  wire popcount32_iick_core_133;
  wire popcount32_iick_core_135;
  wire popcount32_iick_core_136;
  wire popcount32_iick_core_137;
  wire popcount32_iick_core_138;
  wire popcount32_iick_core_139;
  wire popcount32_iick_core_141;
  wire popcount32_iick_core_143;
  wire popcount32_iick_core_144;
  wire popcount32_iick_core_146;
  wire popcount32_iick_core_148;
  wire popcount32_iick_core_150;
  wire popcount32_iick_core_151;
  wire popcount32_iick_core_152;
  wire popcount32_iick_core_153;
  wire popcount32_iick_core_154;
  wire popcount32_iick_core_155;
  wire popcount32_iick_core_156;
  wire popcount32_iick_core_157;
  wire popcount32_iick_core_158;
  wire popcount32_iick_core_159;
  wire popcount32_iick_core_160;
  wire popcount32_iick_core_164;
  wire popcount32_iick_core_165;
  wire popcount32_iick_core_166;
  wire popcount32_iick_core_169;
  wire popcount32_iick_core_170;
  wire popcount32_iick_core_171;
  wire popcount32_iick_core_172;
  wire popcount32_iick_core_174;
  wire popcount32_iick_core_179;
  wire popcount32_iick_core_180;
  wire popcount32_iick_core_184;
  wire popcount32_iick_core_185;
  wire popcount32_iick_core_186;
  wire popcount32_iick_core_187;
  wire popcount32_iick_core_189;
  wire popcount32_iick_core_191;
  wire popcount32_iick_core_193;
  wire popcount32_iick_core_194;
  wire popcount32_iick_core_195;
  wire popcount32_iick_core_196;
  wire popcount32_iick_core_197;
  wire popcount32_iick_core_198;
  wire popcount32_iick_core_203;
  wire popcount32_iick_core_204;
  wire popcount32_iick_core_206;
  wire popcount32_iick_core_207;
  wire popcount32_iick_core_209;
  wire popcount32_iick_core_211;
  wire popcount32_iick_core_212;
  wire popcount32_iick_core_213;
  wire popcount32_iick_core_214;
  wire popcount32_iick_core_215;
  wire popcount32_iick_core_216;
  wire popcount32_iick_core_217;
  wire popcount32_iick_core_218;
  wire popcount32_iick_core_219;
  wire popcount32_iick_core_220;
  wire popcount32_iick_core_221;
  wire popcount32_iick_core_222;
  wire popcount32_iick_core_223;
  wire popcount32_iick_core_225;

  assign popcount32_iick_core_035 = input_a[29] & input_a[19];
  assign popcount32_iick_core_036 = input_a[0] | input_a[19];
  assign popcount32_iick_core_038 = input_a[9] ^ input_a[31];
  assign popcount32_iick_core_040 = popcount32_iick_core_035 | input_a[2];
  assign popcount32_iick_core_041 = ~(input_a[23] ^ input_a[7]);
  assign popcount32_iick_core_042 = popcount32_iick_core_040 | input_a[0];
  assign popcount32_iick_core_043 = ~(input_a[9] ^ input_a[22]);
  assign popcount32_iick_core_045 = input_a[4] ^ input_a[6];
  assign popcount32_iick_core_046 = input_a[4] & input_a[5];
  assign popcount32_iick_core_049 = input_a[13] ^ input_a[3];
  assign popcount32_iick_core_051 = input_a[5] ^ input_a[4];
  assign popcount32_iick_core_052 = popcount32_iick_core_046 & input_a[6];
  assign popcount32_iick_core_053 = popcount32_iick_core_051 | popcount32_iick_core_045;
  assign popcount32_iick_core_056 = ~input_a[19];
  assign popcount32_iick_core_058 = popcount32_iick_core_042 ^ popcount32_iick_core_053;
  assign popcount32_iick_core_059 = popcount32_iick_core_042 & popcount32_iick_core_053;
  assign popcount32_iick_core_061 = input_a[14] | input_a[19];
  assign popcount32_iick_core_064 = input_a[26] & input_a[13];
  assign popcount32_iick_core_065 = popcount32_iick_core_052 | popcount32_iick_core_059;
  assign popcount32_iick_core_066 = input_a[14] ^ input_a[0];
  assign popcount32_iick_core_068 = input_a[8] ^ input_a[9];
  assign popcount32_iick_core_069 = input_a[8] & input_a[9];
  assign popcount32_iick_core_070 = ~(input_a[31] | input_a[23]);
  assign popcount32_iick_core_072 = input_a[15] ^ input_a[26];
  assign popcount32_iick_core_074 = popcount32_iick_core_069 ^ input_a[10];
  assign popcount32_iick_core_075 = input_a[9] & input_a[10];
  assign popcount32_iick_core_076 = popcount32_iick_core_074 ^ popcount32_iick_core_068;
  assign popcount32_iick_core_077 = input_a[10] & input_a[8];
  assign popcount32_iick_core_078 = popcount32_iick_core_075 | popcount32_iick_core_077;
  assign popcount32_iick_core_079 = input_a[12] ^ input_a[13];
  assign popcount32_iick_core_080 = input_a[12] & input_a[13];
  assign popcount32_iick_core_081 = ~input_a[10];
  assign popcount32_iick_core_082 = input_a[18] & input_a[15];
  assign popcount32_iick_core_083 = popcount32_iick_core_079 ^ popcount32_iick_core_081;
  assign popcount32_iick_core_084 = popcount32_iick_core_079 & popcount32_iick_core_081;
  assign popcount32_iick_core_085 = popcount32_iick_core_080 ^ popcount32_iick_core_082;
  assign popcount32_iick_core_086 = popcount32_iick_core_080 & popcount32_iick_core_082;
  assign popcount32_iick_core_087 = popcount32_iick_core_085 ^ popcount32_iick_core_084;
  assign popcount32_iick_core_088 = popcount32_iick_core_085 & popcount32_iick_core_084;
  assign popcount32_iick_core_089 = popcount32_iick_core_086 | popcount32_iick_core_088;
  assign popcount32_iick_core_091 = input_a[30] & popcount32_iick_core_083;
  assign popcount32_iick_core_092 = popcount32_iick_core_076 ^ popcount32_iick_core_087;
  assign popcount32_iick_core_093 = popcount32_iick_core_076 & popcount32_iick_core_087;
  assign popcount32_iick_core_094 = popcount32_iick_core_092 ^ popcount32_iick_core_091;
  assign popcount32_iick_core_095 = popcount32_iick_core_092 & popcount32_iick_core_091;
  assign popcount32_iick_core_096 = popcount32_iick_core_093 | popcount32_iick_core_095;
  assign popcount32_iick_core_097 = popcount32_iick_core_078 ^ popcount32_iick_core_089;
  assign popcount32_iick_core_098 = input_a[10] & popcount32_iick_core_089;
  assign popcount32_iick_core_099 = popcount32_iick_core_097 ^ popcount32_iick_core_096;
  assign popcount32_iick_core_100 = popcount32_iick_core_097 & popcount32_iick_core_096;
  assign popcount32_iick_core_101 = popcount32_iick_core_098 | popcount32_iick_core_100;
  assign popcount32_iick_core_103 = input_a[26] & input_a[6];
  assign popcount32_iick_core_104 = popcount32_iick_core_058 ^ popcount32_iick_core_094;
  assign popcount32_iick_core_105 = popcount32_iick_core_058 & popcount32_iick_core_094;
  assign popcount32_iick_core_106 = input_a[7] & input_a[1];
  assign popcount32_iick_core_109 = popcount32_iick_core_065 ^ popcount32_iick_core_099;
  assign popcount32_iick_core_110 = popcount32_iick_core_065 & popcount32_iick_core_099;
  assign popcount32_iick_core_111 = popcount32_iick_core_109 ^ popcount32_iick_core_105;
  assign popcount32_iick_core_112 = popcount32_iick_core_109 & popcount32_iick_core_105;
  assign popcount32_iick_core_113 = popcount32_iick_core_110 | popcount32_iick_core_112;
  assign popcount32_iick_core_115_not = ~input_a[20];
  assign popcount32_iick_core_116 = popcount32_iick_core_101 | popcount32_iick_core_113;
  assign popcount32_iick_core_118 = input_a[26] & input_a[19];
  assign popcount32_iick_core_119 = input_a[26] | input_a[28];
  assign popcount32_iick_core_120 = ~(input_a[16] ^ input_a[25]);
  assign popcount32_iick_core_121 = ~input_a[19];
  assign popcount32_iick_core_122 = input_a[31] & input_a[25];
  assign popcount32_iick_core_123 = ~(input_a[8] & input_a[1]);
  assign popcount32_iick_core_125 = input_a[16] ^ popcount32_iick_core_122;
  assign popcount32_iick_core_126 = input_a[16] & popcount32_iick_core_122;
  assign popcount32_iick_core_127 = popcount32_iick_core_125 | input_a[3];
  assign popcount32_iick_core_130 = ~(input_a[28] & input_a[15]);
  assign popcount32_iick_core_131 = input_a[20] & input_a[21];
  assign popcount32_iick_core_132 = input_a[22] | input_a[23];
  assign popcount32_iick_core_133 = input_a[22] & input_a[23];
  assign popcount32_iick_core_135 = input_a[14] & popcount32_iick_core_132;
  assign popcount32_iick_core_136 = popcount32_iick_core_131 ^ popcount32_iick_core_133;
  assign popcount32_iick_core_137 = popcount32_iick_core_131 & popcount32_iick_core_133;
  assign popcount32_iick_core_138 = popcount32_iick_core_136 | popcount32_iick_core_135;
  assign popcount32_iick_core_139 = ~(input_a[26] & input_a[11]);
  assign popcount32_iick_core_141 = input_a[15] | input_a[12];
  assign popcount32_iick_core_143 = popcount32_iick_core_127 ^ popcount32_iick_core_138;
  assign popcount32_iick_core_144 = popcount32_iick_core_127 & popcount32_iick_core_138;
  assign popcount32_iick_core_146 = input_a[2] & input_a[4];
  assign popcount32_iick_core_148 = popcount32_iick_core_126 | popcount32_iick_core_137;
  assign popcount32_iick_core_150 = popcount32_iick_core_148 | popcount32_iick_core_144;
  assign popcount32_iick_core_151 = input_a[24] ^ input_a[11];
  assign popcount32_iick_core_152 = ~(input_a[25] & input_a[23]);
  assign popcount32_iick_core_153 = input_a[11] | input_a[20];
  assign popcount32_iick_core_154 = input_a[24] & input_a[28];
  assign popcount32_iick_core_155 = ~(input_a[5] | input_a[15]);
  assign popcount32_iick_core_156 = input_a[26] & input_a[27];
  assign popcount32_iick_core_157 = input_a[11] | input_a[17];
  assign popcount32_iick_core_158 = input_a[3] & input_a[15];
  assign popcount32_iick_core_159 = popcount32_iick_core_154 ^ popcount32_iick_core_156;
  assign popcount32_iick_core_160 = popcount32_iick_core_154 & popcount32_iick_core_156;
  assign popcount32_iick_core_164 = ~input_a[1];
  assign popcount32_iick_core_165 = ~(input_a[3] & input_a[20]);
  assign popcount32_iick_core_166 = ~input_a[13];
  assign popcount32_iick_core_169 = ~(input_a[4] ^ input_a[16]);
  assign popcount32_iick_core_170 = input_a[29] ^ input_a[16];
  assign popcount32_iick_core_171 = ~(input_a[5] ^ input_a[5]);
  assign popcount32_iick_core_172 = ~input_a[31];
  assign popcount32_iick_core_174 = ~input_a[25];
  assign popcount32_iick_core_179 = popcount32_iick_core_159 ^ popcount32_iick_core_157;
  assign popcount32_iick_core_180 = popcount32_iick_core_159 & popcount32_iick_core_157;
  assign popcount32_iick_core_184 = popcount32_iick_core_160 | popcount32_iick_core_180;
  assign popcount32_iick_core_185 = input_a[1] & input_a[12];
  assign popcount32_iick_core_186 = input_a[20] | input_a[27];
  assign popcount32_iick_core_187 = input_a[28] | input_a[21];
  assign popcount32_iick_core_189 = popcount32_iick_core_143 ^ popcount32_iick_core_179;
  assign popcount32_iick_core_191 = ~popcount32_iick_core_189;
  assign popcount32_iick_core_193 = popcount32_iick_core_143 | popcount32_iick_core_189;
  assign popcount32_iick_core_194 = popcount32_iick_core_150 ^ popcount32_iick_core_184;
  assign popcount32_iick_core_195 = popcount32_iick_core_150 & popcount32_iick_core_184;
  assign popcount32_iick_core_196 = popcount32_iick_core_194 ^ popcount32_iick_core_193;
  assign popcount32_iick_core_197 = popcount32_iick_core_194 & popcount32_iick_core_193;
  assign popcount32_iick_core_198 = popcount32_iick_core_195 | popcount32_iick_core_197;
  assign popcount32_iick_core_203 = input_a[27] & input_a[5];
  assign popcount32_iick_core_204 = ~(input_a[4] ^ input_a[29]);
  assign popcount32_iick_core_206 = popcount32_iick_core_106 ^ popcount32_iick_core_191;
  assign popcount32_iick_core_207 = popcount32_iick_core_106 & popcount32_iick_core_191;
  assign popcount32_iick_core_209 = input_a[5] ^ input_a[31];
  assign popcount32_iick_core_211 = popcount32_iick_core_111 ^ popcount32_iick_core_196;
  assign popcount32_iick_core_212 = popcount32_iick_core_111 & popcount32_iick_core_196;
  assign popcount32_iick_core_213 = popcount32_iick_core_211 ^ popcount32_iick_core_207;
  assign popcount32_iick_core_214 = popcount32_iick_core_211 & popcount32_iick_core_207;
  assign popcount32_iick_core_215 = popcount32_iick_core_212 | popcount32_iick_core_214;
  assign popcount32_iick_core_216 = popcount32_iick_core_116 ^ popcount32_iick_core_198;
  assign popcount32_iick_core_217 = popcount32_iick_core_116 & popcount32_iick_core_198;
  assign popcount32_iick_core_218 = popcount32_iick_core_216 ^ popcount32_iick_core_215;
  assign popcount32_iick_core_219 = popcount32_iick_core_216 & popcount32_iick_core_215;
  assign popcount32_iick_core_220 = popcount32_iick_core_217 | popcount32_iick_core_219;
  assign popcount32_iick_core_221 = ~input_a[24];
  assign popcount32_iick_core_222 = input_a[23] & input_a[11];
  assign popcount32_iick_core_223 = input_a[27] & input_a[0];
  assign popcount32_iick_core_225 = ~input_a[25];

  assign popcount32_iick_out[0] = popcount32_iick_core_104;
  assign popcount32_iick_out[1] = popcount32_iick_core_206;
  assign popcount32_iick_out[2] = popcount32_iick_core_213;
  assign popcount32_iick_out[3] = popcount32_iick_core_218;
  assign popcount32_iick_out[4] = popcount32_iick_core_220;
  assign popcount32_iick_out[5] = 1'b0;
endmodule