// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.94958
// WCE=29.0
// EP=0.950328%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_pz4x(input [37:0] input_a, output [5:0] popcount38_pz4x_out);
  wire popcount38_pz4x_core_040;
  wire popcount38_pz4x_core_042;
  wire popcount38_pz4x_core_043;
  wire popcount38_pz4x_core_044;
  wire popcount38_pz4x_core_045;
  wire popcount38_pz4x_core_048;
  wire popcount38_pz4x_core_049;
  wire popcount38_pz4x_core_053;
  wire popcount38_pz4x_core_054;
  wire popcount38_pz4x_core_055;
  wire popcount38_pz4x_core_056;
  wire popcount38_pz4x_core_057;
  wire popcount38_pz4x_core_058;
  wire popcount38_pz4x_core_061;
  wire popcount38_pz4x_core_064;
  wire popcount38_pz4x_core_065;
  wire popcount38_pz4x_core_067;
  wire popcount38_pz4x_core_070;
  wire popcount38_pz4x_core_071;
  wire popcount38_pz4x_core_072;
  wire popcount38_pz4x_core_074;
  wire popcount38_pz4x_core_075;
  wire popcount38_pz4x_core_076;
  wire popcount38_pz4x_core_078;
  wire popcount38_pz4x_core_079;
  wire popcount38_pz4x_core_080;
  wire popcount38_pz4x_core_081;
  wire popcount38_pz4x_core_083;
  wire popcount38_pz4x_core_084;
  wire popcount38_pz4x_core_085;
  wire popcount38_pz4x_core_086;
  wire popcount38_pz4x_core_087;
  wire popcount38_pz4x_core_088;
  wire popcount38_pz4x_core_090;
  wire popcount38_pz4x_core_091;
  wire popcount38_pz4x_core_092;
  wire popcount38_pz4x_core_093;
  wire popcount38_pz4x_core_094;
  wire popcount38_pz4x_core_097;
  wire popcount38_pz4x_core_098;
  wire popcount38_pz4x_core_104;
  wire popcount38_pz4x_core_107;
  wire popcount38_pz4x_core_110;
  wire popcount38_pz4x_core_113;
  wire popcount38_pz4x_core_115;
  wire popcount38_pz4x_core_116;
  wire popcount38_pz4x_core_117;
  wire popcount38_pz4x_core_120;
  wire popcount38_pz4x_core_125;
  wire popcount38_pz4x_core_126;
  wire popcount38_pz4x_core_127;
  wire popcount38_pz4x_core_130;
  wire popcount38_pz4x_core_131;
  wire popcount38_pz4x_core_132;
  wire popcount38_pz4x_core_133;
  wire popcount38_pz4x_core_137;
  wire popcount38_pz4x_core_138;
  wire popcount38_pz4x_core_139;
  wire popcount38_pz4x_core_140;
  wire popcount38_pz4x_core_141;
  wire popcount38_pz4x_core_142_not;
  wire popcount38_pz4x_core_143;
  wire popcount38_pz4x_core_145;
  wire popcount38_pz4x_core_146;
  wire popcount38_pz4x_core_149_not;
  wire popcount38_pz4x_core_151;
  wire popcount38_pz4x_core_152_not;
  wire popcount38_pz4x_core_154;
  wire popcount38_pz4x_core_157;
  wire popcount38_pz4x_core_158;
  wire popcount38_pz4x_core_160;
  wire popcount38_pz4x_core_161;
  wire popcount38_pz4x_core_162;
  wire popcount38_pz4x_core_165;
  wire popcount38_pz4x_core_166;
  wire popcount38_pz4x_core_167;
  wire popcount38_pz4x_core_168;
  wire popcount38_pz4x_core_169;
  wire popcount38_pz4x_core_172;
  wire popcount38_pz4x_core_174;
  wire popcount38_pz4x_core_176;
  wire popcount38_pz4x_core_177;
  wire popcount38_pz4x_core_178;
  wire popcount38_pz4x_core_180;
  wire popcount38_pz4x_core_181;
  wire popcount38_pz4x_core_182;
  wire popcount38_pz4x_core_184;
  wire popcount38_pz4x_core_185;
  wire popcount38_pz4x_core_187;
  wire popcount38_pz4x_core_189;
  wire popcount38_pz4x_core_190;
  wire popcount38_pz4x_core_191;
  wire popcount38_pz4x_core_193_not;
  wire popcount38_pz4x_core_195;
  wire popcount38_pz4x_core_196;
  wire popcount38_pz4x_core_197;
  wire popcount38_pz4x_core_198;
  wire popcount38_pz4x_core_199;
  wire popcount38_pz4x_core_200;
  wire popcount38_pz4x_core_201;
  wire popcount38_pz4x_core_202;
  wire popcount38_pz4x_core_203;
  wire popcount38_pz4x_core_204_not;
  wire popcount38_pz4x_core_205;
  wire popcount38_pz4x_core_209;
  wire popcount38_pz4x_core_211;
  wire popcount38_pz4x_core_213;
  wire popcount38_pz4x_core_214;
  wire popcount38_pz4x_core_215;
  wire popcount38_pz4x_core_216;
  wire popcount38_pz4x_core_217;
  wire popcount38_pz4x_core_218;
  wire popcount38_pz4x_core_219;
  wire popcount38_pz4x_core_220;
  wire popcount38_pz4x_core_221_not;
  wire popcount38_pz4x_core_222;
  wire popcount38_pz4x_core_223;
  wire popcount38_pz4x_core_227;
  wire popcount38_pz4x_core_228;
  wire popcount38_pz4x_core_229;
  wire popcount38_pz4x_core_230;
  wire popcount38_pz4x_core_231;
  wire popcount38_pz4x_core_232;
  wire popcount38_pz4x_core_233;
  wire popcount38_pz4x_core_234;
  wire popcount38_pz4x_core_235;
  wire popcount38_pz4x_core_237;
  wire popcount38_pz4x_core_239;
  wire popcount38_pz4x_core_240;
  wire popcount38_pz4x_core_243;
  wire popcount38_pz4x_core_244;
  wire popcount38_pz4x_core_245;
  wire popcount38_pz4x_core_250;
  wire popcount38_pz4x_core_251;
  wire popcount38_pz4x_core_254;
  wire popcount38_pz4x_core_255;
  wire popcount38_pz4x_core_256;
  wire popcount38_pz4x_core_262;
  wire popcount38_pz4x_core_263;
  wire popcount38_pz4x_core_264;
  wire popcount38_pz4x_core_268;
  wire popcount38_pz4x_core_269;
  wire popcount38_pz4x_core_271;
  wire popcount38_pz4x_core_273;
  wire popcount38_pz4x_core_274;
  wire popcount38_pz4x_core_277;
  wire popcount38_pz4x_core_278;
  wire popcount38_pz4x_core_279;
  wire popcount38_pz4x_core_280;
  wire popcount38_pz4x_core_283;
  wire popcount38_pz4x_core_285;
  wire popcount38_pz4x_core_286;
  wire popcount38_pz4x_core_287;
  wire popcount38_pz4x_core_290;
  wire popcount38_pz4x_core_294;
  wire popcount38_pz4x_core_295;
  wire popcount38_pz4x_core_296;

  assign popcount38_pz4x_core_040 = ~(input_a[24] | input_a[13]);
  assign popcount38_pz4x_core_042 = ~(input_a[33] | input_a[5]);
  assign popcount38_pz4x_core_043 = ~(input_a[13] & input_a[2]);
  assign popcount38_pz4x_core_044 = input_a[0] ^ input_a[9];
  assign popcount38_pz4x_core_045 = ~(input_a[23] & input_a[20]);
  assign popcount38_pz4x_core_048 = ~(input_a[10] ^ input_a[16]);
  assign popcount38_pz4x_core_049 = ~(input_a[27] & input_a[23]);
  assign popcount38_pz4x_core_053 = input_a[27] ^ input_a[1];
  assign popcount38_pz4x_core_054 = ~(input_a[17] | input_a[20]);
  assign popcount38_pz4x_core_055 = ~(input_a[32] ^ input_a[32]);
  assign popcount38_pz4x_core_056 = input_a[19] ^ input_a[5];
  assign popcount38_pz4x_core_057 = ~(input_a[3] | input_a[31]);
  assign popcount38_pz4x_core_058 = input_a[8] & input_a[7];
  assign popcount38_pz4x_core_061 = ~input_a[25];
  assign popcount38_pz4x_core_064 = ~input_a[20];
  assign popcount38_pz4x_core_065 = ~input_a[23];
  assign popcount38_pz4x_core_067 = ~(input_a[27] | input_a[7]);
  assign popcount38_pz4x_core_070 = ~(input_a[6] | input_a[29]);
  assign popcount38_pz4x_core_071 = input_a[13] & input_a[33];
  assign popcount38_pz4x_core_072 = ~(input_a[9] ^ input_a[13]);
  assign popcount38_pz4x_core_074 = ~(input_a[14] ^ input_a[29]);
  assign popcount38_pz4x_core_075 = input_a[2] & input_a[16];
  assign popcount38_pz4x_core_076 = input_a[19] & input_a[3];
  assign popcount38_pz4x_core_078 = input_a[37] | input_a[16];
  assign popcount38_pz4x_core_079 = input_a[33] | input_a[33];
  assign popcount38_pz4x_core_080 = ~(input_a[30] & input_a[2]);
  assign popcount38_pz4x_core_081 = input_a[15] | input_a[29];
  assign popcount38_pz4x_core_083 = input_a[23] ^ input_a[7];
  assign popcount38_pz4x_core_084 = ~input_a[2];
  assign popcount38_pz4x_core_085 = ~(input_a[34] ^ input_a[20]);
  assign popcount38_pz4x_core_086 = input_a[2] ^ input_a[6];
  assign popcount38_pz4x_core_087 = ~(input_a[16] & input_a[36]);
  assign popcount38_pz4x_core_088 = input_a[24] ^ input_a[4];
  assign popcount38_pz4x_core_090 = ~(input_a[33] & input_a[23]);
  assign popcount38_pz4x_core_091 = input_a[23] ^ input_a[23];
  assign popcount38_pz4x_core_092 = ~(input_a[16] ^ input_a[35]);
  assign popcount38_pz4x_core_093 = input_a[32] | input_a[30];
  assign popcount38_pz4x_core_094 = ~input_a[21];
  assign popcount38_pz4x_core_097 = ~input_a[25];
  assign popcount38_pz4x_core_098 = ~(input_a[27] | input_a[30]);
  assign popcount38_pz4x_core_104 = ~(input_a[16] ^ input_a[18]);
  assign popcount38_pz4x_core_107 = input_a[28] & input_a[20];
  assign popcount38_pz4x_core_110 = ~(input_a[8] ^ input_a[16]);
  assign popcount38_pz4x_core_113 = ~(input_a[12] & input_a[20]);
  assign popcount38_pz4x_core_115 = input_a[5] | input_a[16];
  assign popcount38_pz4x_core_116 = input_a[25] ^ input_a[8];
  assign popcount38_pz4x_core_117 = input_a[23] & input_a[10];
  assign popcount38_pz4x_core_120 = ~(input_a[0] ^ input_a[5]);
  assign popcount38_pz4x_core_125 = ~(input_a[7] ^ input_a[32]);
  assign popcount38_pz4x_core_126 = input_a[34] & input_a[8];
  assign popcount38_pz4x_core_127 = ~input_a[10];
  assign popcount38_pz4x_core_130 = input_a[5] & input_a[8];
  assign popcount38_pz4x_core_131 = ~(input_a[28] | input_a[26]);
  assign popcount38_pz4x_core_132 = input_a[7] & input_a[36];
  assign popcount38_pz4x_core_133 = input_a[19] ^ input_a[1];
  assign popcount38_pz4x_core_137 = ~(input_a[7] ^ input_a[23]);
  assign popcount38_pz4x_core_138 = ~(input_a[10] ^ input_a[17]);
  assign popcount38_pz4x_core_139 = ~(input_a[27] | input_a[23]);
  assign popcount38_pz4x_core_140 = input_a[33] ^ input_a[8];
  assign popcount38_pz4x_core_141 = ~(input_a[28] & input_a[17]);
  assign popcount38_pz4x_core_142_not = ~input_a[34];
  assign popcount38_pz4x_core_143 = input_a[21] | input_a[22];
  assign popcount38_pz4x_core_145 = input_a[28] & input_a[15];
  assign popcount38_pz4x_core_146 = input_a[2] & input_a[33];
  assign popcount38_pz4x_core_149_not = ~input_a[6];
  assign popcount38_pz4x_core_151 = ~(input_a[24] | input_a[34]);
  assign popcount38_pz4x_core_152_not = ~input_a[3];
  assign popcount38_pz4x_core_154 = ~(input_a[11] | input_a[21]);
  assign popcount38_pz4x_core_157 = ~(input_a[0] | input_a[8]);
  assign popcount38_pz4x_core_158 = input_a[14] & input_a[36];
  assign popcount38_pz4x_core_160 = ~(input_a[31] | input_a[1]);
  assign popcount38_pz4x_core_161 = ~(input_a[9] ^ input_a[4]);
  assign popcount38_pz4x_core_162 = ~input_a[15];
  assign popcount38_pz4x_core_165 = ~input_a[22];
  assign popcount38_pz4x_core_166 = ~input_a[9];
  assign popcount38_pz4x_core_167 = input_a[18] ^ input_a[3];
  assign popcount38_pz4x_core_168 = ~input_a[13];
  assign popcount38_pz4x_core_169 = ~input_a[20];
  assign popcount38_pz4x_core_172 = ~input_a[27];
  assign popcount38_pz4x_core_174 = ~(input_a[1] ^ input_a[13]);
  assign popcount38_pz4x_core_176 = ~input_a[25];
  assign popcount38_pz4x_core_177 = input_a[22] ^ input_a[22];
  assign popcount38_pz4x_core_178 = input_a[6] & input_a[22];
  assign popcount38_pz4x_core_180 = ~input_a[31];
  assign popcount38_pz4x_core_181 = ~(input_a[35] | input_a[13]);
  assign popcount38_pz4x_core_182 = input_a[14] | input_a[24];
  assign popcount38_pz4x_core_184 = ~(input_a[17] & input_a[25]);
  assign popcount38_pz4x_core_185 = ~(input_a[25] ^ input_a[13]);
  assign popcount38_pz4x_core_187 = ~(input_a[22] & input_a[25]);
  assign popcount38_pz4x_core_189 = input_a[16] ^ input_a[28];
  assign popcount38_pz4x_core_190 = input_a[30] | input_a[8];
  assign popcount38_pz4x_core_191 = ~(input_a[10] & input_a[35]);
  assign popcount38_pz4x_core_193_not = ~input_a[20];
  assign popcount38_pz4x_core_195 = input_a[27] & input_a[20];
  assign popcount38_pz4x_core_196 = input_a[4] | input_a[15];
  assign popcount38_pz4x_core_197 = ~(input_a[0] | input_a[22]);
  assign popcount38_pz4x_core_198 = ~(input_a[12] | input_a[14]);
  assign popcount38_pz4x_core_199 = ~(input_a[8] | input_a[4]);
  assign popcount38_pz4x_core_200 = input_a[7] ^ input_a[19];
  assign popcount38_pz4x_core_201 = input_a[21] ^ input_a[14];
  assign popcount38_pz4x_core_202 = ~(input_a[24] | input_a[1]);
  assign popcount38_pz4x_core_203 = ~(input_a[3] | input_a[2]);
  assign popcount38_pz4x_core_204_not = ~input_a[18];
  assign popcount38_pz4x_core_205 = input_a[31] ^ input_a[13];
  assign popcount38_pz4x_core_209 = ~(input_a[10] ^ input_a[31]);
  assign popcount38_pz4x_core_211 = ~(input_a[23] | input_a[18]);
  assign popcount38_pz4x_core_213 = ~(input_a[34] & input_a[14]);
  assign popcount38_pz4x_core_214 = input_a[7] ^ input_a[14];
  assign popcount38_pz4x_core_215 = ~(input_a[7] ^ input_a[6]);
  assign popcount38_pz4x_core_216 = ~(input_a[12] ^ input_a[9]);
  assign popcount38_pz4x_core_217 = input_a[1] | input_a[32];
  assign popcount38_pz4x_core_218 = ~(input_a[12] & input_a[19]);
  assign popcount38_pz4x_core_219 = ~(input_a[15] | input_a[33]);
  assign popcount38_pz4x_core_220 = ~input_a[37];
  assign popcount38_pz4x_core_221_not = ~input_a[14];
  assign popcount38_pz4x_core_222 = ~(input_a[32] | input_a[14]);
  assign popcount38_pz4x_core_223 = input_a[9] & input_a[10];
  assign popcount38_pz4x_core_227 = input_a[37] & input_a[27];
  assign popcount38_pz4x_core_228 = input_a[1] ^ input_a[21];
  assign popcount38_pz4x_core_229 = ~input_a[15];
  assign popcount38_pz4x_core_230 = ~(input_a[18] & input_a[1]);
  assign popcount38_pz4x_core_231 = input_a[32] ^ input_a[15];
  assign popcount38_pz4x_core_232 = input_a[16] | input_a[20];
  assign popcount38_pz4x_core_233 = input_a[19] | input_a[19];
  assign popcount38_pz4x_core_234 = input_a[22] & input_a[28];
  assign popcount38_pz4x_core_235 = input_a[19] ^ input_a[16];
  assign popcount38_pz4x_core_237 = input_a[31] ^ input_a[24];
  assign popcount38_pz4x_core_239 = ~(input_a[27] ^ input_a[30]);
  assign popcount38_pz4x_core_240 = input_a[4] & input_a[30];
  assign popcount38_pz4x_core_243 = ~(input_a[36] & input_a[12]);
  assign popcount38_pz4x_core_244 = input_a[6] & input_a[19];
  assign popcount38_pz4x_core_245 = ~(input_a[33] ^ input_a[2]);
  assign popcount38_pz4x_core_250 = input_a[5] | input_a[21];
  assign popcount38_pz4x_core_251 = ~(input_a[12] ^ input_a[36]);
  assign popcount38_pz4x_core_254 = input_a[33] ^ input_a[36];
  assign popcount38_pz4x_core_255 = input_a[8] | input_a[17];
  assign popcount38_pz4x_core_256 = ~(input_a[15] ^ input_a[15]);
  assign popcount38_pz4x_core_262 = input_a[31] & input_a[14];
  assign popcount38_pz4x_core_263 = input_a[3] | input_a[0];
  assign popcount38_pz4x_core_264 = ~(input_a[16] ^ input_a[27]);
  assign popcount38_pz4x_core_268 = ~(input_a[12] | input_a[22]);
  assign popcount38_pz4x_core_269 = ~(input_a[12] ^ input_a[10]);
  assign popcount38_pz4x_core_271 = input_a[34] & input_a[10];
  assign popcount38_pz4x_core_273 = input_a[13] & input_a[3];
  assign popcount38_pz4x_core_274 = input_a[19] & input_a[29];
  assign popcount38_pz4x_core_277 = input_a[24] | input_a[1];
  assign popcount38_pz4x_core_278 = ~(input_a[32] ^ input_a[4]);
  assign popcount38_pz4x_core_279 = ~(input_a[12] & input_a[33]);
  assign popcount38_pz4x_core_280 = ~input_a[2];
  assign popcount38_pz4x_core_283 = ~input_a[21];
  assign popcount38_pz4x_core_285 = ~(input_a[4] | input_a[26]);
  assign popcount38_pz4x_core_286 = ~(input_a[12] | input_a[31]);
  assign popcount38_pz4x_core_287 = ~(input_a[15] | input_a[11]);
  assign popcount38_pz4x_core_290 = ~(input_a[10] | input_a[9]);
  assign popcount38_pz4x_core_294 = ~(input_a[2] & input_a[16]);
  assign popcount38_pz4x_core_295 = input_a[15] & input_a[6];
  assign popcount38_pz4x_core_296 = input_a[32] | input_a[23];

  assign popcount38_pz4x_out[0] = 1'b1;
  assign popcount38_pz4x_out[1] = input_a[32];
  assign popcount38_pz4x_out[2] = input_a[32];
  assign popcount38_pz4x_out[3] = input_a[15];
  assign popcount38_pz4x_out[4] = 1'b1;
  assign popcount38_pz4x_out[5] = 1'b0;
endmodule