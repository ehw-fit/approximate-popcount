// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.42922
// WCE=20.0
// EP=0.943987%
// Printed PDK parameters:
//  Area=12118344.0
//  Delay=28491136.0
//  Power=485560.0

module popcount40_kz6j(input [39:0] input_a, output [5:0] popcount40_kz6j_out);
  wire popcount40_kz6j_core_042;
  wire popcount40_kz6j_core_043;
  wire popcount40_kz6j_core_044;
  wire popcount40_kz6j_core_045;
  wire popcount40_kz6j_core_046;
  wire popcount40_kz6j_core_047;
  wire popcount40_kz6j_core_048;
  wire popcount40_kz6j_core_051;
  wire popcount40_kz6j_core_052;
  wire popcount40_kz6j_core_053;
  wire popcount40_kz6j_core_054;
  wire popcount40_kz6j_core_055;
  wire popcount40_kz6j_core_058;
  wire popcount40_kz6j_core_059;
  wire popcount40_kz6j_core_061;
  wire popcount40_kz6j_core_062;
  wire popcount40_kz6j_core_063;
  wire popcount40_kz6j_core_064;
  wire popcount40_kz6j_core_067;
  wire popcount40_kz6j_core_068;
  wire popcount40_kz6j_core_070;
  wire popcount40_kz6j_core_075;
  wire popcount40_kz6j_core_076;
  wire popcount40_kz6j_core_079;
  wire popcount40_kz6j_core_080;
  wire popcount40_kz6j_core_081;
  wire popcount40_kz6j_core_083;
  wire popcount40_kz6j_core_084;
  wire popcount40_kz6j_core_085;
  wire popcount40_kz6j_core_086;
  wire popcount40_kz6j_core_087;
  wire popcount40_kz6j_core_089;
  wire popcount40_kz6j_core_091;
  wire popcount40_kz6j_core_093;
  wire popcount40_kz6j_core_094;
  wire popcount40_kz6j_core_095;
  wire popcount40_kz6j_core_097;
  wire popcount40_kz6j_core_100_not;
  wire popcount40_kz6j_core_101;
  wire popcount40_kz6j_core_102;
  wire popcount40_kz6j_core_105;
  wire popcount40_kz6j_core_107;
  wire popcount40_kz6j_core_109;
  wire popcount40_kz6j_core_112;
  wire popcount40_kz6j_core_115;
  wire popcount40_kz6j_core_116;
  wire popcount40_kz6j_core_119;
  wire popcount40_kz6j_core_120;
  wire popcount40_kz6j_core_121_not;
  wire popcount40_kz6j_core_122;
  wire popcount40_kz6j_core_125;
  wire popcount40_kz6j_core_128;
  wire popcount40_kz6j_core_130;
  wire popcount40_kz6j_core_133;
  wire popcount40_kz6j_core_134;
  wire popcount40_kz6j_core_135;
  wire popcount40_kz6j_core_137;
  wire popcount40_kz6j_core_138;
  wire popcount40_kz6j_core_141;
  wire popcount40_kz6j_core_143;
  wire popcount40_kz6j_core_145;
  wire popcount40_kz6j_core_146;
  wire popcount40_kz6j_core_147;
  wire popcount40_kz6j_core_148;
  wire popcount40_kz6j_core_151;
  wire popcount40_kz6j_core_152;
  wire popcount40_kz6j_core_153;
  wire popcount40_kz6j_core_154;
  wire popcount40_kz6j_core_155;
  wire popcount40_kz6j_core_158;
  wire popcount40_kz6j_core_162;
  wire popcount40_kz6j_core_166;
  wire popcount40_kz6j_core_168;
  wire popcount40_kz6j_core_169;
  wire popcount40_kz6j_core_171;
  wire popcount40_kz6j_core_173;
  wire popcount40_kz6j_core_175;
  wire popcount40_kz6j_core_176;
  wire popcount40_kz6j_core_178;
  wire popcount40_kz6j_core_180;
  wire popcount40_kz6j_core_181;
  wire popcount40_kz6j_core_183;
  wire popcount40_kz6j_core_184;
  wire popcount40_kz6j_core_185;
  wire popcount40_kz6j_core_187;
  wire popcount40_kz6j_core_188;
  wire popcount40_kz6j_core_189;
  wire popcount40_kz6j_core_190;
  wire popcount40_kz6j_core_192;
  wire popcount40_kz6j_core_193;
  wire popcount40_kz6j_core_197;
  wire popcount40_kz6j_core_199;
  wire popcount40_kz6j_core_201;
  wire popcount40_kz6j_core_203;
  wire popcount40_kz6j_core_204;
  wire popcount40_kz6j_core_207;
  wire popcount40_kz6j_core_208;
  wire popcount40_kz6j_core_209;
  wire popcount40_kz6j_core_210;
  wire popcount40_kz6j_core_211;
  wire popcount40_kz6j_core_215;
  wire popcount40_kz6j_core_216;
  wire popcount40_kz6j_core_217;
  wire popcount40_kz6j_core_219;
  wire popcount40_kz6j_core_220;
  wire popcount40_kz6j_core_221;
  wire popcount40_kz6j_core_222;
  wire popcount40_kz6j_core_223;
  wire popcount40_kz6j_core_224;
  wire popcount40_kz6j_core_225;
  wire popcount40_kz6j_core_226;
  wire popcount40_kz6j_core_228;
  wire popcount40_kz6j_core_229;
  wire popcount40_kz6j_core_233;
  wire popcount40_kz6j_core_235;
  wire popcount40_kz6j_core_236;
  wire popcount40_kz6j_core_238;
  wire popcount40_kz6j_core_240_not;
  wire popcount40_kz6j_core_243;
  wire popcount40_kz6j_core_244;
  wire popcount40_kz6j_core_245;
  wire popcount40_kz6j_core_246;
  wire popcount40_kz6j_core_247;
  wire popcount40_kz6j_core_248;
  wire popcount40_kz6j_core_252;
  wire popcount40_kz6j_core_254;
  wire popcount40_kz6j_core_255;
  wire popcount40_kz6j_core_256;
  wire popcount40_kz6j_core_257;
  wire popcount40_kz6j_core_261;
  wire popcount40_kz6j_core_262;
  wire popcount40_kz6j_core_263;
  wire popcount40_kz6j_core_265;
  wire popcount40_kz6j_core_266;
  wire popcount40_kz6j_core_267;
  wire popcount40_kz6j_core_268;
  wire popcount40_kz6j_core_269;
  wire popcount40_kz6j_core_270;
  wire popcount40_kz6j_core_271;
  wire popcount40_kz6j_core_272;
  wire popcount40_kz6j_core_273;
  wire popcount40_kz6j_core_274;
  wire popcount40_kz6j_core_275;
  wire popcount40_kz6j_core_276;
  wire popcount40_kz6j_core_281;
  wire popcount40_kz6j_core_284;
  wire popcount40_kz6j_core_288;
  wire popcount40_kz6j_core_290;
  wire popcount40_kz6j_core_291;
  wire popcount40_kz6j_core_293;
  wire popcount40_kz6j_core_294;
  wire popcount40_kz6j_core_295;
  wire popcount40_kz6j_core_299;
  wire popcount40_kz6j_core_300;
  wire popcount40_kz6j_core_302;
  wire popcount40_kz6j_core_303;
  wire popcount40_kz6j_core_304;
  wire popcount40_kz6j_core_305;
  wire popcount40_kz6j_core_306;
  wire popcount40_kz6j_core_308;
  wire popcount40_kz6j_core_309;
  wire popcount40_kz6j_core_310;
  wire popcount40_kz6j_core_311;
  wire popcount40_kz6j_core_312;
  wire popcount40_kz6j_core_314;
  wire popcount40_kz6j_core_315;
  wire popcount40_kz6j_core_316;

  assign popcount40_kz6j_core_042 = ~(input_a[18] & input_a[25]);
  assign popcount40_kz6j_core_043 = input_a[4] & input_a[18];
  assign popcount40_kz6j_core_044 = input_a[7] ^ input_a[9];
  assign popcount40_kz6j_core_045 = ~(input_a[28] | input_a[13]);
  assign popcount40_kz6j_core_046 = input_a[16] | input_a[16];
  assign popcount40_kz6j_core_047 = ~(input_a[28] | input_a[7]);
  assign popcount40_kz6j_core_048 = ~(input_a[12] ^ input_a[2]);
  assign popcount40_kz6j_core_051 = ~(input_a[4] ^ input_a[23]);
  assign popcount40_kz6j_core_052 = input_a[7] & input_a[27];
  assign popcount40_kz6j_core_053 = popcount40_kz6j_core_043 & input_a[14];
  assign popcount40_kz6j_core_054 = input_a[36] | input_a[18];
  assign popcount40_kz6j_core_055 = ~(input_a[36] ^ input_a[21]);
  assign popcount40_kz6j_core_058 = ~(input_a[31] ^ input_a[19]);
  assign popcount40_kz6j_core_059 = ~(input_a[21] ^ input_a[3]);
  assign popcount40_kz6j_core_061 = input_a[33] ^ input_a[18];
  assign popcount40_kz6j_core_062 = input_a[24] & input_a[27];
  assign popcount40_kz6j_core_063 = input_a[7] | input_a[14];
  assign popcount40_kz6j_core_064 = input_a[17] | input_a[0];
  assign popcount40_kz6j_core_067 = input_a[33] ^ input_a[23];
  assign popcount40_kz6j_core_068 = input_a[1] & input_a[23];
  assign popcount40_kz6j_core_070 = input_a[10] & popcount40_kz6j_core_062;
  assign popcount40_kz6j_core_075 = input_a[21] ^ input_a[28];
  assign popcount40_kz6j_core_076 = ~(input_a[24] & input_a[13]);
  assign popcount40_kz6j_core_079 = input_a[38] & popcount40_kz6j_core_068;
  assign popcount40_kz6j_core_080 = ~input_a[5];
  assign popcount40_kz6j_core_081 = ~input_a[17];
  assign popcount40_kz6j_core_083 = popcount40_kz6j_core_053 | popcount40_kz6j_core_070;
  assign popcount40_kz6j_core_084 = popcount40_kz6j_core_053 & popcount40_kz6j_core_070;
  assign popcount40_kz6j_core_085 = popcount40_kz6j_core_083 | popcount40_kz6j_core_079;
  assign popcount40_kz6j_core_086 = popcount40_kz6j_core_083 & popcount40_kz6j_core_079;
  assign popcount40_kz6j_core_087 = popcount40_kz6j_core_084 | popcount40_kz6j_core_086;
  assign popcount40_kz6j_core_089 = ~input_a[30];
  assign popcount40_kz6j_core_091 = input_a[23] ^ input_a[39];
  assign popcount40_kz6j_core_093 = input_a[4] ^ input_a[19];
  assign popcount40_kz6j_core_094 = ~(input_a[33] | input_a[0]);
  assign popcount40_kz6j_core_095 = input_a[17] ^ input_a[5];
  assign popcount40_kz6j_core_097 = input_a[35] | input_a[12];
  assign popcount40_kz6j_core_100_not = ~input_a[2];
  assign popcount40_kz6j_core_101 = ~(input_a[1] | input_a[2]);
  assign popcount40_kz6j_core_102 = ~(input_a[16] | input_a[12]);
  assign popcount40_kz6j_core_105 = input_a[37] & input_a[17];
  assign popcount40_kz6j_core_107 = ~(input_a[20] | input_a[15]);
  assign popcount40_kz6j_core_109 = input_a[11] | input_a[2];
  assign popcount40_kz6j_core_112 = ~input_a[25];
  assign popcount40_kz6j_core_115 = ~(input_a[1] & input_a[7]);
  assign popcount40_kz6j_core_116 = ~(input_a[15] ^ input_a[17]);
  assign popcount40_kz6j_core_119 = ~input_a[14];
  assign popcount40_kz6j_core_120 = ~(input_a[37] & input_a[28]);
  assign popcount40_kz6j_core_121_not = ~input_a[31];
  assign popcount40_kz6j_core_122 = ~input_a[5];
  assign popcount40_kz6j_core_125 = ~(input_a[24] ^ input_a[4]);
  assign popcount40_kz6j_core_128 = ~(input_a[34] ^ input_a[24]);
  assign popcount40_kz6j_core_130 = input_a[7] & input_a[4];
  assign popcount40_kz6j_core_133 = ~(input_a[35] ^ input_a[38]);
  assign popcount40_kz6j_core_134 = input_a[39] & input_a[14];
  assign popcount40_kz6j_core_135 = input_a[23] ^ input_a[29];
  assign popcount40_kz6j_core_137 = input_a[0] ^ input_a[21];
  assign popcount40_kz6j_core_138 = ~(input_a[30] | input_a[13]);
  assign popcount40_kz6j_core_141 = input_a[32] ^ input_a[21];
  assign popcount40_kz6j_core_143 = input_a[34] & input_a[6];
  assign popcount40_kz6j_core_145 = input_a[27] | input_a[23];
  assign popcount40_kz6j_core_146 = ~(input_a[36] | input_a[23]);
  assign popcount40_kz6j_core_147 = input_a[23] & input_a[7];
  assign popcount40_kz6j_core_148 = ~(input_a[26] | input_a[6]);
  assign popcount40_kz6j_core_151 = ~popcount40_kz6j_core_085;
  assign popcount40_kz6j_core_152 = input_a[16] ^ input_a[21];
  assign popcount40_kz6j_core_153 = ~popcount40_kz6j_core_151;
  assign popcount40_kz6j_core_154 = ~input_a[35];
  assign popcount40_kz6j_core_155 = input_a[8] ^ input_a[29];
  assign popcount40_kz6j_core_158 = ~popcount40_kz6j_core_087;
  assign popcount40_kz6j_core_162 = ~(input_a[24] ^ input_a[20]);
  assign popcount40_kz6j_core_166 = input_a[0] & input_a[38];
  assign popcount40_kz6j_core_168 = ~input_a[29];
  assign popcount40_kz6j_core_169 = input_a[27] | input_a[11];
  assign popcount40_kz6j_core_171 = ~(input_a[37] ^ input_a[0]);
  assign popcount40_kz6j_core_173 = input_a[11] ^ input_a[12];
  assign popcount40_kz6j_core_175 = ~(input_a[3] & input_a[4]);
  assign popcount40_kz6j_core_176 = ~input_a[8];
  assign popcount40_kz6j_core_178 = ~(input_a[36] | input_a[22]);
  assign popcount40_kz6j_core_180 = ~(input_a[30] ^ input_a[33]);
  assign popcount40_kz6j_core_181 = ~(input_a[9] | input_a[39]);
  assign popcount40_kz6j_core_183 = ~(input_a[32] | input_a[31]);
  assign popcount40_kz6j_core_184 = ~(input_a[28] & input_a[12]);
  assign popcount40_kz6j_core_185 = ~input_a[14];
  assign popcount40_kz6j_core_187 = ~(input_a[0] & input_a[25]);
  assign popcount40_kz6j_core_188 = ~(input_a[25] | input_a[7]);
  assign popcount40_kz6j_core_189 = ~(input_a[13] ^ input_a[21]);
  assign popcount40_kz6j_core_190 = input_a[21] & input_a[0];
  assign popcount40_kz6j_core_192 = ~(input_a[19] & input_a[21]);
  assign popcount40_kz6j_core_193 = ~(input_a[18] & input_a[25]);
  assign popcount40_kz6j_core_197 = input_a[39] | input_a[24];
  assign popcount40_kz6j_core_199 = input_a[26] | input_a[15];
  assign popcount40_kz6j_core_201 = input_a[5] | input_a[23];
  assign popcount40_kz6j_core_203 = input_a[27] & input_a[28];
  assign popcount40_kz6j_core_204 = input_a[30] & input_a[35];
  assign popcount40_kz6j_core_207 = input_a[9] | input_a[17];
  assign popcount40_kz6j_core_208 = ~(input_a[29] | input_a[6]);
  assign popcount40_kz6j_core_209 = input_a[34] | input_a[19];
  assign popcount40_kz6j_core_210 = ~input_a[18];
  assign popcount40_kz6j_core_211 = ~input_a[24];
  assign popcount40_kz6j_core_215 = ~(input_a[23] | input_a[7]);
  assign popcount40_kz6j_core_216 = input_a[0] | input_a[8];
  assign popcount40_kz6j_core_217 = input_a[2] | input_a[24];
  assign popcount40_kz6j_core_219 = input_a[15] ^ input_a[28];
  assign popcount40_kz6j_core_220 = input_a[11] & input_a[38];
  assign popcount40_kz6j_core_221 = ~(input_a[21] ^ input_a[5]);
  assign popcount40_kz6j_core_222 = ~(input_a[20] | input_a[5]);
  assign popcount40_kz6j_core_223 = input_a[20] ^ input_a[19];
  assign popcount40_kz6j_core_224 = ~(input_a[21] & input_a[31]);
  assign popcount40_kz6j_core_225 = input_a[11] | input_a[27];
  assign popcount40_kz6j_core_226 = input_a[22] ^ input_a[28];
  assign popcount40_kz6j_core_228 = ~(input_a[19] | input_a[18]);
  assign popcount40_kz6j_core_229 = input_a[31] ^ input_a[27];
  assign popcount40_kz6j_core_233 = ~(input_a[35] ^ input_a[28]);
  assign popcount40_kz6j_core_235 = input_a[3] & input_a[11];
  assign popcount40_kz6j_core_236 = ~(input_a[1] ^ input_a[3]);
  assign popcount40_kz6j_core_238 = input_a[18] ^ input_a[23];
  assign popcount40_kz6j_core_240_not = ~input_a[29];
  assign popcount40_kz6j_core_243 = input_a[16] & input_a[33];
  assign popcount40_kz6j_core_244 = input_a[30] & input_a[2];
  assign popcount40_kz6j_core_245 = popcount40_kz6j_core_235 & input_a[12];
  assign popcount40_kz6j_core_246 = ~(input_a[26] ^ input_a[31]);
  assign popcount40_kz6j_core_247 = input_a[29] & popcount40_kz6j_core_243;
  assign popcount40_kz6j_core_248 = popcount40_kz6j_core_245 | popcount40_kz6j_core_247;
  assign popcount40_kz6j_core_252 = ~(input_a[12] & input_a[36]);
  assign popcount40_kz6j_core_254 = ~input_a[36];
  assign popcount40_kz6j_core_255 = input_a[1] & input_a[31];
  assign popcount40_kz6j_core_256 = input_a[6] & input_a[8];
  assign popcount40_kz6j_core_257 = input_a[7] ^ input_a[12];
  assign popcount40_kz6j_core_261 = input_a[32] ^ input_a[27];
  assign popcount40_kz6j_core_262 = ~(input_a[0] ^ input_a[11]);
  assign popcount40_kz6j_core_263 = ~(input_a[32] ^ input_a[23]);
  assign popcount40_kz6j_core_265 = ~(input_a[16] | input_a[21]);
  assign popcount40_kz6j_core_266 = ~input_a[0];
  assign popcount40_kz6j_core_267 = ~input_a[15];
  assign popcount40_kz6j_core_268 = input_a[38] | input_a[21];
  assign popcount40_kz6j_core_269 = ~(input_a[8] & input_a[4]);
  assign popcount40_kz6j_core_270 = ~(input_a[2] & input_a[9]);
  assign popcount40_kz6j_core_271 = input_a[13] & input_a[17];
  assign popcount40_kz6j_core_272 = input_a[2] & input_a[35];
  assign popcount40_kz6j_core_273 = ~(input_a[0] ^ input_a[3]);
  assign popcount40_kz6j_core_274 = input_a[25] & input_a[35];
  assign popcount40_kz6j_core_275 = ~(input_a[34] | input_a[5]);
  assign popcount40_kz6j_core_276 = popcount40_kz6j_core_209 & popcount40_kz6j_core_248;
  assign popcount40_kz6j_core_281 = input_a[4] ^ input_a[33];
  assign popcount40_kz6j_core_284 = ~(input_a[12] & input_a[31]);
  assign popcount40_kz6j_core_288 = input_a[16] ^ input_a[1];
  assign popcount40_kz6j_core_290 = input_a[15] | input_a[6];
  assign popcount40_kz6j_core_291 = input_a[26] & input_a[13];
  assign popcount40_kz6j_core_293 = input_a[17] & popcount40_kz6j_core_272;
  assign popcount40_kz6j_core_294 = input_a[22] | input_a[21];
  assign popcount40_kz6j_core_295 = input_a[12] & input_a[15];
  assign popcount40_kz6j_core_299 = ~(input_a[31] | input_a[6]);
  assign popcount40_kz6j_core_300 = popcount40_kz6j_core_153 & popcount40_kz6j_core_293;
  assign popcount40_kz6j_core_302 = popcount40_kz6j_core_158 ^ popcount40_kz6j_core_276;
  assign popcount40_kz6j_core_303 = popcount40_kz6j_core_158 & popcount40_kz6j_core_276;
  assign popcount40_kz6j_core_304 = popcount40_kz6j_core_302 ^ popcount40_kz6j_core_300;
  assign popcount40_kz6j_core_305 = input_a[2] & popcount40_kz6j_core_300;
  assign popcount40_kz6j_core_306 = popcount40_kz6j_core_303 | popcount40_kz6j_core_305;
  assign popcount40_kz6j_core_308 = input_a[9] & input_a[7];
  assign popcount40_kz6j_core_309 = popcount40_kz6j_core_087 | popcount40_kz6j_core_306;
  assign popcount40_kz6j_core_310 = ~(input_a[3] | input_a[15]);
  assign popcount40_kz6j_core_311 = input_a[4] ^ input_a[9];
  assign popcount40_kz6j_core_312 = ~(input_a[21] & input_a[39]);
  assign popcount40_kz6j_core_314 = input_a[18] | input_a[2];
  assign popcount40_kz6j_core_315 = input_a[20] & input_a[37];
  assign popcount40_kz6j_core_316 = input_a[0] | input_a[17];

  assign popcount40_kz6j_out[0] = input_a[8];
  assign popcount40_kz6j_out[1] = popcount40_kz6j_core_158;
  assign popcount40_kz6j_out[2] = 1'b1;
  assign popcount40_kz6j_out[3] = popcount40_kz6j_core_304;
  assign popcount40_kz6j_out[4] = popcount40_kz6j_core_309;
  assign popcount40_kz6j_out[5] = 1'b0;
endmodule