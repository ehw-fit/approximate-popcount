// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5001
// WCE=38.0
// EP=0.999876%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_vg2l(input [34:0] input_a, output [5:0] popcount35_vg2l_out);
  wire popcount35_vg2l_core_037;
  wire popcount35_vg2l_core_038;
  wire popcount35_vg2l_core_041;
  wire popcount35_vg2l_core_042;
  wire popcount35_vg2l_core_044;
  wire popcount35_vg2l_core_046;
  wire popcount35_vg2l_core_047;
  wire popcount35_vg2l_core_048_not;
  wire popcount35_vg2l_core_049;
  wire popcount35_vg2l_core_050;
  wire popcount35_vg2l_core_051;
  wire popcount35_vg2l_core_052;
  wire popcount35_vg2l_core_054;
  wire popcount35_vg2l_core_055;
  wire popcount35_vg2l_core_056;
  wire popcount35_vg2l_core_057;
  wire popcount35_vg2l_core_058;
  wire popcount35_vg2l_core_060;
  wire popcount35_vg2l_core_061;
  wire popcount35_vg2l_core_062;
  wire popcount35_vg2l_core_065;
  wire popcount35_vg2l_core_067;
  wire popcount35_vg2l_core_068;
  wire popcount35_vg2l_core_069;
  wire popcount35_vg2l_core_071;
  wire popcount35_vg2l_core_072;
  wire popcount35_vg2l_core_073;
  wire popcount35_vg2l_core_075_not;
  wire popcount35_vg2l_core_076;
  wire popcount35_vg2l_core_077;
  wire popcount35_vg2l_core_079;
  wire popcount35_vg2l_core_080;
  wire popcount35_vg2l_core_081;
  wire popcount35_vg2l_core_083;
  wire popcount35_vg2l_core_084;
  wire popcount35_vg2l_core_085;
  wire popcount35_vg2l_core_088;
  wire popcount35_vg2l_core_089;
  wire popcount35_vg2l_core_090;
  wire popcount35_vg2l_core_093;
  wire popcount35_vg2l_core_097;
  wire popcount35_vg2l_core_098;
  wire popcount35_vg2l_core_100;
  wire popcount35_vg2l_core_103;
  wire popcount35_vg2l_core_104;
  wire popcount35_vg2l_core_105;
  wire popcount35_vg2l_core_107;
  wire popcount35_vg2l_core_108;
  wire popcount35_vg2l_core_109;
  wire popcount35_vg2l_core_112;
  wire popcount35_vg2l_core_113;
  wire popcount35_vg2l_core_117;
  wire popcount35_vg2l_core_119_not;
  wire popcount35_vg2l_core_120;
  wire popcount35_vg2l_core_123;
  wire popcount35_vg2l_core_124;
  wire popcount35_vg2l_core_125;
  wire popcount35_vg2l_core_126;
  wire popcount35_vg2l_core_127;
  wire popcount35_vg2l_core_128;
  wire popcount35_vg2l_core_129;
  wire popcount35_vg2l_core_130;
  wire popcount35_vg2l_core_132;
  wire popcount35_vg2l_core_133;
  wire popcount35_vg2l_core_135;
  wire popcount35_vg2l_core_136_not;
  wire popcount35_vg2l_core_138;
  wire popcount35_vg2l_core_140;
  wire popcount35_vg2l_core_143;
  wire popcount35_vg2l_core_145;
  wire popcount35_vg2l_core_148;
  wire popcount35_vg2l_core_149;
  wire popcount35_vg2l_core_150;
  wire popcount35_vg2l_core_152;
  wire popcount35_vg2l_core_153;
  wire popcount35_vg2l_core_154;
  wire popcount35_vg2l_core_156;
  wire popcount35_vg2l_core_159;
  wire popcount35_vg2l_core_161;
  wire popcount35_vg2l_core_164;
  wire popcount35_vg2l_core_165;
  wire popcount35_vg2l_core_167;
  wire popcount35_vg2l_core_168;
  wire popcount35_vg2l_core_170;
  wire popcount35_vg2l_core_171;
  wire popcount35_vg2l_core_174;
  wire popcount35_vg2l_core_175;
  wire popcount35_vg2l_core_176;
  wire popcount35_vg2l_core_180_not;
  wire popcount35_vg2l_core_181;
  wire popcount35_vg2l_core_182;
  wire popcount35_vg2l_core_183;
  wire popcount35_vg2l_core_184;
  wire popcount35_vg2l_core_185_not;
  wire popcount35_vg2l_core_186;
  wire popcount35_vg2l_core_187;
  wire popcount35_vg2l_core_188;
  wire popcount35_vg2l_core_189;
  wire popcount35_vg2l_core_190;
  wire popcount35_vg2l_core_191;
  wire popcount35_vg2l_core_192;
  wire popcount35_vg2l_core_195;
  wire popcount35_vg2l_core_196_not;
  wire popcount35_vg2l_core_198;
  wire popcount35_vg2l_core_202;
  wire popcount35_vg2l_core_203;
  wire popcount35_vg2l_core_205_not;
  wire popcount35_vg2l_core_206;
  wire popcount35_vg2l_core_207;
  wire popcount35_vg2l_core_208;
  wire popcount35_vg2l_core_209;
  wire popcount35_vg2l_core_212;
  wire popcount35_vg2l_core_214;
  wire popcount35_vg2l_core_215;
  wire popcount35_vg2l_core_216;
  wire popcount35_vg2l_core_217;
  wire popcount35_vg2l_core_219;
  wire popcount35_vg2l_core_220;
  wire popcount35_vg2l_core_222;
  wire popcount35_vg2l_core_223;
  wire popcount35_vg2l_core_224;
  wire popcount35_vg2l_core_225;
  wire popcount35_vg2l_core_226;
  wire popcount35_vg2l_core_227;
  wire popcount35_vg2l_core_229;
  wire popcount35_vg2l_core_230;
  wire popcount35_vg2l_core_231;
  wire popcount35_vg2l_core_232;
  wire popcount35_vg2l_core_233;
  wire popcount35_vg2l_core_235;
  wire popcount35_vg2l_core_236;
  wire popcount35_vg2l_core_237;
  wire popcount35_vg2l_core_241;
  wire popcount35_vg2l_core_242;
  wire popcount35_vg2l_core_244;
  wire popcount35_vg2l_core_245;
  wire popcount35_vg2l_core_246;
  wire popcount35_vg2l_core_247;
  wire popcount35_vg2l_core_250;
  wire popcount35_vg2l_core_252;
  wire popcount35_vg2l_core_253;
  wire popcount35_vg2l_core_254;
  wire popcount35_vg2l_core_255;
  wire popcount35_vg2l_core_256;
  wire popcount35_vg2l_core_257;
  wire popcount35_vg2l_core_259;
  wire popcount35_vg2l_core_260;
  wire popcount35_vg2l_core_261;
  wire popcount35_vg2l_core_264;

  assign popcount35_vg2l_core_037 = ~input_a[18];
  assign popcount35_vg2l_core_038 = ~(input_a[34] ^ input_a[11]);
  assign popcount35_vg2l_core_041 = ~input_a[23];
  assign popcount35_vg2l_core_042 = ~(input_a[27] | input_a[15]);
  assign popcount35_vg2l_core_044 = ~input_a[14];
  assign popcount35_vg2l_core_046 = ~input_a[7];
  assign popcount35_vg2l_core_047 = ~(input_a[30] | input_a[10]);
  assign popcount35_vg2l_core_048_not = ~input_a[3];
  assign popcount35_vg2l_core_049 = input_a[22] | input_a[12];
  assign popcount35_vg2l_core_050 = input_a[16] & input_a[16];
  assign popcount35_vg2l_core_051 = input_a[2] | input_a[15];
  assign popcount35_vg2l_core_052 = input_a[3] ^ input_a[26];
  assign popcount35_vg2l_core_054 = ~(input_a[12] & input_a[23]);
  assign popcount35_vg2l_core_055 = input_a[17] | input_a[0];
  assign popcount35_vg2l_core_056 = ~input_a[22];
  assign popcount35_vg2l_core_057 = input_a[32] | input_a[14];
  assign popcount35_vg2l_core_058 = ~(input_a[13] ^ input_a[34]);
  assign popcount35_vg2l_core_060 = input_a[0] | input_a[9];
  assign popcount35_vg2l_core_061 = input_a[29] & input_a[17];
  assign popcount35_vg2l_core_062 = input_a[18] | input_a[17];
  assign popcount35_vg2l_core_065 = ~input_a[18];
  assign popcount35_vg2l_core_067 = input_a[5] ^ input_a[28];
  assign popcount35_vg2l_core_068 = input_a[26] ^ input_a[2];
  assign popcount35_vg2l_core_069 = ~(input_a[21] | input_a[11]);
  assign popcount35_vg2l_core_071 = input_a[12] ^ input_a[30];
  assign popcount35_vg2l_core_072 = ~(input_a[1] & input_a[31]);
  assign popcount35_vg2l_core_073 = ~(input_a[3] | input_a[10]);
  assign popcount35_vg2l_core_075_not = ~input_a[19];
  assign popcount35_vg2l_core_076 = ~(input_a[34] | input_a[32]);
  assign popcount35_vg2l_core_077 = ~(input_a[16] & input_a[33]);
  assign popcount35_vg2l_core_079 = input_a[31] ^ input_a[30];
  assign popcount35_vg2l_core_080 = ~(input_a[12] ^ input_a[13]);
  assign popcount35_vg2l_core_081 = input_a[15] | input_a[17];
  assign popcount35_vg2l_core_083 = ~input_a[26];
  assign popcount35_vg2l_core_084 = input_a[29] ^ input_a[17];
  assign popcount35_vg2l_core_085 = ~(input_a[13] ^ input_a[24]);
  assign popcount35_vg2l_core_088 = ~(input_a[20] ^ input_a[32]);
  assign popcount35_vg2l_core_089 = input_a[34] & input_a[23];
  assign popcount35_vg2l_core_090 = ~input_a[27];
  assign popcount35_vg2l_core_093 = input_a[24] | input_a[29];
  assign popcount35_vg2l_core_097 = ~input_a[2];
  assign popcount35_vg2l_core_098 = ~input_a[28];
  assign popcount35_vg2l_core_100 = ~(input_a[2] | input_a[26]);
  assign popcount35_vg2l_core_103 = input_a[34] ^ input_a[6];
  assign popcount35_vg2l_core_104 = input_a[19] ^ input_a[26];
  assign popcount35_vg2l_core_105 = input_a[6] & input_a[31];
  assign popcount35_vg2l_core_107 = input_a[32] | input_a[16];
  assign popcount35_vg2l_core_108 = input_a[18] ^ input_a[27];
  assign popcount35_vg2l_core_109 = ~(input_a[4] ^ input_a[23]);
  assign popcount35_vg2l_core_112 = ~(input_a[16] | input_a[32]);
  assign popcount35_vg2l_core_113 = ~(input_a[9] ^ input_a[21]);
  assign popcount35_vg2l_core_117 = ~(input_a[28] | input_a[15]);
  assign popcount35_vg2l_core_119_not = ~input_a[8];
  assign popcount35_vg2l_core_120 = ~(input_a[34] ^ input_a[13]);
  assign popcount35_vg2l_core_123 = input_a[8] ^ input_a[33];
  assign popcount35_vg2l_core_124 = ~(input_a[25] & input_a[6]);
  assign popcount35_vg2l_core_125 = ~input_a[22];
  assign popcount35_vg2l_core_126 = input_a[21] | input_a[14];
  assign popcount35_vg2l_core_127 = ~input_a[15];
  assign popcount35_vg2l_core_128 = ~input_a[13];
  assign popcount35_vg2l_core_129 = ~(input_a[13] & input_a[14]);
  assign popcount35_vg2l_core_130 = ~input_a[10];
  assign popcount35_vg2l_core_132 = input_a[21] & input_a[14];
  assign popcount35_vg2l_core_133 = ~input_a[10];
  assign popcount35_vg2l_core_135 = ~(input_a[25] ^ input_a[24]);
  assign popcount35_vg2l_core_136_not = ~input_a[19];
  assign popcount35_vg2l_core_138 = ~(input_a[27] & input_a[3]);
  assign popcount35_vg2l_core_140 = input_a[30] | input_a[30];
  assign popcount35_vg2l_core_143 = input_a[24] ^ input_a[34];
  assign popcount35_vg2l_core_145 = input_a[23] ^ input_a[10];
  assign popcount35_vg2l_core_148 = ~(input_a[28] | input_a[3]);
  assign popcount35_vg2l_core_149 = input_a[20] | input_a[23];
  assign popcount35_vg2l_core_150 = ~(input_a[7] & input_a[7]);
  assign popcount35_vg2l_core_152 = input_a[4] | input_a[16];
  assign popcount35_vg2l_core_153 = input_a[13] & input_a[16];
  assign popcount35_vg2l_core_154 = ~(input_a[2] & input_a[8]);
  assign popcount35_vg2l_core_156 = input_a[3] & input_a[13];
  assign popcount35_vg2l_core_159 = ~input_a[2];
  assign popcount35_vg2l_core_161 = ~(input_a[26] & input_a[8]);
  assign popcount35_vg2l_core_164 = ~(input_a[16] | input_a[4]);
  assign popcount35_vg2l_core_165 = input_a[5] ^ input_a[4];
  assign popcount35_vg2l_core_167 = input_a[4] ^ input_a[17];
  assign popcount35_vg2l_core_168 = input_a[33] ^ input_a[15];
  assign popcount35_vg2l_core_170 = input_a[20] & input_a[29];
  assign popcount35_vg2l_core_171 = ~(input_a[33] & input_a[33]);
  assign popcount35_vg2l_core_174 = ~input_a[10];
  assign popcount35_vg2l_core_175 = ~(input_a[5] & input_a[15]);
  assign popcount35_vg2l_core_176 = ~(input_a[7] | input_a[6]);
  assign popcount35_vg2l_core_180_not = ~input_a[32];
  assign popcount35_vg2l_core_181 = ~(input_a[22] ^ input_a[20]);
  assign popcount35_vg2l_core_182 = ~(input_a[21] | input_a[23]);
  assign popcount35_vg2l_core_183 = input_a[4] ^ input_a[14];
  assign popcount35_vg2l_core_184 = ~input_a[1];
  assign popcount35_vg2l_core_185_not = ~input_a[10];
  assign popcount35_vg2l_core_186 = ~(input_a[0] & input_a[15]);
  assign popcount35_vg2l_core_187 = ~input_a[16];
  assign popcount35_vg2l_core_188 = ~(input_a[8] & input_a[26]);
  assign popcount35_vg2l_core_189 = ~input_a[20];
  assign popcount35_vg2l_core_190 = input_a[26] | input_a[33];
  assign popcount35_vg2l_core_191 = input_a[8] | input_a[1];
  assign popcount35_vg2l_core_192 = ~(input_a[23] | input_a[16]);
  assign popcount35_vg2l_core_195 = ~(input_a[16] & input_a[9]);
  assign popcount35_vg2l_core_196_not = ~input_a[28];
  assign popcount35_vg2l_core_198 = input_a[21] ^ input_a[25];
  assign popcount35_vg2l_core_202 = input_a[15] ^ input_a[14];
  assign popcount35_vg2l_core_203 = ~input_a[31];
  assign popcount35_vg2l_core_205_not = ~input_a[13];
  assign popcount35_vg2l_core_206 = input_a[1] & input_a[17];
  assign popcount35_vg2l_core_207 = input_a[1] ^ input_a[20];
  assign popcount35_vg2l_core_208 = ~(input_a[2] ^ input_a[22]);
  assign popcount35_vg2l_core_209 = ~input_a[9];
  assign popcount35_vg2l_core_212 = input_a[18] | input_a[34];
  assign popcount35_vg2l_core_214 = input_a[9] ^ input_a[33];
  assign popcount35_vg2l_core_215 = ~(input_a[20] | input_a[30]);
  assign popcount35_vg2l_core_216 = ~(input_a[29] & input_a[32]);
  assign popcount35_vg2l_core_217 = input_a[11] ^ input_a[34];
  assign popcount35_vg2l_core_219 = input_a[6] ^ input_a[19];
  assign popcount35_vg2l_core_220 = input_a[12] | input_a[25];
  assign popcount35_vg2l_core_222 = input_a[7] ^ input_a[31];
  assign popcount35_vg2l_core_223 = ~(input_a[29] ^ input_a[6]);
  assign popcount35_vg2l_core_224 = input_a[27] | input_a[26];
  assign popcount35_vg2l_core_225 = input_a[29] & input_a[12];
  assign popcount35_vg2l_core_226 = ~(input_a[8] ^ input_a[4]);
  assign popcount35_vg2l_core_227 = input_a[6] & input_a[32];
  assign popcount35_vg2l_core_229 = input_a[25] | input_a[33];
  assign popcount35_vg2l_core_230 = ~input_a[5];
  assign popcount35_vg2l_core_231 = ~(input_a[33] & input_a[13]);
  assign popcount35_vg2l_core_232 = input_a[6] ^ input_a[18];
  assign popcount35_vg2l_core_233 = ~(input_a[7] | input_a[1]);
  assign popcount35_vg2l_core_235 = input_a[9] & input_a[30];
  assign popcount35_vg2l_core_236 = ~(input_a[14] | input_a[11]);
  assign popcount35_vg2l_core_237 = ~input_a[31];
  assign popcount35_vg2l_core_241 = input_a[29] | input_a[20];
  assign popcount35_vg2l_core_242 = ~(input_a[30] ^ input_a[18]);
  assign popcount35_vg2l_core_244 = input_a[16] | input_a[19];
  assign popcount35_vg2l_core_245 = ~(input_a[22] ^ input_a[1]);
  assign popcount35_vg2l_core_246 = ~(input_a[24] ^ input_a[4]);
  assign popcount35_vg2l_core_247 = ~(input_a[34] & input_a[2]);
  assign popcount35_vg2l_core_250 = ~(input_a[7] & input_a[20]);
  assign popcount35_vg2l_core_252 = ~(input_a[28] | input_a[21]);
  assign popcount35_vg2l_core_253 = input_a[14] ^ input_a[24];
  assign popcount35_vg2l_core_254 = ~(input_a[29] & input_a[13]);
  assign popcount35_vg2l_core_255 = input_a[34] | input_a[33];
  assign popcount35_vg2l_core_256 = ~(input_a[23] & input_a[10]);
  assign popcount35_vg2l_core_257 = input_a[31] | input_a[31];
  assign popcount35_vg2l_core_259 = input_a[7] ^ input_a[4];
  assign popcount35_vg2l_core_260 = ~input_a[14];
  assign popcount35_vg2l_core_261 = ~(input_a[0] & input_a[32]);
  assign popcount35_vg2l_core_264 = input_a[34] ^ input_a[32];

  assign popcount35_vg2l_out[0] = 1'b0;
  assign popcount35_vg2l_out[1] = 1'b0;
  assign popcount35_vg2l_out[2] = 1'b0;
  assign popcount35_vg2l_out[3] = input_a[3];
  assign popcount35_vg2l_out[4] = 1'b0;
  assign popcount35_vg2l_out[5] = input_a[26];
endmodule