// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.16373
// WCE=20.0
// EP=0.932979%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_6to5(input [23:0] input_a, output [4:0] popcount24_6to5_out);
  wire popcount24_6to5_core_028;
  wire popcount24_6to5_core_030;
  wire popcount24_6to5_core_031_not;
  wire popcount24_6to5_core_032;
  wire popcount24_6to5_core_033;
  wire popcount24_6to5_core_036;
  wire popcount24_6to5_core_038;
  wire popcount24_6to5_core_039;
  wire popcount24_6to5_core_041_not;
  wire popcount24_6to5_core_044;
  wire popcount24_6to5_core_046;
  wire popcount24_6to5_core_048;
  wire popcount24_6to5_core_049;
  wire popcount24_6to5_core_052;
  wire popcount24_6to5_core_053;
  wire popcount24_6to5_core_054;
  wire popcount24_6to5_core_056;
  wire popcount24_6to5_core_059;
  wire popcount24_6to5_core_060;
  wire popcount24_6to5_core_062;
  wire popcount24_6to5_core_064;
  wire popcount24_6to5_core_065;
  wire popcount24_6to5_core_066;
  wire popcount24_6to5_core_067;
  wire popcount24_6to5_core_069;
  wire popcount24_6to5_core_070;
  wire popcount24_6to5_core_071;
  wire popcount24_6to5_core_072;
  wire popcount24_6to5_core_073;
  wire popcount24_6to5_core_074;
  wire popcount24_6to5_core_075;
  wire popcount24_6to5_core_076;
  wire popcount24_6to5_core_078;
  wire popcount24_6to5_core_082;
  wire popcount24_6to5_core_084;
  wire popcount24_6to5_core_086;
  wire popcount24_6to5_core_087;
  wire popcount24_6to5_core_088;
  wire popcount24_6to5_core_089;
  wire popcount24_6to5_core_090;
  wire popcount24_6to5_core_091;
  wire popcount24_6to5_core_092;
  wire popcount24_6to5_core_094;
  wire popcount24_6to5_core_096;
  wire popcount24_6to5_core_098;
  wire popcount24_6to5_core_100;
  wire popcount24_6to5_core_101;
  wire popcount24_6to5_core_102;
  wire popcount24_6to5_core_103;
  wire popcount24_6to5_core_104;
  wire popcount24_6to5_core_105;
  wire popcount24_6to5_core_107;
  wire popcount24_6to5_core_108;
  wire popcount24_6to5_core_109;
  wire popcount24_6to5_core_110;
  wire popcount24_6to5_core_111;
  wire popcount24_6to5_core_116;
  wire popcount24_6to5_core_118;
  wire popcount24_6to5_core_119;
  wire popcount24_6to5_core_120;
  wire popcount24_6to5_core_122;
  wire popcount24_6to5_core_124;
  wire popcount24_6to5_core_127;
  wire popcount24_6to5_core_129;
  wire popcount24_6to5_core_130;
  wire popcount24_6to5_core_133;
  wire popcount24_6to5_core_134_not;
  wire popcount24_6to5_core_135;
  wire popcount24_6to5_core_136;
  wire popcount24_6to5_core_137;
  wire popcount24_6to5_core_138;
  wire popcount24_6to5_core_140;
  wire popcount24_6to5_core_141;
  wire popcount24_6to5_core_143;
  wire popcount24_6to5_core_144;
  wire popcount24_6to5_core_146;
  wire popcount24_6to5_core_147;
  wire popcount24_6to5_core_149;
  wire popcount24_6to5_core_152_not;
  wire popcount24_6to5_core_153;
  wire popcount24_6to5_core_154;
  wire popcount24_6to5_core_156;
  wire popcount24_6to5_core_159;
  wire popcount24_6to5_core_160;
  wire popcount24_6to5_core_161;
  wire popcount24_6to5_core_162;
  wire popcount24_6to5_core_163;
  wire popcount24_6to5_core_164;
  wire popcount24_6to5_core_165;
  wire popcount24_6to5_core_166;
  wire popcount24_6to5_core_167_not;
  wire popcount24_6to5_core_168;
  wire popcount24_6to5_core_169;
  wire popcount24_6to5_core_170;
  wire popcount24_6to5_core_176;
  wire popcount24_6to5_core_177;

  assign popcount24_6to5_core_028 = input_a[6] | input_a[16];
  assign popcount24_6to5_core_030 = ~input_a[6];
  assign popcount24_6to5_core_031_not = ~input_a[9];
  assign popcount24_6to5_core_032 = ~(input_a[12] | input_a[3]);
  assign popcount24_6to5_core_033 = input_a[4] & input_a[22];
  assign popcount24_6to5_core_036 = ~(input_a[22] ^ input_a[20]);
  assign popcount24_6to5_core_038 = input_a[15] & input_a[10];
  assign popcount24_6to5_core_039 = ~(input_a[9] | input_a[22]);
  assign popcount24_6to5_core_041_not = ~input_a[12];
  assign popcount24_6to5_core_044 = ~input_a[12];
  assign popcount24_6to5_core_046 = input_a[3] & input_a[13];
  assign popcount24_6to5_core_048 = ~(input_a[23] & input_a[15]);
  assign popcount24_6to5_core_049 = input_a[15] & input_a[3];
  assign popcount24_6to5_core_052 = ~(input_a[0] | input_a[6]);
  assign popcount24_6to5_core_053 = input_a[15] | input_a[17];
  assign popcount24_6to5_core_054 = ~(input_a[23] & input_a[15]);
  assign popcount24_6to5_core_056 = ~input_a[9];
  assign popcount24_6to5_core_059 = input_a[13] & input_a[11];
  assign popcount24_6to5_core_060 = input_a[18] ^ input_a[12];
  assign popcount24_6to5_core_062 = ~(input_a[4] | input_a[8]);
  assign popcount24_6to5_core_064 = ~(input_a[14] | input_a[7]);
  assign popcount24_6to5_core_065 = ~(input_a[15] | input_a[20]);
  assign popcount24_6to5_core_066 = ~(input_a[22] ^ input_a[21]);
  assign popcount24_6to5_core_067 = input_a[19] | input_a[3];
  assign popcount24_6to5_core_069 = input_a[13] | input_a[15];
  assign popcount24_6to5_core_070 = input_a[4] ^ input_a[8];
  assign popcount24_6to5_core_071 = ~(input_a[8] | input_a[6]);
  assign popcount24_6to5_core_072 = ~(input_a[6] | input_a[11]);
  assign popcount24_6to5_core_073 = input_a[4] & input_a[22];
  assign popcount24_6to5_core_074 = input_a[0] | input_a[7];
  assign popcount24_6to5_core_075 = input_a[18] & input_a[9];
  assign popcount24_6to5_core_076 = ~(input_a[14] & input_a[14]);
  assign popcount24_6to5_core_078 = input_a[12] & input_a[2];
  assign popcount24_6to5_core_082 = ~(input_a[21] | input_a[4]);
  assign popcount24_6to5_core_084 = ~input_a[17];
  assign popcount24_6to5_core_086 = ~(input_a[15] & input_a[20]);
  assign popcount24_6to5_core_087 = ~input_a[6];
  assign popcount24_6to5_core_088 = input_a[15] & input_a[20];
  assign popcount24_6to5_core_089 = ~(input_a[2] & input_a[10]);
  assign popcount24_6to5_core_090 = ~(input_a[11] | input_a[8]);
  assign popcount24_6to5_core_091 = ~(input_a[7] ^ input_a[14]);
  assign popcount24_6to5_core_092 = ~(input_a[18] & input_a[1]);
  assign popcount24_6to5_core_094 = ~(input_a[5] | input_a[22]);
  assign popcount24_6to5_core_096 = input_a[17] ^ input_a[4];
  assign popcount24_6to5_core_098 = ~(input_a[10] | input_a[20]);
  assign popcount24_6to5_core_100 = ~input_a[15];
  assign popcount24_6to5_core_101 = ~(input_a[13] | input_a[3]);
  assign popcount24_6to5_core_102 = ~(input_a[11] | input_a[13]);
  assign popcount24_6to5_core_103 = ~(input_a[5] ^ input_a[7]);
  assign popcount24_6to5_core_104 = input_a[11] | input_a[3];
  assign popcount24_6to5_core_105 = input_a[20] ^ input_a[5];
  assign popcount24_6to5_core_107 = ~(input_a[4] & input_a[4]);
  assign popcount24_6to5_core_108 = input_a[21] | input_a[16];
  assign popcount24_6to5_core_109 = input_a[21] & input_a[5];
  assign popcount24_6to5_core_110 = input_a[10] & input_a[16];
  assign popcount24_6to5_core_111 = input_a[16] & input_a[11];
  assign popcount24_6to5_core_116 = input_a[18] | input_a[14];
  assign popcount24_6to5_core_118 = input_a[21] | input_a[6];
  assign popcount24_6to5_core_119 = ~(input_a[21] | input_a[16]);
  assign popcount24_6to5_core_120 = input_a[14] & input_a[11];
  assign popcount24_6to5_core_122 = input_a[1] | input_a[16];
  assign popcount24_6to5_core_124 = input_a[16] | input_a[15];
  assign popcount24_6to5_core_127 = input_a[1] | input_a[19];
  assign popcount24_6to5_core_129 = input_a[7] | input_a[15];
  assign popcount24_6to5_core_130 = ~input_a[4];
  assign popcount24_6to5_core_133 = input_a[13] ^ input_a[10];
  assign popcount24_6to5_core_134_not = ~input_a[7];
  assign popcount24_6to5_core_135 = ~(input_a[7] ^ input_a[11]);
  assign popcount24_6to5_core_136 = input_a[21] & input_a[0];
  assign popcount24_6to5_core_137 = input_a[15] | input_a[15];
  assign popcount24_6to5_core_138 = input_a[13] | input_a[11];
  assign popcount24_6to5_core_140 = input_a[23] | input_a[7];
  assign popcount24_6to5_core_141 = input_a[1] & input_a[20];
  assign popcount24_6to5_core_143 = input_a[13] | input_a[0];
  assign popcount24_6to5_core_144 = ~(input_a[4] & input_a[4]);
  assign popcount24_6to5_core_146 = ~input_a[22];
  assign popcount24_6to5_core_147 = ~(input_a[3] & input_a[17]);
  assign popcount24_6to5_core_149 = input_a[19] ^ input_a[16];
  assign popcount24_6to5_core_152_not = ~input_a[17];
  assign popcount24_6to5_core_153 = ~(input_a[14] | input_a[23]);
  assign popcount24_6to5_core_154 = input_a[14] & input_a[12];
  assign popcount24_6to5_core_156 = ~(input_a[4] & input_a[10]);
  assign popcount24_6to5_core_159 = ~input_a[18];
  assign popcount24_6to5_core_160 = ~input_a[8];
  assign popcount24_6to5_core_161 = input_a[17] & input_a[16];
  assign popcount24_6to5_core_162 = ~(input_a[6] & input_a[0]);
  assign popcount24_6to5_core_163 = ~(input_a[23] & input_a[2]);
  assign popcount24_6to5_core_164 = ~(input_a[8] ^ input_a[0]);
  assign popcount24_6to5_core_165 = input_a[11] ^ input_a[4];
  assign popcount24_6to5_core_166 = input_a[23] ^ input_a[2];
  assign popcount24_6to5_core_167_not = ~input_a[1];
  assign popcount24_6to5_core_168 = ~(input_a[6] | input_a[13]);
  assign popcount24_6to5_core_169 = input_a[15] | input_a[14];
  assign popcount24_6to5_core_170 = ~(input_a[6] ^ input_a[18]);
  assign popcount24_6to5_core_176 = input_a[9] & input_a[16];
  assign popcount24_6to5_core_177 = ~(input_a[12] | input_a[14]);

  assign popcount24_6to5_out[0] = input_a[5];
  assign popcount24_6to5_out[1] = input_a[6];
  assign popcount24_6to5_out[2] = input_a[21];
  assign popcount24_6to5_out[3] = input_a[0];
  assign popcount24_6to5_out[4] = 1'b0;
endmodule