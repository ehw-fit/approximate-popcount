// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.79266
// WCE=13.0
// EP=0.827212%
// Printed PDK parameters:
//  Area=45850963.0
//  Delay=63942064.0
//  Power=2230000.0

module popcount36_vanw(input [35:0] input_a, output [5:0] popcount36_vanw_out);
  wire popcount36_vanw_core_038;
  wire popcount36_vanw_core_040;
  wire popcount36_vanw_core_041;
  wire popcount36_vanw_core_042;
  wire popcount36_vanw_core_046;
  wire popcount36_vanw_core_047;
  wire popcount36_vanw_core_049;
  wire popcount36_vanw_core_050;
  wire popcount36_vanw_core_051;
  wire popcount36_vanw_core_052;
  wire popcount36_vanw_core_053;
  wire popcount36_vanw_core_054;
  wire popcount36_vanw_core_055;
  wire popcount36_vanw_core_057;
  wire popcount36_vanw_core_058;
  wire popcount36_vanw_core_059;
  wire popcount36_vanw_core_060;
  wire popcount36_vanw_core_061;
  wire popcount36_vanw_core_062;
  wire popcount36_vanw_core_063;
  wire popcount36_vanw_core_065;
  wire popcount36_vanw_core_067;
  wire popcount36_vanw_core_068;
  wire popcount36_vanw_core_069;
  wire popcount36_vanw_core_071;
  wire popcount36_vanw_core_075;
  wire popcount36_vanw_core_076;
  wire popcount36_vanw_core_078;
  wire popcount36_vanw_core_079;
  wire popcount36_vanw_core_080;
  wire popcount36_vanw_core_081;
  wire popcount36_vanw_core_082;
  wire popcount36_vanw_core_083;
  wire popcount36_vanw_core_084;
  wire popcount36_vanw_core_085;
  wire popcount36_vanw_core_086;
  wire popcount36_vanw_core_087;
  wire popcount36_vanw_core_091;
  wire popcount36_vanw_core_092;
  wire popcount36_vanw_core_093;
  wire popcount36_vanw_core_094;
  wire popcount36_vanw_core_095;
  wire popcount36_vanw_core_096;
  wire popcount36_vanw_core_097;
  wire popcount36_vanw_core_099;
  wire popcount36_vanw_core_100;
  wire popcount36_vanw_core_101;
  wire popcount36_vanw_core_102;
  wire popcount36_vanw_core_103;
  wire popcount36_vanw_core_104;
  wire popcount36_vanw_core_105;
  wire popcount36_vanw_core_107;
  wire popcount36_vanw_core_108;
  wire popcount36_vanw_core_109;
  wire popcount36_vanw_core_110;
  wire popcount36_vanw_core_111;
  wire popcount36_vanw_core_112;
  wire popcount36_vanw_core_113;
  wire popcount36_vanw_core_114;
  wire popcount36_vanw_core_117;
  wire popcount36_vanw_core_118;
  wire popcount36_vanw_core_120;
  wire popcount36_vanw_core_121;
  wire popcount36_vanw_core_122;
  wire popcount36_vanw_core_124;
  wire popcount36_vanw_core_126;
  wire popcount36_vanw_core_128;
  wire popcount36_vanw_core_129;
  wire popcount36_vanw_core_130;
  wire popcount36_vanw_core_131;
  wire popcount36_vanw_core_132;
  wire popcount36_vanw_core_133;
  wire popcount36_vanw_core_135;
  wire popcount36_vanw_core_138;
  wire popcount36_vanw_core_139_not;
  wire popcount36_vanw_core_141_not;
  wire popcount36_vanw_core_142;
  wire popcount36_vanw_core_143;
  wire popcount36_vanw_core_146;
  wire popcount36_vanw_core_147;
  wire popcount36_vanw_core_148;
  wire popcount36_vanw_core_149;
  wire popcount36_vanw_core_150;
  wire popcount36_vanw_core_151;
  wire popcount36_vanw_core_155;
  wire popcount36_vanw_core_156;
  wire popcount36_vanw_core_157;
  wire popcount36_vanw_core_158;
  wire popcount36_vanw_core_160;
  wire popcount36_vanw_core_162;
  wire popcount36_vanw_core_164;
  wire popcount36_vanw_core_165;
  wire popcount36_vanw_core_166;
  wire popcount36_vanw_core_168;
  wire popcount36_vanw_core_169;
  wire popcount36_vanw_core_170;
  wire popcount36_vanw_core_171;
  wire popcount36_vanw_core_172;
  wire popcount36_vanw_core_173;
  wire popcount36_vanw_core_174;
  wire popcount36_vanw_core_175;
  wire popcount36_vanw_core_177;
  wire popcount36_vanw_core_181;
  wire popcount36_vanw_core_182;
  wire popcount36_vanw_core_183;
  wire popcount36_vanw_core_184;
  wire popcount36_vanw_core_185;
  wire popcount36_vanw_core_188;
  wire popcount36_vanw_core_189;
  wire popcount36_vanw_core_190;
  wire popcount36_vanw_core_191;
  wire popcount36_vanw_core_192;
  wire popcount36_vanw_core_193;
  wire popcount36_vanw_core_195;
  wire popcount36_vanw_core_198;
  wire popcount36_vanw_core_200;
  wire popcount36_vanw_core_201;
  wire popcount36_vanw_core_202;
  wire popcount36_vanw_core_203;
  wire popcount36_vanw_core_205;
  wire popcount36_vanw_core_206;
  wire popcount36_vanw_core_207;
  wire popcount36_vanw_core_208;
  wire popcount36_vanw_core_209;
  wire popcount36_vanw_core_210;
  wire popcount36_vanw_core_211;
  wire popcount36_vanw_core_213;
  wire popcount36_vanw_core_215;
  wire popcount36_vanw_core_216;
  wire popcount36_vanw_core_217;
  wire popcount36_vanw_core_222_not;
  wire popcount36_vanw_core_223;
  wire popcount36_vanw_core_224;
  wire popcount36_vanw_core_225;
  wire popcount36_vanw_core_227;
  wire popcount36_vanw_core_228;
  wire popcount36_vanw_core_230;
  wire popcount36_vanw_core_235;
  wire popcount36_vanw_core_236;
  wire popcount36_vanw_core_237;
  wire popcount36_vanw_core_238;
  wire popcount36_vanw_core_239;
  wire popcount36_vanw_core_241;
  wire popcount36_vanw_core_243;
  wire popcount36_vanw_core_244;
  wire popcount36_vanw_core_245;
  wire popcount36_vanw_core_247;
  wire popcount36_vanw_core_249;
  wire popcount36_vanw_core_251;
  wire popcount36_vanw_core_257;
  wire popcount36_vanw_core_258;
  wire popcount36_vanw_core_259;
  wire popcount36_vanw_core_260;
  wire popcount36_vanw_core_261;
  wire popcount36_vanw_core_262;
  wire popcount36_vanw_core_263;
  wire popcount36_vanw_core_264;
  wire popcount36_vanw_core_265;
  wire popcount36_vanw_core_266;
  wire popcount36_vanw_core_267;
  wire popcount36_vanw_core_270;
  wire popcount36_vanw_core_275;

  assign popcount36_vanw_core_038 = input_a[0] & input_a[26];
  assign popcount36_vanw_core_040 = input_a[16] ^ input_a[31];
  assign popcount36_vanw_core_041 = input_a[2] & input_a[1];
  assign popcount36_vanw_core_042 = input_a[27] | input_a[1];
  assign popcount36_vanw_core_046 = popcount36_vanw_core_041 | popcount36_vanw_core_038;
  assign popcount36_vanw_core_047 = ~(input_a[1] ^ input_a[3]);
  assign popcount36_vanw_core_049 = input_a[4] ^ input_a[5];
  assign popcount36_vanw_core_050 = input_a[4] & input_a[5];
  assign popcount36_vanw_core_051 = ~(input_a[7] & input_a[8]);
  assign popcount36_vanw_core_052 = input_a[7] & input_a[8];
  assign popcount36_vanw_core_053 = input_a[6] ^ popcount36_vanw_core_051;
  assign popcount36_vanw_core_054 = ~(input_a[27] ^ input_a[15]);
  assign popcount36_vanw_core_055 = popcount36_vanw_core_052 | input_a[6];
  assign popcount36_vanw_core_057 = ~input_a[4];
  assign popcount36_vanw_core_058 = popcount36_vanw_core_049 & popcount36_vanw_core_053;
  assign popcount36_vanw_core_059 = popcount36_vanw_core_050 ^ popcount36_vanw_core_055;
  assign popcount36_vanw_core_060 = popcount36_vanw_core_050 & popcount36_vanw_core_055;
  assign popcount36_vanw_core_061 = popcount36_vanw_core_059 ^ popcount36_vanw_core_058;
  assign popcount36_vanw_core_062 = input_a[6] & popcount36_vanw_core_058;
  assign popcount36_vanw_core_063 = popcount36_vanw_core_060 | popcount36_vanw_core_062;
  assign popcount36_vanw_core_065 = ~input_a[26];
  assign popcount36_vanw_core_067 = ~input_a[14];
  assign popcount36_vanw_core_068 = popcount36_vanw_core_046 ^ popcount36_vanw_core_061;
  assign popcount36_vanw_core_069 = popcount36_vanw_core_046 & popcount36_vanw_core_061;
  assign popcount36_vanw_core_071 = ~(input_a[27] | input_a[33]);
  assign popcount36_vanw_core_075 = popcount36_vanw_core_063 | popcount36_vanw_core_069;
  assign popcount36_vanw_core_076 = input_a[28] | input_a[12];
  assign popcount36_vanw_core_078 = input_a[15] ^ input_a[31];
  assign popcount36_vanw_core_079 = ~(input_a[2] | input_a[28]);
  assign popcount36_vanw_core_080 = ~(input_a[24] ^ input_a[1]);
  assign popcount36_vanw_core_081 = input_a[9] & input_a[10];
  assign popcount36_vanw_core_082 = input_a[6] & input_a[14];
  assign popcount36_vanw_core_083 = input_a[21] & input_a[12];
  assign popcount36_vanw_core_084 = ~(input_a[8] | input_a[35]);
  assign popcount36_vanw_core_085 = ~(input_a[6] & input_a[4]);
  assign popcount36_vanw_core_086 = popcount36_vanw_core_081 | popcount36_vanw_core_083;
  assign popcount36_vanw_core_087 = ~input_a[9];
  assign popcount36_vanw_core_091 = input_a[13] ^ input_a[14];
  assign popcount36_vanw_core_092 = input_a[13] & input_a[14];
  assign popcount36_vanw_core_093 = ~(input_a[16] & input_a[17]);
  assign popcount36_vanw_core_094 = input_a[16] & input_a[17];
  assign popcount36_vanw_core_095 = input_a[15] ^ popcount36_vanw_core_093;
  assign popcount36_vanw_core_096 = input_a[23] & input_a[22];
  assign popcount36_vanw_core_097 = popcount36_vanw_core_094 | input_a[15];
  assign popcount36_vanw_core_099 = popcount36_vanw_core_091 ^ popcount36_vanw_core_095;
  assign popcount36_vanw_core_100 = popcount36_vanw_core_091 & popcount36_vanw_core_095;
  assign popcount36_vanw_core_101 = popcount36_vanw_core_092 ^ popcount36_vanw_core_097;
  assign popcount36_vanw_core_102 = popcount36_vanw_core_092 & popcount36_vanw_core_097;
  assign popcount36_vanw_core_103 = popcount36_vanw_core_101 ^ popcount36_vanw_core_100;
  assign popcount36_vanw_core_104 = input_a[15] & popcount36_vanw_core_100;
  assign popcount36_vanw_core_105 = popcount36_vanw_core_102 | popcount36_vanw_core_104;
  assign popcount36_vanw_core_107 = ~(input_a[7] | input_a[19]);
  assign popcount36_vanw_core_108 = input_a[27] | input_a[1];
  assign popcount36_vanw_core_109 = input_a[28] & popcount36_vanw_core_099;
  assign popcount36_vanw_core_110 = popcount36_vanw_core_086 ^ popcount36_vanw_core_103;
  assign popcount36_vanw_core_111 = popcount36_vanw_core_086 & popcount36_vanw_core_103;
  assign popcount36_vanw_core_112 = popcount36_vanw_core_110 ^ popcount36_vanw_core_109;
  assign popcount36_vanw_core_113 = popcount36_vanw_core_110 & popcount36_vanw_core_109;
  assign popcount36_vanw_core_114 = popcount36_vanw_core_111 | popcount36_vanw_core_113;
  assign popcount36_vanw_core_117 = popcount36_vanw_core_105 | popcount36_vanw_core_114;
  assign popcount36_vanw_core_118 = input_a[7] | input_a[2];
  assign popcount36_vanw_core_120 = ~input_a[35];
  assign popcount36_vanw_core_121 = ~input_a[18];
  assign popcount36_vanw_core_122 = ~input_a[2];
  assign popcount36_vanw_core_124 = popcount36_vanw_core_068 ^ popcount36_vanw_core_112;
  assign popcount36_vanw_core_126 = ~popcount36_vanw_core_124;
  assign popcount36_vanw_core_128 = popcount36_vanw_core_068 | popcount36_vanw_core_124;
  assign popcount36_vanw_core_129 = popcount36_vanw_core_075 ^ popcount36_vanw_core_117;
  assign popcount36_vanw_core_130 = popcount36_vanw_core_075 & popcount36_vanw_core_117;
  assign popcount36_vanw_core_131 = popcount36_vanw_core_129 ^ popcount36_vanw_core_128;
  assign popcount36_vanw_core_132 = popcount36_vanw_core_129 & popcount36_vanw_core_128;
  assign popcount36_vanw_core_133 = popcount36_vanw_core_130 | popcount36_vanw_core_132;
  assign popcount36_vanw_core_135 = ~(input_a[19] ^ input_a[25]);
  assign popcount36_vanw_core_138 = ~(input_a[10] & input_a[11]);
  assign popcount36_vanw_core_139_not = ~input_a[8];
  assign popcount36_vanw_core_141_not = ~input_a[0];
  assign popcount36_vanw_core_142 = input_a[27] | input_a[34];
  assign popcount36_vanw_core_143 = ~(input_a[16] & input_a[5]);
  assign popcount36_vanw_core_146 = ~(input_a[31] ^ input_a[30]);
  assign popcount36_vanw_core_147 = ~(input_a[3] | input_a[20]);
  assign popcount36_vanw_core_148 = input_a[16] & input_a[28];
  assign popcount36_vanw_core_149 = ~input_a[4];
  assign popcount36_vanw_core_150 = ~(input_a[19] & input_a[20]);
  assign popcount36_vanw_core_151 = input_a[19] & input_a[20];
  assign popcount36_vanw_core_155 = ~(input_a[13] ^ input_a[10]);
  assign popcount36_vanw_core_156 = input_a[29] & input_a[23];
  assign popcount36_vanw_core_157 = input_a[5] | input_a[20];
  assign popcount36_vanw_core_158 = input_a[24] & input_a[3];
  assign popcount36_vanw_core_160 = ~input_a[2];
  assign popcount36_vanw_core_162 = input_a[16] & input_a[12];
  assign popcount36_vanw_core_164 = input_a[5] ^ input_a[25];
  assign popcount36_vanw_core_165 = popcount36_vanw_core_156 | popcount36_vanw_core_158;
  assign popcount36_vanw_core_166 = ~(input_a[22] ^ input_a[28]);
  assign popcount36_vanw_core_168 = ~(input_a[18] & input_a[17]);
  assign popcount36_vanw_core_169 = input_a[16] & input_a[5];
  assign popcount36_vanw_core_170 = ~(input_a[20] & input_a[34]);
  assign popcount36_vanw_core_171 = input_a[35] & input_a[26];
  assign popcount36_vanw_core_172 = ~input_a[8];
  assign popcount36_vanw_core_173 = input_a[6] ^ input_a[23];
  assign popcount36_vanw_core_174 = popcount36_vanw_core_150 ^ popcount36_vanw_core_165;
  assign popcount36_vanw_core_175 = popcount36_vanw_core_150 & popcount36_vanw_core_165;
  assign popcount36_vanw_core_177 = input_a[0] & input_a[11];
  assign popcount36_vanw_core_181 = popcount36_vanw_core_151 | popcount36_vanw_core_175;
  assign popcount36_vanw_core_182 = input_a[21] ^ input_a[0];
  assign popcount36_vanw_core_183 = ~(input_a[23] ^ input_a[24]);
  assign popcount36_vanw_core_184 = input_a[15] & input_a[5];
  assign popcount36_vanw_core_185 = ~(input_a[3] & input_a[20]);
  assign popcount36_vanw_core_188 = ~(input_a[4] | input_a[24]);
  assign popcount36_vanw_core_189 = input_a[11] & input_a[30];
  assign popcount36_vanw_core_190 = ~(input_a[35] ^ input_a[5]);
  assign popcount36_vanw_core_191 = input_a[24] & input_a[31];
  assign popcount36_vanw_core_192 = input_a[27] | popcount36_vanw_core_189;
  assign popcount36_vanw_core_193 = ~(input_a[11] ^ input_a[5]);
  assign popcount36_vanw_core_195 = ~(input_a[14] & input_a[24]);
  assign popcount36_vanw_core_198 = input_a[31] & input_a[32];
  assign popcount36_vanw_core_200 = input_a[25] & input_a[35];
  assign popcount36_vanw_core_201 = input_a[3] & input_a[10];
  assign popcount36_vanw_core_202 = input_a[33] & input_a[34];
  assign popcount36_vanw_core_203 = popcount36_vanw_core_200 | popcount36_vanw_core_202;
  assign popcount36_vanw_core_205 = input_a[35] | input_a[29];
  assign popcount36_vanw_core_206 = input_a[22] & input_a[18];
  assign popcount36_vanw_core_207 = popcount36_vanw_core_198 ^ popcount36_vanw_core_203;
  assign popcount36_vanw_core_208 = popcount36_vanw_core_198 & popcount36_vanw_core_203;
  assign popcount36_vanw_core_209 = popcount36_vanw_core_207 ^ popcount36_vanw_core_206;
  assign popcount36_vanw_core_210 = popcount36_vanw_core_207 & popcount36_vanw_core_206;
  assign popcount36_vanw_core_211 = popcount36_vanw_core_208 | popcount36_vanw_core_210;
  assign popcount36_vanw_core_213 = ~(input_a[2] | input_a[8]);
  assign popcount36_vanw_core_215 = input_a[29] ^ input_a[11];
  assign popcount36_vanw_core_216 = popcount36_vanw_core_192 ^ popcount36_vanw_core_209;
  assign popcount36_vanw_core_217 = popcount36_vanw_core_192 & popcount36_vanw_core_209;
  assign popcount36_vanw_core_222_not = ~input_a[26];
  assign popcount36_vanw_core_223 = popcount36_vanw_core_211 | popcount36_vanw_core_217;
  assign popcount36_vanw_core_224 = input_a[20] & input_a[9];
  assign popcount36_vanw_core_225 = ~input_a[15];
  assign popcount36_vanw_core_227 = ~(input_a[27] ^ input_a[22]);
  assign popcount36_vanw_core_228 = ~(input_a[33] ^ input_a[32]);
  assign popcount36_vanw_core_230 = popcount36_vanw_core_174 | popcount36_vanw_core_216;
  assign popcount36_vanw_core_235 = popcount36_vanw_core_181 ^ popcount36_vanw_core_223;
  assign popcount36_vanw_core_236 = popcount36_vanw_core_181 & popcount36_vanw_core_223;
  assign popcount36_vanw_core_237 = popcount36_vanw_core_235 ^ popcount36_vanw_core_230;
  assign popcount36_vanw_core_238 = popcount36_vanw_core_235 & popcount36_vanw_core_230;
  assign popcount36_vanw_core_239 = popcount36_vanw_core_236 | popcount36_vanw_core_238;
  assign popcount36_vanw_core_241 = ~input_a[6];
  assign popcount36_vanw_core_243 = ~(input_a[19] & input_a[21]);
  assign popcount36_vanw_core_244 = ~(input_a[21] | input_a[12]);
  assign popcount36_vanw_core_245 = ~(input_a[26] | input_a[23]);
  assign popcount36_vanw_core_247 = ~(input_a[25] & input_a[23]);
  assign popcount36_vanw_core_249 = ~(input_a[34] ^ input_a[23]);
  assign popcount36_vanw_core_251 = ~input_a[35];
  assign popcount36_vanw_core_257 = popcount36_vanw_core_131 ^ popcount36_vanw_core_237;
  assign popcount36_vanw_core_258 = popcount36_vanw_core_131 & popcount36_vanw_core_237;
  assign popcount36_vanw_core_259 = popcount36_vanw_core_257 ^ popcount36_vanw_core_126;
  assign popcount36_vanw_core_260 = popcount36_vanw_core_257 & popcount36_vanw_core_126;
  assign popcount36_vanw_core_261 = popcount36_vanw_core_258 | popcount36_vanw_core_260;
  assign popcount36_vanw_core_262 = popcount36_vanw_core_133 ^ popcount36_vanw_core_239;
  assign popcount36_vanw_core_263 = popcount36_vanw_core_133 & popcount36_vanw_core_239;
  assign popcount36_vanw_core_264 = popcount36_vanw_core_262 ^ popcount36_vanw_core_261;
  assign popcount36_vanw_core_265 = popcount36_vanw_core_262 & popcount36_vanw_core_261;
  assign popcount36_vanw_core_266 = popcount36_vanw_core_263 | popcount36_vanw_core_265;
  assign popcount36_vanw_core_267 = ~(input_a[12] ^ input_a[10]);
  assign popcount36_vanw_core_270 = ~(input_a[10] ^ input_a[23]);
  assign popcount36_vanw_core_275 = ~(input_a[26] | input_a[21]);

  assign popcount36_vanw_out[0] = 1'b0;
  assign popcount36_vanw_out[1] = popcount36_vanw_core_124;
  assign popcount36_vanw_out[2] = popcount36_vanw_core_259;
  assign popcount36_vanw_out[3] = popcount36_vanw_core_264;
  assign popcount36_vanw_out[4] = popcount36_vanw_core_266;
  assign popcount36_vanw_out[5] = 1'b0;
endmodule