// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.30917
// WCE=17.0
// EP=0.864166%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_3lws(input [34:0] input_a, output [5:0] popcount35_3lws_out);
  wire popcount35_3lws_core_038;
  wire popcount35_3lws_core_040;
  wire popcount35_3lws_core_042;
  wire popcount35_3lws_core_043;
  wire popcount35_3lws_core_044;
  wire popcount35_3lws_core_045;
  wire popcount35_3lws_core_046_not;
  wire popcount35_3lws_core_048;
  wire popcount35_3lws_core_049;
  wire popcount35_3lws_core_050;
  wire popcount35_3lws_core_055;
  wire popcount35_3lws_core_056;
  wire popcount35_3lws_core_057;
  wire popcount35_3lws_core_058;
  wire popcount35_3lws_core_059;
  wire popcount35_3lws_core_060;
  wire popcount35_3lws_core_063;
  wire popcount35_3lws_core_068;
  wire popcount35_3lws_core_069;
  wire popcount35_3lws_core_070;
  wire popcount35_3lws_core_071;
  wire popcount35_3lws_core_072;
  wire popcount35_3lws_core_074;
  wire popcount35_3lws_core_075;
  wire popcount35_3lws_core_078;
  wire popcount35_3lws_core_079_not;
  wire popcount35_3lws_core_080;
  wire popcount35_3lws_core_082;
  wire popcount35_3lws_core_084;
  wire popcount35_3lws_core_085;
  wire popcount35_3lws_core_087;
  wire popcount35_3lws_core_088;
  wire popcount35_3lws_core_089;
  wire popcount35_3lws_core_091;
  wire popcount35_3lws_core_092;
  wire popcount35_3lws_core_093;
  wire popcount35_3lws_core_094;
  wire popcount35_3lws_core_095;
  wire popcount35_3lws_core_096;
  wire popcount35_3lws_core_098;
  wire popcount35_3lws_core_099;
  wire popcount35_3lws_core_103;
  wire popcount35_3lws_core_104;
  wire popcount35_3lws_core_107;
  wire popcount35_3lws_core_108;
  wire popcount35_3lws_core_111;
  wire popcount35_3lws_core_112;
  wire popcount35_3lws_core_113;
  wire popcount35_3lws_core_115;
  wire popcount35_3lws_core_118;
  wire popcount35_3lws_core_119;
  wire popcount35_3lws_core_120;
  wire popcount35_3lws_core_121;
  wire popcount35_3lws_core_122;
  wire popcount35_3lws_core_123;
  wire popcount35_3lws_core_124;
  wire popcount35_3lws_core_125;
  wire popcount35_3lws_core_126;
  wire popcount35_3lws_core_127;
  wire popcount35_3lws_core_128;
  wire popcount35_3lws_core_129;
  wire popcount35_3lws_core_130;
  wire popcount35_3lws_core_131;
  wire popcount35_3lws_core_132;
  wire popcount35_3lws_core_133;
  wire popcount35_3lws_core_134;
  wire popcount35_3lws_core_135;
  wire popcount35_3lws_core_138;
  wire popcount35_3lws_core_139;
  wire popcount35_3lws_core_140;
  wire popcount35_3lws_core_144;
  wire popcount35_3lws_core_146;
  wire popcount35_3lws_core_147;
  wire popcount35_3lws_core_150;
  wire popcount35_3lws_core_151;
  wire popcount35_3lws_core_154;
  wire popcount35_3lws_core_155;
  wire popcount35_3lws_core_157;
  wire popcount35_3lws_core_158;
  wire popcount35_3lws_core_159;
  wire popcount35_3lws_core_160;
  wire popcount35_3lws_core_161;
  wire popcount35_3lws_core_168;
  wire popcount35_3lws_core_169;
  wire popcount35_3lws_core_170;
  wire popcount35_3lws_core_172;
  wire popcount35_3lws_core_173;
  wire popcount35_3lws_core_175;
  wire popcount35_3lws_core_176;
  wire popcount35_3lws_core_179;
  wire popcount35_3lws_core_181;
  wire popcount35_3lws_core_183;
  wire popcount35_3lws_core_184;
  wire popcount35_3lws_core_185;
  wire popcount35_3lws_core_186;
  wire popcount35_3lws_core_187;
  wire popcount35_3lws_core_188;
  wire popcount35_3lws_core_190;
  wire popcount35_3lws_core_192;
  wire popcount35_3lws_core_193;
  wire popcount35_3lws_core_195;
  wire popcount35_3lws_core_196;
  wire popcount35_3lws_core_197;
  wire popcount35_3lws_core_199;
  wire popcount35_3lws_core_200;
  wire popcount35_3lws_core_202;
  wire popcount35_3lws_core_203;
  wire popcount35_3lws_core_205;
  wire popcount35_3lws_core_208;
  wire popcount35_3lws_core_209;
  wire popcount35_3lws_core_212;
  wire popcount35_3lws_core_213;
  wire popcount35_3lws_core_214;
  wire popcount35_3lws_core_215;
  wire popcount35_3lws_core_216;
  wire popcount35_3lws_core_217;
  wire popcount35_3lws_core_218;
  wire popcount35_3lws_core_219;
  wire popcount35_3lws_core_222;
  wire popcount35_3lws_core_223;
  wire popcount35_3lws_core_224;
  wire popcount35_3lws_core_227;
  wire popcount35_3lws_core_228;
  wire popcount35_3lws_core_229;
  wire popcount35_3lws_core_230;
  wire popcount35_3lws_core_233;
  wire popcount35_3lws_core_234;
  wire popcount35_3lws_core_235;
  wire popcount35_3lws_core_236;
  wire popcount35_3lws_core_237;
  wire popcount35_3lws_core_238;
  wire popcount35_3lws_core_239;
  wire popcount35_3lws_core_240;
  wire popcount35_3lws_core_241;
  wire popcount35_3lws_core_242;
  wire popcount35_3lws_core_243;
  wire popcount35_3lws_core_246_not;
  wire popcount35_3lws_core_247;
  wire popcount35_3lws_core_249;
  wire popcount35_3lws_core_251;
  wire popcount35_3lws_core_253;
  wire popcount35_3lws_core_256;
  wire popcount35_3lws_core_257;
  wire popcount35_3lws_core_259;
  wire popcount35_3lws_core_261;
  wire popcount35_3lws_core_262;
  wire popcount35_3lws_core_263;
  wire popcount35_3lws_core_264;

  assign popcount35_3lws_core_038 = input_a[19] | input_a[27];
  assign popcount35_3lws_core_040 = input_a[0] ^ input_a[8];
  assign popcount35_3lws_core_042 = ~(input_a[21] & input_a[33]);
  assign popcount35_3lws_core_043 = input_a[18] ^ input_a[18];
  assign popcount35_3lws_core_044 = input_a[21] & input_a[15];
  assign popcount35_3lws_core_045 = input_a[26] & input_a[16];
  assign popcount35_3lws_core_046_not = ~input_a[24];
  assign popcount35_3lws_core_048 = input_a[3] | input_a[18];
  assign popcount35_3lws_core_049 = ~(input_a[27] & input_a[19]);
  assign popcount35_3lws_core_050 = ~(input_a[31] | input_a[10]);
  assign popcount35_3lws_core_055 = ~(input_a[28] & input_a[28]);
  assign popcount35_3lws_core_056 = input_a[21] | input_a[33];
  assign popcount35_3lws_core_057 = ~(input_a[3] ^ input_a[6]);
  assign popcount35_3lws_core_058 = ~(input_a[29] & input_a[6]);
  assign popcount35_3lws_core_059 = ~(input_a[10] ^ input_a[2]);
  assign popcount35_3lws_core_060 = ~input_a[2];
  assign popcount35_3lws_core_063 = ~input_a[34];
  assign popcount35_3lws_core_068 = ~(input_a[15] & input_a[5]);
  assign popcount35_3lws_core_069 = ~(input_a[24] ^ input_a[2]);
  assign popcount35_3lws_core_070 = ~(input_a[34] ^ input_a[24]);
  assign popcount35_3lws_core_071 = input_a[13] | input_a[18];
  assign popcount35_3lws_core_072 = ~(input_a[14] | input_a[33]);
  assign popcount35_3lws_core_074 = input_a[14] | input_a[30];
  assign popcount35_3lws_core_075 = ~input_a[17];
  assign popcount35_3lws_core_078 = ~(input_a[27] | input_a[3]);
  assign popcount35_3lws_core_079_not = ~input_a[22];
  assign popcount35_3lws_core_080 = input_a[2] | input_a[6];
  assign popcount35_3lws_core_082 = input_a[21] | input_a[24];
  assign popcount35_3lws_core_084 = input_a[17] & input_a[25];
  assign popcount35_3lws_core_085 = input_a[2] | input_a[23];
  assign popcount35_3lws_core_087 = input_a[13] ^ input_a[34];
  assign popcount35_3lws_core_088 = ~input_a[25];
  assign popcount35_3lws_core_089 = input_a[14] & input_a[12];
  assign popcount35_3lws_core_091 = ~(input_a[28] | input_a[14]);
  assign popcount35_3lws_core_092 = ~(input_a[5] ^ input_a[18]);
  assign popcount35_3lws_core_093 = ~(input_a[1] | input_a[29]);
  assign popcount35_3lws_core_094 = input_a[34] & input_a[33];
  assign popcount35_3lws_core_095 = ~(input_a[22] & input_a[17]);
  assign popcount35_3lws_core_096 = input_a[18] ^ input_a[7];
  assign popcount35_3lws_core_098 = ~(input_a[0] | input_a[29]);
  assign popcount35_3lws_core_099 = ~(input_a[34] & input_a[17]);
  assign popcount35_3lws_core_103 = input_a[26] | input_a[4];
  assign popcount35_3lws_core_104 = input_a[26] & input_a[1];
  assign popcount35_3lws_core_107 = ~input_a[26];
  assign popcount35_3lws_core_108 = input_a[20] | input_a[16];
  assign popcount35_3lws_core_111 = input_a[16] | input_a[12];
  assign popcount35_3lws_core_112 = input_a[16] | input_a[21];
  assign popcount35_3lws_core_113 = input_a[5] & input_a[6];
  assign popcount35_3lws_core_115 = input_a[23] | input_a[17];
  assign popcount35_3lws_core_118 = ~(input_a[11] ^ input_a[14]);
  assign popcount35_3lws_core_119 = input_a[26] ^ input_a[15];
  assign popcount35_3lws_core_120 = input_a[14] | input_a[4];
  assign popcount35_3lws_core_121 = ~input_a[28];
  assign popcount35_3lws_core_122 = input_a[33] & input_a[25];
  assign popcount35_3lws_core_123 = input_a[17] ^ input_a[8];
  assign popcount35_3lws_core_124 = input_a[10] ^ input_a[11];
  assign popcount35_3lws_core_125 = input_a[24] ^ input_a[9];
  assign popcount35_3lws_core_126 = input_a[16] & input_a[11];
  assign popcount35_3lws_core_127 = ~(input_a[7] & input_a[2]);
  assign popcount35_3lws_core_128 = ~input_a[0];
  assign popcount35_3lws_core_129 = input_a[3] ^ input_a[19];
  assign popcount35_3lws_core_130 = input_a[34] | input_a[12];
  assign popcount35_3lws_core_131 = input_a[12] | input_a[33];
  assign popcount35_3lws_core_132 = ~input_a[32];
  assign popcount35_3lws_core_133 = ~(input_a[21] | input_a[26]);
  assign popcount35_3lws_core_134 = input_a[30] & input_a[25];
  assign popcount35_3lws_core_135 = input_a[7] ^ input_a[32];
  assign popcount35_3lws_core_138 = input_a[30] & input_a[33];
  assign popcount35_3lws_core_139 = input_a[13] ^ input_a[10];
  assign popcount35_3lws_core_140 = ~(input_a[32] | input_a[11]);
  assign popcount35_3lws_core_144 = input_a[20] | input_a[24];
  assign popcount35_3lws_core_146 = ~input_a[0];
  assign popcount35_3lws_core_147 = input_a[7] ^ input_a[12];
  assign popcount35_3lws_core_150 = ~(input_a[6] & input_a[30]);
  assign popcount35_3lws_core_151 = input_a[10] | input_a[19];
  assign popcount35_3lws_core_154 = ~(input_a[5] ^ input_a[13]);
  assign popcount35_3lws_core_155 = input_a[18] & input_a[19];
  assign popcount35_3lws_core_157 = input_a[25] | input_a[27];
  assign popcount35_3lws_core_158 = input_a[4] | input_a[7];
  assign popcount35_3lws_core_159 = ~input_a[19];
  assign popcount35_3lws_core_160 = ~input_a[17];
  assign popcount35_3lws_core_161 = input_a[6] & input_a[18];
  assign popcount35_3lws_core_168 = ~(input_a[18] ^ input_a[22]);
  assign popcount35_3lws_core_169 = ~(input_a[5] | input_a[17]);
  assign popcount35_3lws_core_170 = ~(input_a[17] | input_a[22]);
  assign popcount35_3lws_core_172 = ~(input_a[30] ^ input_a[16]);
  assign popcount35_3lws_core_173 = input_a[2] & input_a[12];
  assign popcount35_3lws_core_175 = input_a[17] | input_a[31];
  assign popcount35_3lws_core_176 = ~(input_a[24] | input_a[28]);
  assign popcount35_3lws_core_179 = ~(input_a[8] | input_a[5]);
  assign popcount35_3lws_core_181 = ~input_a[10];
  assign popcount35_3lws_core_183 = input_a[27] & input_a[34];
  assign popcount35_3lws_core_184 = ~(input_a[8] & input_a[30]);
  assign popcount35_3lws_core_185 = ~(input_a[18] & input_a[4]);
  assign popcount35_3lws_core_186 = ~(input_a[30] ^ input_a[4]);
  assign popcount35_3lws_core_187 = ~(input_a[30] | input_a[7]);
  assign popcount35_3lws_core_188 = ~input_a[13];
  assign popcount35_3lws_core_190 = input_a[30] ^ input_a[8];
  assign popcount35_3lws_core_192 = ~(input_a[14] ^ input_a[10]);
  assign popcount35_3lws_core_193 = input_a[17] ^ input_a[30];
  assign popcount35_3lws_core_195 = input_a[28] & input_a[34];
  assign popcount35_3lws_core_196 = ~(input_a[25] & input_a[5]);
  assign popcount35_3lws_core_197 = input_a[29] & input_a[28];
  assign popcount35_3lws_core_199 = ~(input_a[13] & input_a[25]);
  assign popcount35_3lws_core_200 = ~(input_a[6] & input_a[34]);
  assign popcount35_3lws_core_202 = ~input_a[21];
  assign popcount35_3lws_core_203 = ~(input_a[22] | input_a[32]);
  assign popcount35_3lws_core_205 = input_a[22] | input_a[22];
  assign popcount35_3lws_core_208 = ~(input_a[12] ^ input_a[7]);
  assign popcount35_3lws_core_209 = ~input_a[2];
  assign popcount35_3lws_core_212 = input_a[5] ^ input_a[5];
  assign popcount35_3lws_core_213 = input_a[29] ^ input_a[24];
  assign popcount35_3lws_core_214 = input_a[21] ^ input_a[31];
  assign popcount35_3lws_core_215 = input_a[14] | input_a[7];
  assign popcount35_3lws_core_216 = input_a[5] | input_a[20];
  assign popcount35_3lws_core_217 = input_a[11] & input_a[4];
  assign popcount35_3lws_core_218 = input_a[24] & input_a[3];
  assign popcount35_3lws_core_219 = ~input_a[0];
  assign popcount35_3lws_core_222 = input_a[3] & input_a[12];
  assign popcount35_3lws_core_223 = ~(input_a[17] ^ input_a[25]);
  assign popcount35_3lws_core_224 = ~(input_a[7] ^ input_a[30]);
  assign popcount35_3lws_core_227 = ~input_a[23];
  assign popcount35_3lws_core_228 = ~(input_a[19] & input_a[10]);
  assign popcount35_3lws_core_229 = ~(input_a[20] & input_a[15]);
  assign popcount35_3lws_core_230 = input_a[31] & input_a[9];
  assign popcount35_3lws_core_233 = ~(input_a[1] & input_a[10]);
  assign popcount35_3lws_core_234 = ~(input_a[5] & input_a[18]);
  assign popcount35_3lws_core_235 = ~(input_a[1] ^ input_a[34]);
  assign popcount35_3lws_core_236 = input_a[12] ^ input_a[22];
  assign popcount35_3lws_core_237 = input_a[10] | input_a[27];
  assign popcount35_3lws_core_238 = input_a[10] ^ input_a[15];
  assign popcount35_3lws_core_239 = ~(input_a[8] & input_a[5]);
  assign popcount35_3lws_core_240 = input_a[28] & input_a[2];
  assign popcount35_3lws_core_241 = ~input_a[31];
  assign popcount35_3lws_core_242 = input_a[8] ^ input_a[15];
  assign popcount35_3lws_core_243 = ~(input_a[3] ^ input_a[11]);
  assign popcount35_3lws_core_246_not = ~input_a[5];
  assign popcount35_3lws_core_247 = ~(input_a[6] & input_a[7]);
  assign popcount35_3lws_core_249 = ~(input_a[15] & input_a[23]);
  assign popcount35_3lws_core_251 = ~input_a[33];
  assign popcount35_3lws_core_253 = ~(input_a[14] ^ input_a[10]);
  assign popcount35_3lws_core_256 = ~input_a[29];
  assign popcount35_3lws_core_257 = ~(input_a[10] ^ input_a[25]);
  assign popcount35_3lws_core_259 = ~(input_a[26] ^ input_a[29]);
  assign popcount35_3lws_core_261 = input_a[19] & input_a[1];
  assign popcount35_3lws_core_262 = ~(input_a[12] ^ input_a[32]);
  assign popcount35_3lws_core_263 = input_a[3] | input_a[12];
  assign popcount35_3lws_core_264 = ~(input_a[17] | input_a[28]);

  assign popcount35_3lws_out[0] = input_a[13];
  assign popcount35_3lws_out[1] = input_a[30];
  assign popcount35_3lws_out[2] = 1'b0;
  assign popcount35_3lws_out[3] = 1'b0;
  assign popcount35_3lws_out[4] = 1'b1;
  assign popcount35_3lws_out[5] = 1'b0;
endmodule