// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.19788
// WCE=20.0
// EP=0.907496%
// Printed PDK parameters:
//  Area=1638800.0
//  Delay=3352434.5
//  Power=75843.0

module popcount40_2dxt(input [39:0] input_a, output [5:0] popcount40_2dxt_out);
  wire popcount40_2dxt_core_042;
  wire popcount40_2dxt_core_047;
  wire popcount40_2dxt_core_048;
  wire popcount40_2dxt_core_049;
  wire popcount40_2dxt_core_050;
  wire popcount40_2dxt_core_051;
  wire popcount40_2dxt_core_053;
  wire popcount40_2dxt_core_054;
  wire popcount40_2dxt_core_056;
  wire popcount40_2dxt_core_057;
  wire popcount40_2dxt_core_059;
  wire popcount40_2dxt_core_061;
  wire popcount40_2dxt_core_062;
  wire popcount40_2dxt_core_063;
  wire popcount40_2dxt_core_064;
  wire popcount40_2dxt_core_065;
  wire popcount40_2dxt_core_068;
  wire popcount40_2dxt_core_071;
  wire popcount40_2dxt_core_072;
  wire popcount40_2dxt_core_074;
  wire popcount40_2dxt_core_075;
  wire popcount40_2dxt_core_076;
  wire popcount40_2dxt_core_077;
  wire popcount40_2dxt_core_080;
  wire popcount40_2dxt_core_081;
  wire popcount40_2dxt_core_083;
  wire popcount40_2dxt_core_086;
  wire popcount40_2dxt_core_088;
  wire popcount40_2dxt_core_089;
  wire popcount40_2dxt_core_091;
  wire popcount40_2dxt_core_092;
  wire popcount40_2dxt_core_093;
  wire popcount40_2dxt_core_095;
  wire popcount40_2dxt_core_096;
  wire popcount40_2dxt_core_097;
  wire popcount40_2dxt_core_098;
  wire popcount40_2dxt_core_099;
  wire popcount40_2dxt_core_100;
  wire popcount40_2dxt_core_101;
  wire popcount40_2dxt_core_102;
  wire popcount40_2dxt_core_103;
  wire popcount40_2dxt_core_104;
  wire popcount40_2dxt_core_105;
  wire popcount40_2dxt_core_106;
  wire popcount40_2dxt_core_107;
  wire popcount40_2dxt_core_110;
  wire popcount40_2dxt_core_111;
  wire popcount40_2dxt_core_112;
  wire popcount40_2dxt_core_115;
  wire popcount40_2dxt_core_117;
  wire popcount40_2dxt_core_118;
  wire popcount40_2dxt_core_119;
  wire popcount40_2dxt_core_120;
  wire popcount40_2dxt_core_125;
  wire popcount40_2dxt_core_126;
  wire popcount40_2dxt_core_127;
  wire popcount40_2dxt_core_128;
  wire popcount40_2dxt_core_130;
  wire popcount40_2dxt_core_131;
  wire popcount40_2dxt_core_132;
  wire popcount40_2dxt_core_134;
  wire popcount40_2dxt_core_136;
  wire popcount40_2dxt_core_137;
  wire popcount40_2dxt_core_138;
  wire popcount40_2dxt_core_139;
  wire popcount40_2dxt_core_140;
  wire popcount40_2dxt_core_143_not;
  wire popcount40_2dxt_core_146;
  wire popcount40_2dxt_core_147;
  wire popcount40_2dxt_core_148;
  wire popcount40_2dxt_core_150;
  wire popcount40_2dxt_core_151;
  wire popcount40_2dxt_core_155;
  wire popcount40_2dxt_core_156;
  wire popcount40_2dxt_core_158;
  wire popcount40_2dxt_core_159;
  wire popcount40_2dxt_core_161;
  wire popcount40_2dxt_core_162;
  wire popcount40_2dxt_core_164;
  wire popcount40_2dxt_core_165;
  wire popcount40_2dxt_core_170;
  wire popcount40_2dxt_core_171;
  wire popcount40_2dxt_core_173;
  wire popcount40_2dxt_core_174;
  wire popcount40_2dxt_core_177;
  wire popcount40_2dxt_core_178;
  wire popcount40_2dxt_core_179;
  wire popcount40_2dxt_core_180;
  wire popcount40_2dxt_core_181;
  wire popcount40_2dxt_core_182;
  wire popcount40_2dxt_core_183;
  wire popcount40_2dxt_core_187;
  wire popcount40_2dxt_core_188;
  wire popcount40_2dxt_core_190;
  wire popcount40_2dxt_core_191;
  wire popcount40_2dxt_core_192;
  wire popcount40_2dxt_core_193;
  wire popcount40_2dxt_core_194;
  wire popcount40_2dxt_core_197;
  wire popcount40_2dxt_core_199;
  wire popcount40_2dxt_core_203;
  wire popcount40_2dxt_core_204;
  wire popcount40_2dxt_core_205;
  wire popcount40_2dxt_core_206;
  wire popcount40_2dxt_core_207;
  wire popcount40_2dxt_core_208;
  wire popcount40_2dxt_core_211;
  wire popcount40_2dxt_core_212;
  wire popcount40_2dxt_core_213;
  wire popcount40_2dxt_core_214;
  wire popcount40_2dxt_core_215;
  wire popcount40_2dxt_core_216;
  wire popcount40_2dxt_core_217;
  wire popcount40_2dxt_core_220;
  wire popcount40_2dxt_core_222;
  wire popcount40_2dxt_core_223;
  wire popcount40_2dxt_core_227;
  wire popcount40_2dxt_core_229_not;
  wire popcount40_2dxt_core_230;
  wire popcount40_2dxt_core_232;
  wire popcount40_2dxt_core_234;
  wire popcount40_2dxt_core_236;
  wire popcount40_2dxt_core_237;
  wire popcount40_2dxt_core_238;
  wire popcount40_2dxt_core_239;
  wire popcount40_2dxt_core_240;
  wire popcount40_2dxt_core_242;
  wire popcount40_2dxt_core_244_not;
  wire popcount40_2dxt_core_245;
  wire popcount40_2dxt_core_246;
  wire popcount40_2dxt_core_247;
  wire popcount40_2dxt_core_248;
  wire popcount40_2dxt_core_251;
  wire popcount40_2dxt_core_252;
  wire popcount40_2dxt_core_254;
  wire popcount40_2dxt_core_255;
  wire popcount40_2dxt_core_256;
  wire popcount40_2dxt_core_258;
  wire popcount40_2dxt_core_259;
  wire popcount40_2dxt_core_261;
  wire popcount40_2dxt_core_262;
  wire popcount40_2dxt_core_266;
  wire popcount40_2dxt_core_270;
  wire popcount40_2dxt_core_271;
  wire popcount40_2dxt_core_272;
  wire popcount40_2dxt_core_273;
  wire popcount40_2dxt_core_274;
  wire popcount40_2dxt_core_276;
  wire popcount40_2dxt_core_278;
  wire popcount40_2dxt_core_280;
  wire popcount40_2dxt_core_281;
  wire popcount40_2dxt_core_282;
  wire popcount40_2dxt_core_283;
  wire popcount40_2dxt_core_284;
  wire popcount40_2dxt_core_285;
  wire popcount40_2dxt_core_288;
  wire popcount40_2dxt_core_290;
  wire popcount40_2dxt_core_291;
  wire popcount40_2dxt_core_292;
  wire popcount40_2dxt_core_294;
  wire popcount40_2dxt_core_296;
  wire popcount40_2dxt_core_298;
  wire popcount40_2dxt_core_299;
  wire popcount40_2dxt_core_300;
  wire popcount40_2dxt_core_301;
  wire popcount40_2dxt_core_302;
  wire popcount40_2dxt_core_303;
  wire popcount40_2dxt_core_306;
  wire popcount40_2dxt_core_307;
  wire popcount40_2dxt_core_308;
  wire popcount40_2dxt_core_312;
  wire popcount40_2dxt_core_313;
  wire popcount40_2dxt_core_314;
  wire popcount40_2dxt_core_316;

  assign popcount40_2dxt_core_042 = ~(input_a[24] ^ input_a[4]);
  assign popcount40_2dxt_core_047 = ~input_a[11];
  assign popcount40_2dxt_core_048 = input_a[5] | input_a[21];
  assign popcount40_2dxt_core_049 = input_a[32] & input_a[25];
  assign popcount40_2dxt_core_050 = ~(input_a[0] | input_a[17]);
  assign popcount40_2dxt_core_051 = ~(input_a[28] ^ input_a[36]);
  assign popcount40_2dxt_core_053 = input_a[39] | input_a[34];
  assign popcount40_2dxt_core_054 = ~input_a[22];
  assign popcount40_2dxt_core_056 = ~(input_a[18] | input_a[13]);
  assign popcount40_2dxt_core_057 = input_a[25] & input_a[27];
  assign popcount40_2dxt_core_059 = ~(input_a[33] & input_a[35]);
  assign popcount40_2dxt_core_061 = ~(input_a[5] ^ input_a[0]);
  assign popcount40_2dxt_core_062 = input_a[8] | input_a[6];
  assign popcount40_2dxt_core_063 = ~(input_a[39] ^ input_a[12]);
  assign popcount40_2dxt_core_064 = input_a[20] | input_a[35];
  assign popcount40_2dxt_core_065 = ~(input_a[27] & input_a[22]);
  assign popcount40_2dxt_core_068 = input_a[21] ^ input_a[2];
  assign popcount40_2dxt_core_071 = ~(input_a[4] | input_a[21]);
  assign popcount40_2dxt_core_072 = ~(input_a[1] ^ input_a[30]);
  assign popcount40_2dxt_core_074 = input_a[20] & input_a[30];
  assign popcount40_2dxt_core_075 = ~input_a[10];
  assign popcount40_2dxt_core_076 = input_a[1] | input_a[2];
  assign popcount40_2dxt_core_077 = input_a[35] ^ input_a[10];
  assign popcount40_2dxt_core_080 = input_a[37] & input_a[38];
  assign popcount40_2dxt_core_081 = ~input_a[33];
  assign popcount40_2dxt_core_083 = input_a[23] | input_a[14];
  assign popcount40_2dxt_core_086 = input_a[4] ^ input_a[13];
  assign popcount40_2dxt_core_088 = ~(input_a[14] & input_a[1]);
  assign popcount40_2dxt_core_089 = input_a[31] ^ input_a[8];
  assign popcount40_2dxt_core_091 = ~input_a[28];
  assign popcount40_2dxt_core_092 = ~(input_a[2] & input_a[0]);
  assign popcount40_2dxt_core_093 = ~input_a[27];
  assign popcount40_2dxt_core_095 = ~(input_a[30] ^ input_a[27]);
  assign popcount40_2dxt_core_096 = ~(input_a[6] | input_a[21]);
  assign popcount40_2dxt_core_097 = ~(input_a[5] ^ input_a[20]);
  assign popcount40_2dxt_core_098 = input_a[5] & input_a[18];
  assign popcount40_2dxt_core_099 = input_a[28] | input_a[24];
  assign popcount40_2dxt_core_100 = input_a[5] ^ input_a[38];
  assign popcount40_2dxt_core_101 = ~(input_a[38] & input_a[17]);
  assign popcount40_2dxt_core_102 = input_a[10] & input_a[8];
  assign popcount40_2dxt_core_103 = ~(input_a[39] & input_a[33]);
  assign popcount40_2dxt_core_104 = ~(input_a[19] | input_a[28]);
  assign popcount40_2dxt_core_105 = input_a[34] | input_a[0];
  assign popcount40_2dxt_core_106 = input_a[2] ^ input_a[11];
  assign popcount40_2dxt_core_107 = ~(input_a[20] ^ input_a[31]);
  assign popcount40_2dxt_core_110 = ~(input_a[24] ^ input_a[10]);
  assign popcount40_2dxt_core_111 = input_a[14] | input_a[19];
  assign popcount40_2dxt_core_112 = input_a[15] | input_a[5];
  assign popcount40_2dxt_core_115 = input_a[22] & input_a[14];
  assign popcount40_2dxt_core_117 = input_a[20] & input_a[34];
  assign popcount40_2dxt_core_118 = ~(input_a[19] | input_a[29]);
  assign popcount40_2dxt_core_119 = ~(input_a[4] | input_a[37]);
  assign popcount40_2dxt_core_120 = input_a[35] ^ input_a[38];
  assign popcount40_2dxt_core_125 = ~(input_a[33] | input_a[16]);
  assign popcount40_2dxt_core_126 = ~input_a[30];
  assign popcount40_2dxt_core_127 = input_a[26] | input_a[17];
  assign popcount40_2dxt_core_128 = input_a[35] & input_a[1];
  assign popcount40_2dxt_core_130 = ~(input_a[24] | input_a[31]);
  assign popcount40_2dxt_core_131 = input_a[1] & input_a[30];
  assign popcount40_2dxt_core_132 = ~(input_a[3] | input_a[5]);
  assign popcount40_2dxt_core_134 = ~(input_a[33] ^ input_a[24]);
  assign popcount40_2dxt_core_136 = ~input_a[16];
  assign popcount40_2dxt_core_137 = ~(input_a[7] ^ input_a[4]);
  assign popcount40_2dxt_core_138 = ~input_a[4];
  assign popcount40_2dxt_core_139 = ~(input_a[15] ^ input_a[22]);
  assign popcount40_2dxt_core_140 = ~(input_a[36] & input_a[32]);
  assign popcount40_2dxt_core_143_not = ~input_a[35];
  assign popcount40_2dxt_core_146 = ~(input_a[16] | input_a[30]);
  assign popcount40_2dxt_core_147 = input_a[17] & input_a[36];
  assign popcount40_2dxt_core_148 = ~(input_a[12] | input_a[11]);
  assign popcount40_2dxt_core_150 = ~(input_a[14] | input_a[27]);
  assign popcount40_2dxt_core_151 = ~input_a[4];
  assign popcount40_2dxt_core_155 = ~(input_a[28] ^ input_a[6]);
  assign popcount40_2dxt_core_156 = input_a[17] | input_a[23];
  assign popcount40_2dxt_core_158 = ~(input_a[31] ^ input_a[26]);
  assign popcount40_2dxt_core_159 = input_a[17] ^ input_a[10];
  assign popcount40_2dxt_core_161 = ~input_a[35];
  assign popcount40_2dxt_core_162 = ~(input_a[25] | input_a[37]);
  assign popcount40_2dxt_core_164 = ~(input_a[30] ^ input_a[8]);
  assign popcount40_2dxt_core_165 = input_a[0] & input_a[32];
  assign popcount40_2dxt_core_170 = ~input_a[1];
  assign popcount40_2dxt_core_171 = ~(input_a[0] & input_a[2]);
  assign popcount40_2dxt_core_173 = input_a[0] | input_a[1];
  assign popcount40_2dxt_core_174 = input_a[15] | input_a[9];
  assign popcount40_2dxt_core_177 = input_a[39] & input_a[1];
  assign popcount40_2dxt_core_178 = ~(input_a[16] | input_a[14]);
  assign popcount40_2dxt_core_179 = input_a[28] & input_a[37];
  assign popcount40_2dxt_core_180 = popcount40_2dxt_core_177 | popcount40_2dxt_core_179;
  assign popcount40_2dxt_core_181 = input_a[30] & input_a[24];
  assign popcount40_2dxt_core_182 = ~input_a[2];
  assign popcount40_2dxt_core_183 = ~(input_a[28] ^ input_a[0]);
  assign popcount40_2dxt_core_187 = ~(input_a[11] | input_a[26]);
  assign popcount40_2dxt_core_188 = ~(input_a[3] ^ input_a[22]);
  assign popcount40_2dxt_core_190 = ~(input_a[29] | input_a[8]);
  assign popcount40_2dxt_core_191 = ~(input_a[15] ^ input_a[17]);
  assign popcount40_2dxt_core_192 = input_a[2] ^ input_a[8];
  assign popcount40_2dxt_core_193 = ~(input_a[6] | input_a[27]);
  assign popcount40_2dxt_core_194 = ~(input_a[25] ^ input_a[13]);
  assign popcount40_2dxt_core_197 = ~(input_a[27] | input_a[19]);
  assign popcount40_2dxt_core_199 = input_a[10] ^ input_a[29];
  assign popcount40_2dxt_core_203 = input_a[26] ^ input_a[19];
  assign popcount40_2dxt_core_204 = input_a[11] & input_a[13];
  assign popcount40_2dxt_core_205 = ~(input_a[35] | input_a[17]);
  assign popcount40_2dxt_core_206 = input_a[20] ^ input_a[1];
  assign popcount40_2dxt_core_207 = input_a[0] & input_a[30];
  assign popcount40_2dxt_core_208 = ~(input_a[0] & input_a[22]);
  assign popcount40_2dxt_core_211 = ~input_a[15];
  assign popcount40_2dxt_core_212 = ~input_a[32];
  assign popcount40_2dxt_core_213 = input_a[2] ^ input_a[27];
  assign popcount40_2dxt_core_214 = ~(input_a[12] | input_a[7]);
  assign popcount40_2dxt_core_215 = input_a[32] | input_a[13];
  assign popcount40_2dxt_core_216 = ~(input_a[21] ^ input_a[15]);
  assign popcount40_2dxt_core_217 = ~input_a[39];
  assign popcount40_2dxt_core_220 = ~(input_a[37] ^ input_a[26]);
  assign popcount40_2dxt_core_222 = input_a[1] ^ input_a[13];
  assign popcount40_2dxt_core_223 = ~input_a[18];
  assign popcount40_2dxt_core_227 = ~(input_a[33] & input_a[20]);
  assign popcount40_2dxt_core_229_not = ~input_a[18];
  assign popcount40_2dxt_core_230 = ~(input_a[3] & input_a[29]);
  assign popcount40_2dxt_core_232 = input_a[17] & input_a[15];
  assign popcount40_2dxt_core_234 = ~(input_a[20] & input_a[7]);
  assign popcount40_2dxt_core_236 = ~input_a[21];
  assign popcount40_2dxt_core_237 = ~(input_a[39] & input_a[3]);
  assign popcount40_2dxt_core_238 = ~input_a[30];
  assign popcount40_2dxt_core_239 = ~input_a[16];
  assign popcount40_2dxt_core_240 = ~(input_a[22] | input_a[23]);
  assign popcount40_2dxt_core_242 = input_a[17] ^ input_a[14];
  assign popcount40_2dxt_core_244_not = ~input_a[7];
  assign popcount40_2dxt_core_245 = ~(input_a[22] | input_a[7]);
  assign popcount40_2dxt_core_246 = ~(input_a[16] | input_a[33]);
  assign popcount40_2dxt_core_247 = input_a[2] & input_a[22];
  assign popcount40_2dxt_core_248 = input_a[8] ^ input_a[35];
  assign popcount40_2dxt_core_251 = ~(input_a[19] | input_a[18]);
  assign popcount40_2dxt_core_252 = ~input_a[20];
  assign popcount40_2dxt_core_254 = input_a[35] ^ input_a[36];
  assign popcount40_2dxt_core_255 = ~(input_a[11] | input_a[13]);
  assign popcount40_2dxt_core_256 = input_a[39] ^ input_a[18];
  assign popcount40_2dxt_core_258 = ~(input_a[32] & input_a[13]);
  assign popcount40_2dxt_core_259 = input_a[7] | input_a[14];
  assign popcount40_2dxt_core_261 = input_a[11] ^ input_a[1];
  assign popcount40_2dxt_core_262 = input_a[8] ^ input_a[19];
  assign popcount40_2dxt_core_266 = ~(input_a[16] & input_a[17]);
  assign popcount40_2dxt_core_270 = ~(input_a[12] & input_a[20]);
  assign popcount40_2dxt_core_271 = input_a[20] & input_a[11];
  assign popcount40_2dxt_core_272 = ~(input_a[1] ^ input_a[4]);
  assign popcount40_2dxt_core_273 = ~(input_a[4] ^ input_a[12]);
  assign popcount40_2dxt_core_274 = input_a[29] & input_a[21];
  assign popcount40_2dxt_core_276 = input_a[24] ^ input_a[15];
  assign popcount40_2dxt_core_278 = input_a[27] | input_a[37];
  assign popcount40_2dxt_core_280 = ~input_a[28];
  assign popcount40_2dxt_core_281 = ~(input_a[16] & input_a[13]);
  assign popcount40_2dxt_core_282 = input_a[13] ^ input_a[15];
  assign popcount40_2dxt_core_283 = input_a[13] & input_a[17];
  assign popcount40_2dxt_core_284 = ~(input_a[8] & input_a[23]);
  assign popcount40_2dxt_core_285 = ~(input_a[31] ^ input_a[34]);
  assign popcount40_2dxt_core_288 = input_a[12] ^ input_a[2];
  assign popcount40_2dxt_core_290 = ~input_a[16];
  assign popcount40_2dxt_core_291 = input_a[33] & input_a[35];
  assign popcount40_2dxt_core_292 = input_a[22] & input_a[28];
  assign popcount40_2dxt_core_294 = ~(input_a[20] ^ input_a[0]);
  assign popcount40_2dxt_core_296 = input_a[31] & input_a[9];
  assign popcount40_2dxt_core_298 = ~(input_a[11] & input_a[18]);
  assign popcount40_2dxt_core_299 = input_a[27] ^ input_a[31];
  assign popcount40_2dxt_core_300 = popcount40_2dxt_core_274 & popcount40_2dxt_core_296;
  assign popcount40_2dxt_core_301 = input_a[25] | input_a[0];
  assign popcount40_2dxt_core_302 = input_a[28] ^ input_a[11];
  assign popcount40_2dxt_core_303 = ~input_a[28];
  assign popcount40_2dxt_core_306 = input_a[29] | input_a[4];
  assign popcount40_2dxt_core_307 = input_a[4] ^ input_a[31];
  assign popcount40_2dxt_core_308 = ~(input_a[9] & input_a[21]);
  assign popcount40_2dxt_core_312 = input_a[2] ^ input_a[3];
  assign popcount40_2dxt_core_313 = ~(input_a[14] | input_a[1]);
  assign popcount40_2dxt_core_314 = input_a[0] & input_a[25];
  assign popcount40_2dxt_core_316 = ~(input_a[28] ^ input_a[32]);

  assign popcount40_2dxt_out[0] = input_a[0];
  assign popcount40_2dxt_out[1] = popcount40_2dxt_core_180;
  assign popcount40_2dxt_out[2] = 1'b0;
  assign popcount40_2dxt_out[3] = popcount40_2dxt_core_300;
  assign popcount40_2dxt_out[4] = 1'b1;
  assign popcount40_2dxt_out[5] = 1'b0;
endmodule