// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.82588
// WCE=30.0
// EP=0.96744%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_7qyk(input [32:0] input_a, output [5:0] popcount33_7qyk_out);
  wire popcount33_7qyk_core_035;
  wire popcount33_7qyk_core_036;
  wire popcount33_7qyk_core_037;
  wire popcount33_7qyk_core_041;
  wire popcount33_7qyk_core_043;
  wire popcount33_7qyk_core_044;
  wire popcount33_7qyk_core_046;
  wire popcount33_7qyk_core_048;
  wire popcount33_7qyk_core_049;
  wire popcount33_7qyk_core_055;
  wire popcount33_7qyk_core_056;
  wire popcount33_7qyk_core_057;
  wire popcount33_7qyk_core_058;
  wire popcount33_7qyk_core_059_not;
  wire popcount33_7qyk_core_060;
  wire popcount33_7qyk_core_061;
  wire popcount33_7qyk_core_063;
  wire popcount33_7qyk_core_064;
  wire popcount33_7qyk_core_065_not;
  wire popcount33_7qyk_core_066;
  wire popcount33_7qyk_core_067;
  wire popcount33_7qyk_core_068;
  wire popcount33_7qyk_core_069;
  wire popcount33_7qyk_core_070;
  wire popcount33_7qyk_core_072;
  wire popcount33_7qyk_core_074;
  wire popcount33_7qyk_core_075;
  wire popcount33_7qyk_core_076;
  wire popcount33_7qyk_core_077;
  wire popcount33_7qyk_core_078;
  wire popcount33_7qyk_core_079;
  wire popcount33_7qyk_core_083;
  wire popcount33_7qyk_core_084;
  wire popcount33_7qyk_core_086;
  wire popcount33_7qyk_core_089;
  wire popcount33_7qyk_core_090;
  wire popcount33_7qyk_core_091;
  wire popcount33_7qyk_core_093;
  wire popcount33_7qyk_core_094;
  wire popcount33_7qyk_core_095;
  wire popcount33_7qyk_core_096;
  wire popcount33_7qyk_core_098;
  wire popcount33_7qyk_core_100;
  wire popcount33_7qyk_core_101;
  wire popcount33_7qyk_core_102;
  wire popcount33_7qyk_core_103;
  wire popcount33_7qyk_core_106;
  wire popcount33_7qyk_core_108;
  wire popcount33_7qyk_core_110;
  wire popcount33_7qyk_core_112;
  wire popcount33_7qyk_core_113;
  wire popcount33_7qyk_core_115;
  wire popcount33_7qyk_core_118;
  wire popcount33_7qyk_core_119;
  wire popcount33_7qyk_core_120;
  wire popcount33_7qyk_core_122;
  wire popcount33_7qyk_core_125;
  wire popcount33_7qyk_core_126;
  wire popcount33_7qyk_core_127;
  wire popcount33_7qyk_core_128;
  wire popcount33_7qyk_core_131;
  wire popcount33_7qyk_core_132;
  wire popcount33_7qyk_core_134;
  wire popcount33_7qyk_core_137;
  wire popcount33_7qyk_core_138;
  wire popcount33_7qyk_core_139;
  wire popcount33_7qyk_core_141;
  wire popcount33_7qyk_core_142;
  wire popcount33_7qyk_core_143;
  wire popcount33_7qyk_core_144;
  wire popcount33_7qyk_core_148;
  wire popcount33_7qyk_core_149;
  wire popcount33_7qyk_core_151;
  wire popcount33_7qyk_core_153;
  wire popcount33_7qyk_core_155;
  wire popcount33_7qyk_core_156;
  wire popcount33_7qyk_core_157;
  wire popcount33_7qyk_core_160;
  wire popcount33_7qyk_core_161;
  wire popcount33_7qyk_core_162;
  wire popcount33_7qyk_core_163;
  wire popcount33_7qyk_core_164;
  wire popcount33_7qyk_core_165;
  wire popcount33_7qyk_core_166;
  wire popcount33_7qyk_core_167;
  wire popcount33_7qyk_core_168;
  wire popcount33_7qyk_core_170;
  wire popcount33_7qyk_core_171;
  wire popcount33_7qyk_core_172;
  wire popcount33_7qyk_core_176;
  wire popcount33_7qyk_core_177;
  wire popcount33_7qyk_core_178;
  wire popcount33_7qyk_core_179;
  wire popcount33_7qyk_core_180;
  wire popcount33_7qyk_core_182;
  wire popcount33_7qyk_core_184;
  wire popcount33_7qyk_core_185;
  wire popcount33_7qyk_core_186;
  wire popcount33_7qyk_core_187;
  wire popcount33_7qyk_core_188;
  wire popcount33_7qyk_core_190;
  wire popcount33_7qyk_core_191;
  wire popcount33_7qyk_core_193;
  wire popcount33_7qyk_core_195;
  wire popcount33_7qyk_core_197;
  wire popcount33_7qyk_core_198;
  wire popcount33_7qyk_core_201;
  wire popcount33_7qyk_core_202;
  wire popcount33_7qyk_core_204;
  wire popcount33_7qyk_core_206;
  wire popcount33_7qyk_core_208;
  wire popcount33_7qyk_core_209;
  wire popcount33_7qyk_core_212;
  wire popcount33_7qyk_core_213;
  wire popcount33_7qyk_core_214;
  wire popcount33_7qyk_core_215;
  wire popcount33_7qyk_core_217;
  wire popcount33_7qyk_core_219;
  wire popcount33_7qyk_core_221;
  wire popcount33_7qyk_core_222;
  wire popcount33_7qyk_core_223;
  wire popcount33_7qyk_core_225;
  wire popcount33_7qyk_core_226_not;
  wire popcount33_7qyk_core_227;
  wire popcount33_7qyk_core_228;
  wire popcount33_7qyk_core_229;
  wire popcount33_7qyk_core_231;
  wire popcount33_7qyk_core_234;
  wire popcount33_7qyk_core_235;
  wire popcount33_7qyk_core_236;
  wire popcount33_7qyk_core_237;
  wire popcount33_7qyk_core_238_not;

  assign popcount33_7qyk_core_035 = ~(input_a[19] | input_a[2]);
  assign popcount33_7qyk_core_036 = ~(input_a[20] & input_a[12]);
  assign popcount33_7qyk_core_037 = ~input_a[15];
  assign popcount33_7qyk_core_041 = ~(input_a[19] ^ input_a[31]);
  assign popcount33_7qyk_core_043 = ~input_a[8];
  assign popcount33_7qyk_core_044 = ~input_a[7];
  assign popcount33_7qyk_core_046 = ~input_a[19];
  assign popcount33_7qyk_core_048 = ~input_a[2];
  assign popcount33_7qyk_core_049 = ~(input_a[27] ^ input_a[28]);
  assign popcount33_7qyk_core_055 = input_a[16] ^ input_a[8];
  assign popcount33_7qyk_core_056 = input_a[30] | input_a[32];
  assign popcount33_7qyk_core_057 = ~(input_a[6] ^ input_a[19]);
  assign popcount33_7qyk_core_058 = ~(input_a[17] ^ input_a[17]);
  assign popcount33_7qyk_core_059_not = ~input_a[30];
  assign popcount33_7qyk_core_060 = input_a[5] | input_a[8];
  assign popcount33_7qyk_core_061 = input_a[18] ^ input_a[8];
  assign popcount33_7qyk_core_063 = ~(input_a[31] | input_a[12]);
  assign popcount33_7qyk_core_064 = input_a[31] & input_a[3];
  assign popcount33_7qyk_core_065_not = ~input_a[9];
  assign popcount33_7qyk_core_066 = input_a[11] & input_a[22];
  assign popcount33_7qyk_core_067 = ~(input_a[14] & input_a[28]);
  assign popcount33_7qyk_core_068 = input_a[29] & input_a[29];
  assign popcount33_7qyk_core_069 = ~input_a[11];
  assign popcount33_7qyk_core_070 = ~(input_a[32] | input_a[23]);
  assign popcount33_7qyk_core_072 = input_a[9] ^ input_a[7];
  assign popcount33_7qyk_core_074 = ~(input_a[25] & input_a[7]);
  assign popcount33_7qyk_core_075 = ~(input_a[32] & input_a[30]);
  assign popcount33_7qyk_core_076 = input_a[16] | input_a[9];
  assign popcount33_7qyk_core_077 = input_a[21] | input_a[31];
  assign popcount33_7qyk_core_078 = input_a[6] | input_a[1];
  assign popcount33_7qyk_core_079 = ~input_a[30];
  assign popcount33_7qyk_core_083 = ~(input_a[27] ^ input_a[7]);
  assign popcount33_7qyk_core_084 = ~(input_a[7] ^ input_a[23]);
  assign popcount33_7qyk_core_086 = ~(input_a[0] ^ input_a[17]);
  assign popcount33_7qyk_core_089 = input_a[2] | input_a[0];
  assign popcount33_7qyk_core_090 = ~(input_a[7] & input_a[8]);
  assign popcount33_7qyk_core_091 = input_a[11] | input_a[27];
  assign popcount33_7qyk_core_093 = ~(input_a[21] & input_a[0]);
  assign popcount33_7qyk_core_094 = input_a[13] | input_a[30];
  assign popcount33_7qyk_core_095 = input_a[16] ^ input_a[20];
  assign popcount33_7qyk_core_096 = ~input_a[24];
  assign popcount33_7qyk_core_098 = ~(input_a[11] & input_a[19]);
  assign popcount33_7qyk_core_100 = input_a[30] ^ input_a[30];
  assign popcount33_7qyk_core_101 = ~(input_a[11] | input_a[12]);
  assign popcount33_7qyk_core_102 = input_a[26] ^ input_a[6];
  assign popcount33_7qyk_core_103 = ~(input_a[7] | input_a[4]);
  assign popcount33_7qyk_core_106 = input_a[12] & input_a[9];
  assign popcount33_7qyk_core_108 = input_a[32] | input_a[21];
  assign popcount33_7qyk_core_110 = ~input_a[18];
  assign popcount33_7qyk_core_112 = input_a[22] | input_a[28];
  assign popcount33_7qyk_core_113 = input_a[30] ^ input_a[16];
  assign popcount33_7qyk_core_115 = input_a[0] ^ input_a[15];
  assign popcount33_7qyk_core_118 = ~input_a[4];
  assign popcount33_7qyk_core_119 = ~input_a[17];
  assign popcount33_7qyk_core_120 = input_a[6] & input_a[7];
  assign popcount33_7qyk_core_122 = ~(input_a[24] | input_a[5]);
  assign popcount33_7qyk_core_125 = ~(input_a[16] & input_a[4]);
  assign popcount33_7qyk_core_126 = ~(input_a[7] & input_a[7]);
  assign popcount33_7qyk_core_127 = ~(input_a[9] & input_a[13]);
  assign popcount33_7qyk_core_128 = input_a[32] ^ input_a[21];
  assign popcount33_7qyk_core_131 = ~(input_a[9] ^ input_a[4]);
  assign popcount33_7qyk_core_132 = input_a[21] | input_a[10];
  assign popcount33_7qyk_core_134 = ~(input_a[2] ^ input_a[2]);
  assign popcount33_7qyk_core_137 = input_a[30] & input_a[15];
  assign popcount33_7qyk_core_138 = input_a[15] ^ input_a[8];
  assign popcount33_7qyk_core_139 = ~(input_a[0] & input_a[3]);
  assign popcount33_7qyk_core_141 = ~(input_a[31] ^ input_a[8]);
  assign popcount33_7qyk_core_142 = ~(input_a[24] ^ input_a[16]);
  assign popcount33_7qyk_core_143 = input_a[4] | input_a[5];
  assign popcount33_7qyk_core_144 = input_a[11] & input_a[23];
  assign popcount33_7qyk_core_148 = ~(input_a[27] | input_a[9]);
  assign popcount33_7qyk_core_149 = input_a[8] | input_a[25];
  assign popcount33_7qyk_core_151 = ~input_a[22];
  assign popcount33_7qyk_core_153 = ~input_a[28];
  assign popcount33_7qyk_core_155 = input_a[22] | input_a[9];
  assign popcount33_7qyk_core_156 = input_a[5] & input_a[0];
  assign popcount33_7qyk_core_157 = ~(input_a[13] | input_a[15]);
  assign popcount33_7qyk_core_160 = ~(input_a[26] & input_a[13]);
  assign popcount33_7qyk_core_161 = ~(input_a[3] ^ input_a[3]);
  assign popcount33_7qyk_core_162 = ~input_a[28];
  assign popcount33_7qyk_core_163 = input_a[29] ^ input_a[1];
  assign popcount33_7qyk_core_164 = ~input_a[31];
  assign popcount33_7qyk_core_165 = input_a[4] | input_a[10];
  assign popcount33_7qyk_core_166 = input_a[32] ^ input_a[31];
  assign popcount33_7qyk_core_167 = input_a[32] ^ input_a[24];
  assign popcount33_7qyk_core_168 = ~input_a[4];
  assign popcount33_7qyk_core_170 = input_a[10] ^ input_a[20];
  assign popcount33_7qyk_core_171 = ~input_a[24];
  assign popcount33_7qyk_core_172 = ~(input_a[2] & input_a[21]);
  assign popcount33_7qyk_core_176 = input_a[25] & input_a[13];
  assign popcount33_7qyk_core_177 = ~(input_a[13] | input_a[10]);
  assign popcount33_7qyk_core_178 = input_a[1] & input_a[11];
  assign popcount33_7qyk_core_179 = ~(input_a[16] & input_a[28]);
  assign popcount33_7qyk_core_180 = ~(input_a[3] | input_a[1]);
  assign popcount33_7qyk_core_182 = ~(input_a[28] | input_a[14]);
  assign popcount33_7qyk_core_184 = ~(input_a[6] | input_a[21]);
  assign popcount33_7qyk_core_185 = ~(input_a[7] & input_a[29]);
  assign popcount33_7qyk_core_186 = input_a[29] | input_a[2];
  assign popcount33_7qyk_core_187 = input_a[20] | input_a[9];
  assign popcount33_7qyk_core_188 = ~(input_a[6] | input_a[29]);
  assign popcount33_7qyk_core_190 = ~(input_a[1] ^ input_a[20]);
  assign popcount33_7qyk_core_191 = input_a[20] ^ input_a[21];
  assign popcount33_7qyk_core_193 = input_a[15] | input_a[16];
  assign popcount33_7qyk_core_195 = input_a[0] & input_a[30];
  assign popcount33_7qyk_core_197 = input_a[18] ^ input_a[19];
  assign popcount33_7qyk_core_198 = input_a[30] ^ input_a[4];
  assign popcount33_7qyk_core_201 = input_a[11] & input_a[19];
  assign popcount33_7qyk_core_202 = ~(input_a[0] & input_a[2]);
  assign popcount33_7qyk_core_204 = ~(input_a[26] | input_a[23]);
  assign popcount33_7qyk_core_206 = ~(input_a[8] ^ input_a[32]);
  assign popcount33_7qyk_core_208 = ~(input_a[9] | input_a[22]);
  assign popcount33_7qyk_core_209 = ~(input_a[26] | input_a[14]);
  assign popcount33_7qyk_core_212 = input_a[22] ^ input_a[12];
  assign popcount33_7qyk_core_213 = ~(input_a[13] ^ input_a[26]);
  assign popcount33_7qyk_core_214 = ~input_a[30];
  assign popcount33_7qyk_core_215 = input_a[29] | input_a[28];
  assign popcount33_7qyk_core_217 = ~(input_a[23] | input_a[20]);
  assign popcount33_7qyk_core_219 = input_a[20] ^ input_a[0];
  assign popcount33_7qyk_core_221 = ~input_a[19];
  assign popcount33_7qyk_core_222 = ~(input_a[23] & input_a[22]);
  assign popcount33_7qyk_core_223 = input_a[13] & input_a[24];
  assign popcount33_7qyk_core_225 = ~input_a[27];
  assign popcount33_7qyk_core_226_not = ~input_a[2];
  assign popcount33_7qyk_core_227 = input_a[15] | input_a[5];
  assign popcount33_7qyk_core_228 = input_a[14] ^ input_a[10];
  assign popcount33_7qyk_core_229 = ~(input_a[13] & input_a[22]);
  assign popcount33_7qyk_core_231 = ~(input_a[8] | input_a[27]);
  assign popcount33_7qyk_core_234 = ~(input_a[10] & input_a[4]);
  assign popcount33_7qyk_core_235 = input_a[10] & input_a[17];
  assign popcount33_7qyk_core_236 = input_a[13] & input_a[11];
  assign popcount33_7qyk_core_237 = ~(input_a[21] ^ input_a[21]);
  assign popcount33_7qyk_core_238_not = ~input_a[32];

  assign popcount33_7qyk_out[0] = 1'b0;
  assign popcount33_7qyk_out[1] = 1'b0;
  assign popcount33_7qyk_out[2] = input_a[17];
  assign popcount33_7qyk_out[3] = input_a[5];
  assign popcount33_7qyk_out[4] = input_a[1];
  assign popcount33_7qyk_out[5] = 1'b0;
endmodule