// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=16.2853
// WCE=50.0
// EP=0.97046%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_75jl(input [37:0] input_a, output [5:0] popcount38_75jl_out);
  wire popcount38_75jl_core_040;
  wire popcount38_75jl_core_041;
  wire popcount38_75jl_core_042;
  wire popcount38_75jl_core_044;
  wire popcount38_75jl_core_047;
  wire popcount38_75jl_core_048;
  wire popcount38_75jl_core_049;
  wire popcount38_75jl_core_050;
  wire popcount38_75jl_core_051;
  wire popcount38_75jl_core_052;
  wire popcount38_75jl_core_054;
  wire popcount38_75jl_core_058;
  wire popcount38_75jl_core_060;
  wire popcount38_75jl_core_061;
  wire popcount38_75jl_core_063;
  wire popcount38_75jl_core_066;
  wire popcount38_75jl_core_068;
  wire popcount38_75jl_core_069;
  wire popcount38_75jl_core_070;
  wire popcount38_75jl_core_071;
  wire popcount38_75jl_core_072;
  wire popcount38_75jl_core_073;
  wire popcount38_75jl_core_075;
  wire popcount38_75jl_core_077;
  wire popcount38_75jl_core_078;
  wire popcount38_75jl_core_082;
  wire popcount38_75jl_core_084;
  wire popcount38_75jl_core_088;
  wire popcount38_75jl_core_089;
  wire popcount38_75jl_core_091;
  wire popcount38_75jl_core_092;
  wire popcount38_75jl_core_095;
  wire popcount38_75jl_core_096;
  wire popcount38_75jl_core_098;
  wire popcount38_75jl_core_099;
  wire popcount38_75jl_core_101;
  wire popcount38_75jl_core_104;
  wire popcount38_75jl_core_105;
  wire popcount38_75jl_core_108;
  wire popcount38_75jl_core_109;
  wire popcount38_75jl_core_110;
  wire popcount38_75jl_core_111;
  wire popcount38_75jl_core_112;
  wire popcount38_75jl_core_114;
  wire popcount38_75jl_core_115;
  wire popcount38_75jl_core_117;
  wire popcount38_75jl_core_118;
  wire popcount38_75jl_core_119;
  wire popcount38_75jl_core_120;
  wire popcount38_75jl_core_122;
  wire popcount38_75jl_core_125;
  wire popcount38_75jl_core_126;
  wire popcount38_75jl_core_127_not;
  wire popcount38_75jl_core_128;
  wire popcount38_75jl_core_130;
  wire popcount38_75jl_core_131;
  wire popcount38_75jl_core_132;
  wire popcount38_75jl_core_133;
  wire popcount38_75jl_core_134;
  wire popcount38_75jl_core_135;
  wire popcount38_75jl_core_137;
  wire popcount38_75jl_core_139;
  wire popcount38_75jl_core_140_not;
  wire popcount38_75jl_core_141_not;
  wire popcount38_75jl_core_142;
  wire popcount38_75jl_core_143;
  wire popcount38_75jl_core_144;
  wire popcount38_75jl_core_146;
  wire popcount38_75jl_core_147;
  wire popcount38_75jl_core_149;
  wire popcount38_75jl_core_152;
  wire popcount38_75jl_core_153;
  wire popcount38_75jl_core_155;
  wire popcount38_75jl_core_156;
  wire popcount38_75jl_core_158;
  wire popcount38_75jl_core_159;
  wire popcount38_75jl_core_161;
  wire popcount38_75jl_core_162;
  wire popcount38_75jl_core_163;
  wire popcount38_75jl_core_166;
  wire popcount38_75jl_core_167;
  wire popcount38_75jl_core_170;
  wire popcount38_75jl_core_171;
  wire popcount38_75jl_core_172;
  wire popcount38_75jl_core_173;
  wire popcount38_75jl_core_174;
  wire popcount38_75jl_core_175;
  wire popcount38_75jl_core_176;
  wire popcount38_75jl_core_179;
  wire popcount38_75jl_core_180;
  wire popcount38_75jl_core_181;
  wire popcount38_75jl_core_182;
  wire popcount38_75jl_core_183;
  wire popcount38_75jl_core_184;
  wire popcount38_75jl_core_185;
  wire popcount38_75jl_core_186;
  wire popcount38_75jl_core_187;
  wire popcount38_75jl_core_188;
  wire popcount38_75jl_core_191;
  wire popcount38_75jl_core_193;
  wire popcount38_75jl_core_194;
  wire popcount38_75jl_core_195;
  wire popcount38_75jl_core_199;
  wire popcount38_75jl_core_200;
  wire popcount38_75jl_core_201;
  wire popcount38_75jl_core_202;
  wire popcount38_75jl_core_204;
  wire popcount38_75jl_core_205;
  wire popcount38_75jl_core_206;
  wire popcount38_75jl_core_208;
  wire popcount38_75jl_core_209;
  wire popcount38_75jl_core_211;
  wire popcount38_75jl_core_212;
  wire popcount38_75jl_core_213;
  wire popcount38_75jl_core_214;
  wire popcount38_75jl_core_215;
  wire popcount38_75jl_core_216;
  wire popcount38_75jl_core_218;
  wire popcount38_75jl_core_219;
  wire popcount38_75jl_core_220;
  wire popcount38_75jl_core_221;
  wire popcount38_75jl_core_224;
  wire popcount38_75jl_core_225_not;
  wire popcount38_75jl_core_226;
  wire popcount38_75jl_core_228;
  wire popcount38_75jl_core_230;
  wire popcount38_75jl_core_232;
  wire popcount38_75jl_core_233;
  wire popcount38_75jl_core_235;
  wire popcount38_75jl_core_236;
  wire popcount38_75jl_core_239;
  wire popcount38_75jl_core_240;
  wire popcount38_75jl_core_242;
  wire popcount38_75jl_core_243;
  wire popcount38_75jl_core_244;
  wire popcount38_75jl_core_245;
  wire popcount38_75jl_core_246;
  wire popcount38_75jl_core_247;
  wire popcount38_75jl_core_249;
  wire popcount38_75jl_core_250;
  wire popcount38_75jl_core_251;
  wire popcount38_75jl_core_253;
  wire popcount38_75jl_core_254;
  wire popcount38_75jl_core_256;
  wire popcount38_75jl_core_258;
  wire popcount38_75jl_core_259;
  wire popcount38_75jl_core_260;
  wire popcount38_75jl_core_261;
  wire popcount38_75jl_core_262;
  wire popcount38_75jl_core_263;
  wire popcount38_75jl_core_264;
  wire popcount38_75jl_core_265;
  wire popcount38_75jl_core_266;
  wire popcount38_75jl_core_267;
  wire popcount38_75jl_core_268;
  wire popcount38_75jl_core_271;
  wire popcount38_75jl_core_272;
  wire popcount38_75jl_core_274;
  wire popcount38_75jl_core_276;
  wire popcount38_75jl_core_277;
  wire popcount38_75jl_core_278;
  wire popcount38_75jl_core_280;
  wire popcount38_75jl_core_281;
  wire popcount38_75jl_core_283;
  wire popcount38_75jl_core_285;
  wire popcount38_75jl_core_286;
  wire popcount38_75jl_core_290;
  wire popcount38_75jl_core_291;
  wire popcount38_75jl_core_292;
  wire popcount38_75jl_core_293;

  assign popcount38_75jl_core_040 = ~input_a[3];
  assign popcount38_75jl_core_041 = ~(input_a[34] ^ input_a[37]);
  assign popcount38_75jl_core_042 = input_a[28] | input_a[31];
  assign popcount38_75jl_core_044 = ~input_a[7];
  assign popcount38_75jl_core_047 = input_a[35] ^ input_a[22];
  assign popcount38_75jl_core_048 = ~(input_a[28] | input_a[18]);
  assign popcount38_75jl_core_049 = input_a[21] | input_a[28];
  assign popcount38_75jl_core_050 = ~(input_a[22] ^ input_a[33]);
  assign popcount38_75jl_core_051 = ~(input_a[26] | input_a[19]);
  assign popcount38_75jl_core_052 = input_a[36] ^ input_a[22];
  assign popcount38_75jl_core_054 = ~(input_a[24] & input_a[18]);
  assign popcount38_75jl_core_058 = input_a[34] ^ input_a[25];
  assign popcount38_75jl_core_060 = ~(input_a[30] | input_a[24]);
  assign popcount38_75jl_core_061 = ~(input_a[18] | input_a[22]);
  assign popcount38_75jl_core_063 = input_a[24] | input_a[31];
  assign popcount38_75jl_core_066 = ~(input_a[8] ^ input_a[7]);
  assign popcount38_75jl_core_068 = input_a[24] & input_a[25];
  assign popcount38_75jl_core_069 = ~input_a[7];
  assign popcount38_75jl_core_070 = input_a[19] | input_a[10];
  assign popcount38_75jl_core_071 = input_a[14] ^ input_a[6];
  assign popcount38_75jl_core_072 = ~input_a[22];
  assign popcount38_75jl_core_073 = input_a[23] ^ input_a[6];
  assign popcount38_75jl_core_075 = ~(input_a[26] & input_a[17]);
  assign popcount38_75jl_core_077 = input_a[6] | input_a[7];
  assign popcount38_75jl_core_078 = ~(input_a[14] | input_a[27]);
  assign popcount38_75jl_core_082 = ~input_a[34];
  assign popcount38_75jl_core_084 = input_a[17] | input_a[27];
  assign popcount38_75jl_core_088 = ~(input_a[4] | input_a[14]);
  assign popcount38_75jl_core_089 = ~(input_a[6] | input_a[14]);
  assign popcount38_75jl_core_091 = ~(input_a[34] | input_a[37]);
  assign popcount38_75jl_core_092 = ~input_a[18];
  assign popcount38_75jl_core_095 = ~(input_a[15] & input_a[27]);
  assign popcount38_75jl_core_096 = ~(input_a[34] ^ input_a[1]);
  assign popcount38_75jl_core_098 = input_a[7] & input_a[22];
  assign popcount38_75jl_core_099 = ~(input_a[14] & input_a[5]);
  assign popcount38_75jl_core_101 = ~(input_a[17] ^ input_a[32]);
  assign popcount38_75jl_core_104 = ~(input_a[6] ^ input_a[19]);
  assign popcount38_75jl_core_105 = ~input_a[28];
  assign popcount38_75jl_core_108 = ~input_a[7];
  assign popcount38_75jl_core_109 = ~(input_a[0] & input_a[7]);
  assign popcount38_75jl_core_110 = input_a[28] ^ input_a[7];
  assign popcount38_75jl_core_111 = ~(input_a[37] ^ input_a[29]);
  assign popcount38_75jl_core_112 = ~(input_a[9] ^ input_a[25]);
  assign popcount38_75jl_core_114 = input_a[33] ^ input_a[30];
  assign popcount38_75jl_core_115 = input_a[15] & input_a[3];
  assign popcount38_75jl_core_117 = ~(input_a[17] | input_a[19]);
  assign popcount38_75jl_core_118 = input_a[29] ^ input_a[12];
  assign popcount38_75jl_core_119 = ~(input_a[14] | input_a[36]);
  assign popcount38_75jl_core_120 = ~(input_a[8] & input_a[16]);
  assign popcount38_75jl_core_122 = input_a[37] ^ input_a[32];
  assign popcount38_75jl_core_125 = input_a[19] ^ input_a[12];
  assign popcount38_75jl_core_126 = ~(input_a[29] ^ input_a[2]);
  assign popcount38_75jl_core_127_not = ~input_a[5];
  assign popcount38_75jl_core_128 = ~(input_a[27] & input_a[33]);
  assign popcount38_75jl_core_130 = ~(input_a[28] | input_a[1]);
  assign popcount38_75jl_core_131 = input_a[34] | input_a[20];
  assign popcount38_75jl_core_132 = ~(input_a[33] ^ input_a[4]);
  assign popcount38_75jl_core_133 = ~(input_a[11] | input_a[13]);
  assign popcount38_75jl_core_134 = ~(input_a[22] | input_a[20]);
  assign popcount38_75jl_core_135 = ~input_a[6];
  assign popcount38_75jl_core_137 = input_a[32] & input_a[19];
  assign popcount38_75jl_core_139 = input_a[20] | input_a[32];
  assign popcount38_75jl_core_140_not = ~input_a[15];
  assign popcount38_75jl_core_141_not = ~input_a[33];
  assign popcount38_75jl_core_142 = ~(input_a[2] | input_a[9]);
  assign popcount38_75jl_core_143 = ~(input_a[34] | input_a[26]);
  assign popcount38_75jl_core_144 = ~input_a[16];
  assign popcount38_75jl_core_146 = input_a[2] | input_a[19];
  assign popcount38_75jl_core_147 = input_a[9] ^ input_a[18];
  assign popcount38_75jl_core_149 = input_a[5] | input_a[15];
  assign popcount38_75jl_core_152 = input_a[29] & input_a[10];
  assign popcount38_75jl_core_153 = input_a[14] | input_a[10];
  assign popcount38_75jl_core_155 = ~(input_a[18] & input_a[34]);
  assign popcount38_75jl_core_156 = ~(input_a[25] | input_a[29]);
  assign popcount38_75jl_core_158 = ~(input_a[3] ^ input_a[25]);
  assign popcount38_75jl_core_159 = ~input_a[14];
  assign popcount38_75jl_core_161 = input_a[12] | input_a[16];
  assign popcount38_75jl_core_162 = input_a[24] ^ input_a[29];
  assign popcount38_75jl_core_163 = ~(input_a[19] & input_a[22]);
  assign popcount38_75jl_core_166 = ~input_a[20];
  assign popcount38_75jl_core_167 = ~(input_a[2] ^ input_a[20]);
  assign popcount38_75jl_core_170 = input_a[17] | input_a[15];
  assign popcount38_75jl_core_171 = ~(input_a[7] & input_a[37]);
  assign popcount38_75jl_core_172 = ~(input_a[37] | input_a[37]);
  assign popcount38_75jl_core_173 = ~(input_a[15] | input_a[8]);
  assign popcount38_75jl_core_174 = ~(input_a[19] ^ input_a[0]);
  assign popcount38_75jl_core_175 = ~(input_a[17] ^ input_a[29]);
  assign popcount38_75jl_core_176 = ~input_a[22];
  assign popcount38_75jl_core_179 = ~(input_a[6] & input_a[26]);
  assign popcount38_75jl_core_180 = ~(input_a[30] | input_a[17]);
  assign popcount38_75jl_core_181 = input_a[35] | input_a[22];
  assign popcount38_75jl_core_182 = input_a[32] & input_a[30];
  assign popcount38_75jl_core_183 = ~(input_a[30] & input_a[16]);
  assign popcount38_75jl_core_184 = ~(input_a[5] & input_a[28]);
  assign popcount38_75jl_core_185 = ~(input_a[8] ^ input_a[16]);
  assign popcount38_75jl_core_186 = input_a[15] | input_a[34];
  assign popcount38_75jl_core_187 = ~(input_a[15] | input_a[37]);
  assign popcount38_75jl_core_188 = ~(input_a[13] & input_a[0]);
  assign popcount38_75jl_core_191 = ~(input_a[35] & input_a[29]);
  assign popcount38_75jl_core_193 = ~(input_a[4] & input_a[28]);
  assign popcount38_75jl_core_194 = ~input_a[1];
  assign popcount38_75jl_core_195 = input_a[0] | input_a[23];
  assign popcount38_75jl_core_199 = input_a[9] | input_a[34];
  assign popcount38_75jl_core_200 = input_a[13] & input_a[28];
  assign popcount38_75jl_core_201 = ~(input_a[34] ^ input_a[19]);
  assign popcount38_75jl_core_202 = ~(input_a[9] ^ input_a[6]);
  assign popcount38_75jl_core_204 = ~(input_a[37] ^ input_a[1]);
  assign popcount38_75jl_core_205 = input_a[6] & input_a[31];
  assign popcount38_75jl_core_206 = input_a[19] | input_a[27];
  assign popcount38_75jl_core_208 = ~(input_a[32] | input_a[3]);
  assign popcount38_75jl_core_209 = ~(input_a[25] & input_a[13]);
  assign popcount38_75jl_core_211 = ~input_a[19];
  assign popcount38_75jl_core_212 = ~(input_a[12] ^ input_a[37]);
  assign popcount38_75jl_core_213 = ~(input_a[9] | input_a[25]);
  assign popcount38_75jl_core_214 = input_a[37] | input_a[31];
  assign popcount38_75jl_core_215 = ~(input_a[2] & input_a[7]);
  assign popcount38_75jl_core_216 = input_a[33] ^ input_a[33];
  assign popcount38_75jl_core_218 = input_a[9] | input_a[17];
  assign popcount38_75jl_core_219 = input_a[23] ^ input_a[3];
  assign popcount38_75jl_core_220 = input_a[35] ^ input_a[1];
  assign popcount38_75jl_core_221 = input_a[34] & input_a[16];
  assign popcount38_75jl_core_224 = input_a[31] & input_a[28];
  assign popcount38_75jl_core_225_not = ~input_a[23];
  assign popcount38_75jl_core_226 = input_a[14] & input_a[27];
  assign popcount38_75jl_core_228 = ~(input_a[18] & input_a[33]);
  assign popcount38_75jl_core_230 = input_a[10] & input_a[3];
  assign popcount38_75jl_core_232 = ~(input_a[12] ^ input_a[1]);
  assign popcount38_75jl_core_233 = ~(input_a[35] ^ input_a[0]);
  assign popcount38_75jl_core_235 = ~(input_a[31] | input_a[9]);
  assign popcount38_75jl_core_236 = input_a[8] | input_a[10];
  assign popcount38_75jl_core_239 = ~input_a[5];
  assign popcount38_75jl_core_240 = ~input_a[17];
  assign popcount38_75jl_core_242 = input_a[37] | input_a[33];
  assign popcount38_75jl_core_243 = input_a[4] | input_a[31];
  assign popcount38_75jl_core_244 = ~(input_a[5] ^ input_a[9]);
  assign popcount38_75jl_core_245 = input_a[16] | input_a[30];
  assign popcount38_75jl_core_246 = ~input_a[34];
  assign popcount38_75jl_core_247 = input_a[27] | input_a[4];
  assign popcount38_75jl_core_249 = ~(input_a[24] & input_a[20]);
  assign popcount38_75jl_core_250 = ~(input_a[8] & input_a[35]);
  assign popcount38_75jl_core_251 = input_a[26] & input_a[27];
  assign popcount38_75jl_core_253 = ~(input_a[10] ^ input_a[10]);
  assign popcount38_75jl_core_254 = input_a[29] ^ input_a[3];
  assign popcount38_75jl_core_256 = ~(input_a[24] & input_a[2]);
  assign popcount38_75jl_core_258 = ~(input_a[26] ^ input_a[32]);
  assign popcount38_75jl_core_259 = ~(input_a[11] & input_a[20]);
  assign popcount38_75jl_core_260 = ~input_a[15];
  assign popcount38_75jl_core_261 = ~(input_a[16] & input_a[37]);
  assign popcount38_75jl_core_262 = input_a[34] & input_a[9];
  assign popcount38_75jl_core_263 = input_a[18] ^ input_a[10];
  assign popcount38_75jl_core_264 = ~(input_a[22] | input_a[3]);
  assign popcount38_75jl_core_265 = ~input_a[4];
  assign popcount38_75jl_core_266 = input_a[33] | input_a[5];
  assign popcount38_75jl_core_267 = input_a[5] | input_a[3];
  assign popcount38_75jl_core_268 = ~(input_a[9] & input_a[4]);
  assign popcount38_75jl_core_271 = input_a[20] & input_a[31];
  assign popcount38_75jl_core_272 = input_a[32] & input_a[24];
  assign popcount38_75jl_core_274 = ~(input_a[21] | input_a[28]);
  assign popcount38_75jl_core_276 = input_a[20] | input_a[4];
  assign popcount38_75jl_core_277 = input_a[17] & input_a[18];
  assign popcount38_75jl_core_278 = input_a[37] ^ input_a[35];
  assign popcount38_75jl_core_280 = ~(input_a[2] ^ input_a[12]);
  assign popcount38_75jl_core_281 = ~(input_a[16] | input_a[3]);
  assign popcount38_75jl_core_283 = input_a[14] ^ input_a[0];
  assign popcount38_75jl_core_285 = input_a[37] | input_a[26];
  assign popcount38_75jl_core_286 = ~(input_a[2] & input_a[34]);
  assign popcount38_75jl_core_290 = ~(input_a[0] & input_a[28]);
  assign popcount38_75jl_core_291 = input_a[35] | input_a[12];
  assign popcount38_75jl_core_292 = ~input_a[30];
  assign popcount38_75jl_core_293 = input_a[25] & input_a[27];

  assign popcount38_75jl_out[0] = input_a[18];
  assign popcount38_75jl_out[1] = input_a[20];
  assign popcount38_75jl_out[2] = input_a[26];
  assign popcount38_75jl_out[3] = 1'b0;
  assign popcount38_75jl_out[4] = input_a[37];
  assign popcount38_75jl_out[5] = input_a[33];
endmodule