// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.5904
// WCE=15.0
// EP=0.880443%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_2mwl(input [24:0] input_a, output [4:0] popcount25_2mwl_out);
  wire popcount25_2mwl_core_028;
  wire popcount25_2mwl_core_029_not;
  wire popcount25_2mwl_core_030;
  wire popcount25_2mwl_core_031;
  wire popcount25_2mwl_core_032;
  wire popcount25_2mwl_core_033;
  wire popcount25_2mwl_core_034;
  wire popcount25_2mwl_core_035;
  wire popcount25_2mwl_core_036;
  wire popcount25_2mwl_core_037;
  wire popcount25_2mwl_core_038;
  wire popcount25_2mwl_core_040;
  wire popcount25_2mwl_core_041;
  wire popcount25_2mwl_core_042;
  wire popcount25_2mwl_core_043;
  wire popcount25_2mwl_core_044;
  wire popcount25_2mwl_core_045;
  wire popcount25_2mwl_core_046;
  wire popcount25_2mwl_core_047;
  wire popcount25_2mwl_core_049;
  wire popcount25_2mwl_core_052;
  wire popcount25_2mwl_core_057;
  wire popcount25_2mwl_core_058;
  wire popcount25_2mwl_core_059;
  wire popcount25_2mwl_core_060;
  wire popcount25_2mwl_core_061;
  wire popcount25_2mwl_core_063;
  wire popcount25_2mwl_core_067;
  wire popcount25_2mwl_core_069;
  wire popcount25_2mwl_core_071;
  wire popcount25_2mwl_core_072;
  wire popcount25_2mwl_core_073;
  wire popcount25_2mwl_core_076;
  wire popcount25_2mwl_core_078;
  wire popcount25_2mwl_core_079_not;
  wire popcount25_2mwl_core_081;
  wire popcount25_2mwl_core_082;
  wire popcount25_2mwl_core_083;
  wire popcount25_2mwl_core_085;
  wire popcount25_2mwl_core_090;
  wire popcount25_2mwl_core_091;
  wire popcount25_2mwl_core_096_not;
  wire popcount25_2mwl_core_097;
  wire popcount25_2mwl_core_098;
  wire popcount25_2mwl_core_099;
  wire popcount25_2mwl_core_100;
  wire popcount25_2mwl_core_101;
  wire popcount25_2mwl_core_102;
  wire popcount25_2mwl_core_103;
  wire popcount25_2mwl_core_104;
  wire popcount25_2mwl_core_105_not;
  wire popcount25_2mwl_core_106;
  wire popcount25_2mwl_core_107;
  wire popcount25_2mwl_core_110;
  wire popcount25_2mwl_core_111;
  wire popcount25_2mwl_core_112;
  wire popcount25_2mwl_core_113;
  wire popcount25_2mwl_core_114;
  wire popcount25_2mwl_core_115;
  wire popcount25_2mwl_core_118;
  wire popcount25_2mwl_core_119;
  wire popcount25_2mwl_core_121;
  wire popcount25_2mwl_core_124;
  wire popcount25_2mwl_core_129;
  wire popcount25_2mwl_core_131;
  wire popcount25_2mwl_core_132;
  wire popcount25_2mwl_core_133;
  wire popcount25_2mwl_core_134;
  wire popcount25_2mwl_core_135;
  wire popcount25_2mwl_core_136;
  wire popcount25_2mwl_core_139;
  wire popcount25_2mwl_core_143;
  wire popcount25_2mwl_core_146;
  wire popcount25_2mwl_core_155;
  wire popcount25_2mwl_core_156;
  wire popcount25_2mwl_core_159;
  wire popcount25_2mwl_core_160;
  wire popcount25_2mwl_core_161;
  wire popcount25_2mwl_core_162;
  wire popcount25_2mwl_core_164;
  wire popcount25_2mwl_core_167;
  wire popcount25_2mwl_core_169;
  wire popcount25_2mwl_core_171;
  wire popcount25_2mwl_core_172;
  wire popcount25_2mwl_core_173;
  wire popcount25_2mwl_core_174_not;
  wire popcount25_2mwl_core_175;
  wire popcount25_2mwl_core_177;
  wire popcount25_2mwl_core_178;
  wire popcount25_2mwl_core_179;
  wire popcount25_2mwl_core_181;
  wire popcount25_2mwl_core_183;

  assign popcount25_2mwl_core_028 = ~(input_a[9] | input_a[18]);
  assign popcount25_2mwl_core_029_not = ~input_a[7];
  assign popcount25_2mwl_core_030 = ~(input_a[20] & input_a[9]);
  assign popcount25_2mwl_core_031 = ~(input_a[17] & input_a[14]);
  assign popcount25_2mwl_core_032 = input_a[3] ^ input_a[9];
  assign popcount25_2mwl_core_033 = input_a[3] ^ input_a[2];
  assign popcount25_2mwl_core_034 = input_a[2] & input_a[23];
  assign popcount25_2mwl_core_035 = ~(input_a[4] ^ input_a[4]);
  assign popcount25_2mwl_core_036 = ~(input_a[0] ^ input_a[10]);
  assign popcount25_2mwl_core_037 = ~(input_a[24] ^ input_a[1]);
  assign popcount25_2mwl_core_038 = ~(input_a[17] ^ input_a[24]);
  assign popcount25_2mwl_core_040 = ~(input_a[22] & input_a[23]);
  assign popcount25_2mwl_core_041 = input_a[2] ^ input_a[7];
  assign popcount25_2mwl_core_042 = ~(input_a[8] | input_a[19]);
  assign popcount25_2mwl_core_043 = input_a[1] | input_a[22];
  assign popcount25_2mwl_core_044 = ~input_a[4];
  assign popcount25_2mwl_core_045 = input_a[12] ^ input_a[11];
  assign popcount25_2mwl_core_046 = ~input_a[4];
  assign popcount25_2mwl_core_047 = ~input_a[1];
  assign popcount25_2mwl_core_049 = ~(input_a[23] | input_a[22]);
  assign popcount25_2mwl_core_052 = ~(input_a[3] ^ input_a[17]);
  assign popcount25_2mwl_core_057 = input_a[2] & input_a[23];
  assign popcount25_2mwl_core_058 = input_a[24] ^ input_a[1];
  assign popcount25_2mwl_core_059 = input_a[3] ^ input_a[17];
  assign popcount25_2mwl_core_060 = input_a[3] & input_a[3];
  assign popcount25_2mwl_core_061 = input_a[2] | input_a[3];
  assign popcount25_2mwl_core_063 = ~(input_a[14] | input_a[17]);
  assign popcount25_2mwl_core_067 = input_a[18] | input_a[19];
  assign popcount25_2mwl_core_069 = ~(input_a[3] | input_a[24]);
  assign popcount25_2mwl_core_071 = ~(input_a[8] & input_a[14]);
  assign popcount25_2mwl_core_072 = input_a[13] ^ input_a[21];
  assign popcount25_2mwl_core_073 = ~(input_a[15] & input_a[19]);
  assign popcount25_2mwl_core_076 = ~(input_a[3] & input_a[18]);
  assign popcount25_2mwl_core_078 = input_a[8] ^ input_a[14];
  assign popcount25_2mwl_core_079_not = ~input_a[18];
  assign popcount25_2mwl_core_081 = ~input_a[6];
  assign popcount25_2mwl_core_082 = ~input_a[3];
  assign popcount25_2mwl_core_083 = ~(input_a[10] ^ input_a[9]);
  assign popcount25_2mwl_core_085 = ~(input_a[22] ^ input_a[6]);
  assign popcount25_2mwl_core_090 = ~(input_a[8] & input_a[1]);
  assign popcount25_2mwl_core_091 = ~(input_a[16] & input_a[17]);
  assign popcount25_2mwl_core_096_not = ~input_a[11];
  assign popcount25_2mwl_core_097 = input_a[18] | input_a[12];
  assign popcount25_2mwl_core_098 = ~(input_a[24] & input_a[11]);
  assign popcount25_2mwl_core_099 = ~(input_a[0] ^ input_a[18]);
  assign popcount25_2mwl_core_100 = ~(input_a[15] ^ input_a[17]);
  assign popcount25_2mwl_core_101 = ~(input_a[1] ^ input_a[15]);
  assign popcount25_2mwl_core_102 = ~(input_a[3] & input_a[7]);
  assign popcount25_2mwl_core_103 = input_a[16] & input_a[3];
  assign popcount25_2mwl_core_104 = ~(input_a[4] & input_a[7]);
  assign popcount25_2mwl_core_105_not = ~input_a[4];
  assign popcount25_2mwl_core_106 = input_a[5] | input_a[18];
  assign popcount25_2mwl_core_107 = ~(input_a[23] ^ input_a[7]);
  assign popcount25_2mwl_core_110 = ~(input_a[19] & input_a[7]);
  assign popcount25_2mwl_core_111 = input_a[4] ^ input_a[10];
  assign popcount25_2mwl_core_112 = ~(input_a[3] | input_a[12]);
  assign popcount25_2mwl_core_113 = ~(input_a[4] | input_a[6]);
  assign popcount25_2mwl_core_114 = ~input_a[1];
  assign popcount25_2mwl_core_115 = input_a[20] | input_a[22];
  assign popcount25_2mwl_core_118 = ~(input_a[21] | input_a[5]);
  assign popcount25_2mwl_core_119 = input_a[0] & input_a[16];
  assign popcount25_2mwl_core_121 = ~(input_a[5] & input_a[15]);
  assign popcount25_2mwl_core_124 = input_a[24] ^ input_a[11];
  assign popcount25_2mwl_core_129 = ~(input_a[18] ^ input_a[22]);
  assign popcount25_2mwl_core_131 = ~(input_a[9] | input_a[21]);
  assign popcount25_2mwl_core_132 = input_a[5] & input_a[22];
  assign popcount25_2mwl_core_133 = ~input_a[12];
  assign popcount25_2mwl_core_134 = input_a[21] ^ input_a[14];
  assign popcount25_2mwl_core_135 = input_a[13] | input_a[4];
  assign popcount25_2mwl_core_136 = ~(input_a[8] ^ input_a[12]);
  assign popcount25_2mwl_core_139 = input_a[4] & input_a[16];
  assign popcount25_2mwl_core_143 = input_a[15] | input_a[5];
  assign popcount25_2mwl_core_146 = ~(input_a[22] | input_a[12]);
  assign popcount25_2mwl_core_155 = ~(input_a[18] ^ input_a[9]);
  assign popcount25_2mwl_core_156 = ~(input_a[10] ^ input_a[18]);
  assign popcount25_2mwl_core_159 = ~(input_a[18] | input_a[20]);
  assign popcount25_2mwl_core_160 = ~(input_a[15] & input_a[19]);
  assign popcount25_2mwl_core_161 = ~(input_a[1] ^ input_a[24]);
  assign popcount25_2mwl_core_162 = ~(input_a[21] ^ input_a[18]);
  assign popcount25_2mwl_core_164 = ~(input_a[8] & input_a[9]);
  assign popcount25_2mwl_core_167 = input_a[20] | input_a[13];
  assign popcount25_2mwl_core_169 = ~(input_a[21] ^ input_a[23]);
  assign popcount25_2mwl_core_171 = input_a[17] | input_a[6];
  assign popcount25_2mwl_core_172 = input_a[5] & input_a[10];
  assign popcount25_2mwl_core_173 = ~(input_a[24] ^ input_a[11]);
  assign popcount25_2mwl_core_174_not = ~input_a[9];
  assign popcount25_2mwl_core_175 = input_a[14] ^ input_a[4];
  assign popcount25_2mwl_core_177 = input_a[22] | input_a[13];
  assign popcount25_2mwl_core_178 = ~(input_a[16] & input_a[5]);
  assign popcount25_2mwl_core_179 = input_a[24] ^ input_a[14];
  assign popcount25_2mwl_core_181 = ~(input_a[18] ^ input_a[7]);
  assign popcount25_2mwl_core_183 = ~(input_a[4] | input_a[24]);

  assign popcount25_2mwl_out[0] = 1'b0;
  assign popcount25_2mwl_out[1] = input_a[23];
  assign popcount25_2mwl_out[2] = input_a[24];
  assign popcount25_2mwl_out[3] = 1'b1;
  assign popcount25_2mwl_out[4] = 1'b0;
endmodule