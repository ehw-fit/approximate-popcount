// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.16973
// WCE=14.0
// EP=0.856089%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_5jsl(input [26:0] input_a, output [4:0] popcount27_5jsl_out);
  wire popcount27_5jsl_core_029;
  wire popcount27_5jsl_core_031;
  wire popcount27_5jsl_core_033;
  wire popcount27_5jsl_core_034;
  wire popcount27_5jsl_core_036;
  wire popcount27_5jsl_core_037;
  wire popcount27_5jsl_core_038;
  wire popcount27_5jsl_core_041;
  wire popcount27_5jsl_core_043;
  wire popcount27_5jsl_core_044;
  wire popcount27_5jsl_core_045;
  wire popcount27_5jsl_core_046;
  wire popcount27_5jsl_core_047;
  wire popcount27_5jsl_core_048;
  wire popcount27_5jsl_core_049;
  wire popcount27_5jsl_core_050;
  wire popcount27_5jsl_core_052;
  wire popcount27_5jsl_core_053;
  wire popcount27_5jsl_core_054;
  wire popcount27_5jsl_core_056;
  wire popcount27_5jsl_core_057;
  wire popcount27_5jsl_core_058;
  wire popcount27_5jsl_core_060;
  wire popcount27_5jsl_core_061;
  wire popcount27_5jsl_core_062;
  wire popcount27_5jsl_core_064;
  wire popcount27_5jsl_core_065;
  wire popcount27_5jsl_core_066;
  wire popcount27_5jsl_core_067;
  wire popcount27_5jsl_core_071;
  wire popcount27_5jsl_core_072;
  wire popcount27_5jsl_core_073;
  wire popcount27_5jsl_core_074;
  wire popcount27_5jsl_core_075;
  wire popcount27_5jsl_core_076;
  wire popcount27_5jsl_core_077;
  wire popcount27_5jsl_core_079;
  wire popcount27_5jsl_core_080;
  wire popcount27_5jsl_core_081;
  wire popcount27_5jsl_core_083;
  wire popcount27_5jsl_core_085;
  wire popcount27_5jsl_core_088;
  wire popcount27_5jsl_core_089;
  wire popcount27_5jsl_core_090;
  wire popcount27_5jsl_core_092;
  wire popcount27_5jsl_core_093;
  wire popcount27_5jsl_core_095;
  wire popcount27_5jsl_core_102;
  wire popcount27_5jsl_core_104;
  wire popcount27_5jsl_core_106_not;
  wire popcount27_5jsl_core_107;
  wire popcount27_5jsl_core_108;
  wire popcount27_5jsl_core_111;
  wire popcount27_5jsl_core_113;
  wire popcount27_5jsl_core_114;
  wire popcount27_5jsl_core_117;
  wire popcount27_5jsl_core_118;
  wire popcount27_5jsl_core_119;
  wire popcount27_5jsl_core_120;
  wire popcount27_5jsl_core_121;
  wire popcount27_5jsl_core_123;
  wire popcount27_5jsl_core_124;
  wire popcount27_5jsl_core_126;
  wire popcount27_5jsl_core_127;
  wire popcount27_5jsl_core_129;
  wire popcount27_5jsl_core_130;
  wire popcount27_5jsl_core_132;
  wire popcount27_5jsl_core_133;
  wire popcount27_5jsl_core_134;
  wire popcount27_5jsl_core_135;
  wire popcount27_5jsl_core_136;
  wire popcount27_5jsl_core_138;
  wire popcount27_5jsl_core_139;
  wire popcount27_5jsl_core_141;
  wire popcount27_5jsl_core_143;
  wire popcount27_5jsl_core_144;
  wire popcount27_5jsl_core_146;
  wire popcount27_5jsl_core_147;
  wire popcount27_5jsl_core_148;
  wire popcount27_5jsl_core_149;
  wire popcount27_5jsl_core_151;
  wire popcount27_5jsl_core_153;
  wire popcount27_5jsl_core_155;
  wire popcount27_5jsl_core_156_not;
  wire popcount27_5jsl_core_157;
  wire popcount27_5jsl_core_158;
  wire popcount27_5jsl_core_159;
  wire popcount27_5jsl_core_161;
  wire popcount27_5jsl_core_162;
  wire popcount27_5jsl_core_163;
  wire popcount27_5jsl_core_164;
  wire popcount27_5jsl_core_165;
  wire popcount27_5jsl_core_167;
  wire popcount27_5jsl_core_170;
  wire popcount27_5jsl_core_171;
  wire popcount27_5jsl_core_172;
  wire popcount27_5jsl_core_173;
  wire popcount27_5jsl_core_174;
  wire popcount27_5jsl_core_175;
  wire popcount27_5jsl_core_176;
  wire popcount27_5jsl_core_177;
  wire popcount27_5jsl_core_178;
  wire popcount27_5jsl_core_179;
  wire popcount27_5jsl_core_180;
  wire popcount27_5jsl_core_181;
  wire popcount27_5jsl_core_182;
  wire popcount27_5jsl_core_183;
  wire popcount27_5jsl_core_184;
  wire popcount27_5jsl_core_186;
  wire popcount27_5jsl_core_188;
  wire popcount27_5jsl_core_189;
  wire popcount27_5jsl_core_190;
  wire popcount27_5jsl_core_192;
  wire popcount27_5jsl_core_194;

  assign popcount27_5jsl_core_029 = ~(input_a[22] | input_a[7]);
  assign popcount27_5jsl_core_031 = ~(input_a[13] | input_a[3]);
  assign popcount27_5jsl_core_033 = input_a[3] | input_a[8];
  assign popcount27_5jsl_core_034 = ~(input_a[14] & input_a[17]);
  assign popcount27_5jsl_core_036 = ~input_a[1];
  assign popcount27_5jsl_core_037 = ~(input_a[25] ^ input_a[13]);
  assign popcount27_5jsl_core_038 = input_a[18] | input_a[1];
  assign popcount27_5jsl_core_041 = ~input_a[21];
  assign popcount27_5jsl_core_043 = input_a[21] | input_a[0];
  assign popcount27_5jsl_core_044 = input_a[22] & input_a[6];
  assign popcount27_5jsl_core_045 = ~input_a[5];
  assign popcount27_5jsl_core_046 = ~(input_a[24] & input_a[19]);
  assign popcount27_5jsl_core_047 = ~(input_a[23] ^ input_a[10]);
  assign popcount27_5jsl_core_048 = input_a[3] | input_a[1];
  assign popcount27_5jsl_core_049 = ~(input_a[17] | input_a[23]);
  assign popcount27_5jsl_core_050 = ~(input_a[16] & input_a[16]);
  assign popcount27_5jsl_core_052 = ~(input_a[2] ^ input_a[11]);
  assign popcount27_5jsl_core_053 = input_a[4] ^ input_a[11];
  assign popcount27_5jsl_core_054 = input_a[3] ^ input_a[0];
  assign popcount27_5jsl_core_056 = ~(input_a[5] | input_a[26]);
  assign popcount27_5jsl_core_057 = ~(input_a[20] & input_a[2]);
  assign popcount27_5jsl_core_058 = ~(input_a[21] & input_a[5]);
  assign popcount27_5jsl_core_060 = input_a[18] | input_a[23];
  assign popcount27_5jsl_core_061 = ~(input_a[7] & input_a[22]);
  assign popcount27_5jsl_core_062 = input_a[15] | input_a[12];
  assign popcount27_5jsl_core_064 = ~input_a[2];
  assign popcount27_5jsl_core_065 = ~input_a[22];
  assign popcount27_5jsl_core_066 = ~(input_a[18] & input_a[7]);
  assign popcount27_5jsl_core_067 = ~(input_a[25] ^ input_a[1]);
  assign popcount27_5jsl_core_071 = input_a[15] ^ input_a[6];
  assign popcount27_5jsl_core_072 = input_a[12] & input_a[25];
  assign popcount27_5jsl_core_073 = ~input_a[11];
  assign popcount27_5jsl_core_074 = ~(input_a[20] | input_a[0]);
  assign popcount27_5jsl_core_075 = ~(input_a[24] & input_a[10]);
  assign popcount27_5jsl_core_076 = input_a[19] & input_a[21];
  assign popcount27_5jsl_core_077 = ~(input_a[18] | input_a[15]);
  assign popcount27_5jsl_core_079 = input_a[8] & input_a[19];
  assign popcount27_5jsl_core_080 = ~(input_a[23] & input_a[20]);
  assign popcount27_5jsl_core_081 = ~input_a[2];
  assign popcount27_5jsl_core_083 = input_a[24] | input_a[1];
  assign popcount27_5jsl_core_085 = input_a[16] | input_a[18];
  assign popcount27_5jsl_core_088 = input_a[10] ^ input_a[22];
  assign popcount27_5jsl_core_089 = input_a[8] ^ input_a[10];
  assign popcount27_5jsl_core_090 = ~(input_a[17] & input_a[0]);
  assign popcount27_5jsl_core_092 = input_a[5] | input_a[6];
  assign popcount27_5jsl_core_093 = input_a[24] | input_a[3];
  assign popcount27_5jsl_core_095 = ~(input_a[24] ^ input_a[19]);
  assign popcount27_5jsl_core_102 = ~(input_a[22] ^ input_a[4]);
  assign popcount27_5jsl_core_104 = ~(input_a[20] & input_a[10]);
  assign popcount27_5jsl_core_106_not = ~input_a[6];
  assign popcount27_5jsl_core_107 = input_a[17] & input_a[1];
  assign popcount27_5jsl_core_108 = ~(input_a[24] ^ input_a[11]);
  assign popcount27_5jsl_core_111 = input_a[3] | input_a[26];
  assign popcount27_5jsl_core_113 = ~input_a[12];
  assign popcount27_5jsl_core_114 = ~input_a[22];
  assign popcount27_5jsl_core_117 = ~(input_a[7] & input_a[19]);
  assign popcount27_5jsl_core_118 = input_a[19] & input_a[10];
  assign popcount27_5jsl_core_119 = ~(input_a[6] ^ input_a[11]);
  assign popcount27_5jsl_core_120 = input_a[23] ^ input_a[21];
  assign popcount27_5jsl_core_121 = ~(input_a[1] ^ input_a[23]);
  assign popcount27_5jsl_core_123 = input_a[12] | input_a[26];
  assign popcount27_5jsl_core_124 = ~(input_a[15] | input_a[7]);
  assign popcount27_5jsl_core_126 = input_a[7] & input_a[24];
  assign popcount27_5jsl_core_127 = ~(input_a[15] | input_a[20]);
  assign popcount27_5jsl_core_129 = input_a[8] | input_a[12];
  assign popcount27_5jsl_core_130 = ~input_a[18];
  assign popcount27_5jsl_core_132 = ~(input_a[24] | input_a[17]);
  assign popcount27_5jsl_core_133 = input_a[16] | input_a[18];
  assign popcount27_5jsl_core_134 = ~(input_a[9] | input_a[2]);
  assign popcount27_5jsl_core_135 = input_a[23] ^ input_a[26];
  assign popcount27_5jsl_core_136 = ~(input_a[19] ^ input_a[14]);
  assign popcount27_5jsl_core_138 = input_a[9] & input_a[22];
  assign popcount27_5jsl_core_139 = input_a[15] ^ input_a[5];
  assign popcount27_5jsl_core_141 = ~input_a[14];
  assign popcount27_5jsl_core_143 = input_a[23] & input_a[23];
  assign popcount27_5jsl_core_144 = ~(input_a[5] & input_a[23]);
  assign popcount27_5jsl_core_146 = input_a[8] ^ input_a[14];
  assign popcount27_5jsl_core_147 = input_a[13] | input_a[12];
  assign popcount27_5jsl_core_148 = ~(input_a[19] | input_a[16]);
  assign popcount27_5jsl_core_149 = ~(input_a[11] & input_a[20]);
  assign popcount27_5jsl_core_151 = ~(input_a[13] | input_a[12]);
  assign popcount27_5jsl_core_153 = ~input_a[5];
  assign popcount27_5jsl_core_155 = input_a[0] | input_a[25];
  assign popcount27_5jsl_core_156_not = ~input_a[11];
  assign popcount27_5jsl_core_157 = ~input_a[9];
  assign popcount27_5jsl_core_158 = input_a[9] | input_a[8];
  assign popcount27_5jsl_core_159 = ~(input_a[20] ^ input_a[18]);
  assign popcount27_5jsl_core_161 = ~(input_a[26] ^ input_a[14]);
  assign popcount27_5jsl_core_162 = input_a[4] & input_a[16];
  assign popcount27_5jsl_core_163 = ~input_a[1];
  assign popcount27_5jsl_core_164 = ~input_a[13];
  assign popcount27_5jsl_core_165 = input_a[18] | input_a[10];
  assign popcount27_5jsl_core_167 = input_a[2] | input_a[2];
  assign popcount27_5jsl_core_170 = ~input_a[20];
  assign popcount27_5jsl_core_171 = input_a[1] ^ input_a[11];
  assign popcount27_5jsl_core_172 = input_a[24] & input_a[6];
  assign popcount27_5jsl_core_173 = ~(input_a[5] | input_a[1]);
  assign popcount27_5jsl_core_174 = ~(input_a[8] | input_a[1]);
  assign popcount27_5jsl_core_175 = input_a[8] | input_a[26];
  assign popcount27_5jsl_core_176 = ~(input_a[15] & input_a[1]);
  assign popcount27_5jsl_core_177 = input_a[9] | input_a[12];
  assign popcount27_5jsl_core_178 = ~input_a[13];
  assign popcount27_5jsl_core_179 = ~(input_a[14] | input_a[0]);
  assign popcount27_5jsl_core_180 = ~(input_a[4] & input_a[1]);
  assign popcount27_5jsl_core_181 = input_a[25] ^ input_a[13];
  assign popcount27_5jsl_core_182 = input_a[10] & input_a[16];
  assign popcount27_5jsl_core_183 = ~(input_a[1] ^ input_a[11]);
  assign popcount27_5jsl_core_184 = ~(input_a[19] ^ input_a[13]);
  assign popcount27_5jsl_core_186 = input_a[14] ^ input_a[12];
  assign popcount27_5jsl_core_188 = input_a[21] ^ input_a[25];
  assign popcount27_5jsl_core_189 = input_a[23] ^ input_a[9];
  assign popcount27_5jsl_core_190 = ~(input_a[5] | input_a[5]);
  assign popcount27_5jsl_core_192 = input_a[22] ^ input_a[19];
  assign popcount27_5jsl_core_194 = input_a[26] & input_a[5];

  assign popcount27_5jsl_out[0] = input_a[15];
  assign popcount27_5jsl_out[1] = 1'b0;
  assign popcount27_5jsl_out[2] = 1'b1;
  assign popcount27_5jsl_out[3] = 1'b1;
  assign popcount27_5jsl_out[4] = 1'b0;
endmodule