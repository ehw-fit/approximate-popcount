// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.25652
// WCE=13.0
// EP=0.863617%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_fkj6(input [23:0] input_a, output [4:0] popcount24_fkj6_out);
  wire popcount24_fkj6_core_027;
  wire popcount24_fkj6_core_029;
  wire popcount24_fkj6_core_030;
  wire popcount24_fkj6_core_031;
  wire popcount24_fkj6_core_033;
  wire popcount24_fkj6_core_034;
  wire popcount24_fkj6_core_037;
  wire popcount24_fkj6_core_038;
  wire popcount24_fkj6_core_039;
  wire popcount24_fkj6_core_040;
  wire popcount24_fkj6_core_042;
  wire popcount24_fkj6_core_043;
  wire popcount24_fkj6_core_046;
  wire popcount24_fkj6_core_047;
  wire popcount24_fkj6_core_048;
  wire popcount24_fkj6_core_050;
  wire popcount24_fkj6_core_052;
  wire popcount24_fkj6_core_053;
  wire popcount24_fkj6_core_054;
  wire popcount24_fkj6_core_055;
  wire popcount24_fkj6_core_056;
  wire popcount24_fkj6_core_058;
  wire popcount24_fkj6_core_061;
  wire popcount24_fkj6_core_062;
  wire popcount24_fkj6_core_063;
  wire popcount24_fkj6_core_064;
  wire popcount24_fkj6_core_066;
  wire popcount24_fkj6_core_067;
  wire popcount24_fkj6_core_069;
  wire popcount24_fkj6_core_072;
  wire popcount24_fkj6_core_075;
  wire popcount24_fkj6_core_076;
  wire popcount24_fkj6_core_077;
  wire popcount24_fkj6_core_080;
  wire popcount24_fkj6_core_081;
  wire popcount24_fkj6_core_084;
  wire popcount24_fkj6_core_085;
  wire popcount24_fkj6_core_086_not;
  wire popcount24_fkj6_core_090;
  wire popcount24_fkj6_core_092;
  wire popcount24_fkj6_core_094;
  wire popcount24_fkj6_core_097;
  wire popcount24_fkj6_core_098;
  wire popcount24_fkj6_core_100;
  wire popcount24_fkj6_core_101;
  wire popcount24_fkj6_core_102;
  wire popcount24_fkj6_core_104;
  wire popcount24_fkj6_core_105;
  wire popcount24_fkj6_core_106;
  wire popcount24_fkj6_core_107;
  wire popcount24_fkj6_core_108;
  wire popcount24_fkj6_core_111;
  wire popcount24_fkj6_core_112;
  wire popcount24_fkj6_core_114;
  wire popcount24_fkj6_core_115;
  wire popcount24_fkj6_core_116;
  wire popcount24_fkj6_core_117;
  wire popcount24_fkj6_core_120;
  wire popcount24_fkj6_core_125;
  wire popcount24_fkj6_core_127;
  wire popcount24_fkj6_core_128;
  wire popcount24_fkj6_core_130;
  wire popcount24_fkj6_core_131;
  wire popcount24_fkj6_core_135;
  wire popcount24_fkj6_core_136_not;
  wire popcount24_fkj6_core_139;
  wire popcount24_fkj6_core_140_not;
  wire popcount24_fkj6_core_142;
  wire popcount24_fkj6_core_145;
  wire popcount24_fkj6_core_147;
  wire popcount24_fkj6_core_149;
  wire popcount24_fkj6_core_150;
  wire popcount24_fkj6_core_151;
  wire popcount24_fkj6_core_152;
  wire popcount24_fkj6_core_153;
  wire popcount24_fkj6_core_156;
  wire popcount24_fkj6_core_157;
  wire popcount24_fkj6_core_161;
  wire popcount24_fkj6_core_162;
  wire popcount24_fkj6_core_163;
  wire popcount24_fkj6_core_164;
  wire popcount24_fkj6_core_165;
  wire popcount24_fkj6_core_166;
  wire popcount24_fkj6_core_169;
  wire popcount24_fkj6_core_172_not;
  wire popcount24_fkj6_core_175;
  wire popcount24_fkj6_core_176;

  assign popcount24_fkj6_core_027 = ~(input_a[0] & input_a[13]);
  assign popcount24_fkj6_core_029 = ~input_a[7];
  assign popcount24_fkj6_core_030 = ~input_a[16];
  assign popcount24_fkj6_core_031 = ~(input_a[7] ^ input_a[10]);
  assign popcount24_fkj6_core_033 = ~input_a[6];
  assign popcount24_fkj6_core_034 = ~(input_a[11] | input_a[13]);
  assign popcount24_fkj6_core_037 = ~input_a[15];
  assign popcount24_fkj6_core_038 = ~input_a[11];
  assign popcount24_fkj6_core_039 = input_a[15] & input_a[6];
  assign popcount24_fkj6_core_040 = input_a[20] ^ input_a[8];
  assign popcount24_fkj6_core_042 = ~input_a[19];
  assign popcount24_fkj6_core_043 = input_a[21] & input_a[1];
  assign popcount24_fkj6_core_046 = ~(input_a[23] | input_a[15]);
  assign popcount24_fkj6_core_047 = input_a[17] | input_a[11];
  assign popcount24_fkj6_core_048 = ~input_a[15];
  assign popcount24_fkj6_core_050 = input_a[3] | input_a[10];
  assign popcount24_fkj6_core_052 = input_a[19] ^ input_a[18];
  assign popcount24_fkj6_core_053 = input_a[11] | input_a[17];
  assign popcount24_fkj6_core_054 = ~(input_a[11] & input_a[2]);
  assign popcount24_fkj6_core_055 = ~input_a[8];
  assign popcount24_fkj6_core_056 = input_a[20] | input_a[1];
  assign popcount24_fkj6_core_058 = ~input_a[7];
  assign popcount24_fkj6_core_061 = input_a[4] & input_a[7];
  assign popcount24_fkj6_core_062 = ~(input_a[5] | input_a[17]);
  assign popcount24_fkj6_core_063 = input_a[13] | input_a[11];
  assign popcount24_fkj6_core_064 = ~(input_a[22] ^ input_a[14]);
  assign popcount24_fkj6_core_066 = ~(input_a[6] & input_a[13]);
  assign popcount24_fkj6_core_067 = input_a[15] & input_a[3];
  assign popcount24_fkj6_core_069 = ~input_a[2];
  assign popcount24_fkj6_core_072 = input_a[16] | input_a[20];
  assign popcount24_fkj6_core_075 = ~(input_a[20] | input_a[5]);
  assign popcount24_fkj6_core_076 = input_a[15] | input_a[0];
  assign popcount24_fkj6_core_077 = input_a[21] ^ input_a[21];
  assign popcount24_fkj6_core_080 = input_a[4] ^ input_a[22];
  assign popcount24_fkj6_core_081 = input_a[19] | input_a[13];
  assign popcount24_fkj6_core_084 = input_a[4] | input_a[14];
  assign popcount24_fkj6_core_085 = ~input_a[15];
  assign popcount24_fkj6_core_086_not = ~input_a[4];
  assign popcount24_fkj6_core_090 = input_a[23] & input_a[13];
  assign popcount24_fkj6_core_092 = ~(input_a[14] & input_a[5]);
  assign popcount24_fkj6_core_094 = ~(input_a[7] & input_a[10]);
  assign popcount24_fkj6_core_097 = input_a[11] ^ input_a[8];
  assign popcount24_fkj6_core_098 = input_a[17] ^ input_a[0];
  assign popcount24_fkj6_core_100 = ~(input_a[16] & input_a[13]);
  assign popcount24_fkj6_core_101 = input_a[0] & input_a[15];
  assign popcount24_fkj6_core_102 = input_a[15] ^ input_a[3];
  assign popcount24_fkj6_core_104 = ~(input_a[13] | input_a[12]);
  assign popcount24_fkj6_core_105 = ~input_a[0];
  assign popcount24_fkj6_core_106 = input_a[4] & input_a[16];
  assign popcount24_fkj6_core_107 = ~(input_a[2] | input_a[12]);
  assign popcount24_fkj6_core_108 = ~input_a[20];
  assign popcount24_fkj6_core_111 = input_a[5] | input_a[0];
  assign popcount24_fkj6_core_112 = ~(input_a[4] & input_a[17]);
  assign popcount24_fkj6_core_114 = input_a[23] ^ input_a[1];
  assign popcount24_fkj6_core_115 = ~(input_a[17] ^ input_a[23]);
  assign popcount24_fkj6_core_116 = ~input_a[12];
  assign popcount24_fkj6_core_117 = input_a[22] & input_a[5];
  assign popcount24_fkj6_core_120 = ~(input_a[12] & input_a[11]);
  assign popcount24_fkj6_core_125 = ~(input_a[6] | input_a[10]);
  assign popcount24_fkj6_core_127 = ~input_a[3];
  assign popcount24_fkj6_core_128 = input_a[8] | input_a[11];
  assign popcount24_fkj6_core_130 = input_a[13] & input_a[10];
  assign popcount24_fkj6_core_131 = input_a[17] & input_a[23];
  assign popcount24_fkj6_core_135 = input_a[13] ^ input_a[20];
  assign popcount24_fkj6_core_136_not = ~input_a[6];
  assign popcount24_fkj6_core_139 = ~input_a[9];
  assign popcount24_fkj6_core_140_not = ~input_a[9];
  assign popcount24_fkj6_core_142 = ~(input_a[1] ^ input_a[0]);
  assign popcount24_fkj6_core_145 = ~(input_a[21] | input_a[18]);
  assign popcount24_fkj6_core_147 = ~(input_a[3] ^ input_a[11]);
  assign popcount24_fkj6_core_149 = ~input_a[12];
  assign popcount24_fkj6_core_150 = input_a[20] & input_a[12];
  assign popcount24_fkj6_core_151 = input_a[2] & input_a[21];
  assign popcount24_fkj6_core_152 = input_a[7] ^ input_a[11];
  assign popcount24_fkj6_core_153 = input_a[17] ^ input_a[19];
  assign popcount24_fkj6_core_156 = input_a[16] & input_a[7];
  assign popcount24_fkj6_core_157 = input_a[23] & input_a[14];
  assign popcount24_fkj6_core_161 = input_a[20] | input_a[15];
  assign popcount24_fkj6_core_162 = input_a[17] | input_a[15];
  assign popcount24_fkj6_core_163 = input_a[14] ^ input_a[15];
  assign popcount24_fkj6_core_164 = input_a[3] & input_a[12];
  assign popcount24_fkj6_core_165 = ~input_a[17];
  assign popcount24_fkj6_core_166 = ~(input_a[6] ^ input_a[2]);
  assign popcount24_fkj6_core_169 = input_a[5] & input_a[22];
  assign popcount24_fkj6_core_172_not = ~input_a[21];
  assign popcount24_fkj6_core_175 = ~(input_a[4] ^ input_a[5]);
  assign popcount24_fkj6_core_176 = ~(input_a[4] ^ input_a[18]);

  assign popcount24_fkj6_out[0] = input_a[12];
  assign popcount24_fkj6_out[1] = 1'b1;
  assign popcount24_fkj6_out[2] = 1'b0;
  assign popcount24_fkj6_out[3] = 1'b1;
  assign popcount24_fkj6_out[4] = 1'b0;
endmodule