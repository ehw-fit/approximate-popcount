// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.67128
// WCE=20.0
// EP=0.954212%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_hn6m(input [28:0] input_a, output [4:0] popcount29_hn6m_out);
  wire popcount29_hn6m_core_031;
  wire popcount29_hn6m_core_032;
  wire popcount29_hn6m_core_033;
  wire popcount29_hn6m_core_037;
  wire popcount29_hn6m_core_038;
  wire popcount29_hn6m_core_039;
  wire popcount29_hn6m_core_042;
  wire popcount29_hn6m_core_043;
  wire popcount29_hn6m_core_045;
  wire popcount29_hn6m_core_047;
  wire popcount29_hn6m_core_049;
  wire popcount29_hn6m_core_050;
  wire popcount29_hn6m_core_051;
  wire popcount29_hn6m_core_054;
  wire popcount29_hn6m_core_055;
  wire popcount29_hn6m_core_056;
  wire popcount29_hn6m_core_057;
  wire popcount29_hn6m_core_058;
  wire popcount29_hn6m_core_059;
  wire popcount29_hn6m_core_061;
  wire popcount29_hn6m_core_062;
  wire popcount29_hn6m_core_064;
  wire popcount29_hn6m_core_067;
  wire popcount29_hn6m_core_068;
  wire popcount29_hn6m_core_071;
  wire popcount29_hn6m_core_072;
  wire popcount29_hn6m_core_073;
  wire popcount29_hn6m_core_074;
  wire popcount29_hn6m_core_075;
  wire popcount29_hn6m_core_076;
  wire popcount29_hn6m_core_078;
  wire popcount29_hn6m_core_081;
  wire popcount29_hn6m_core_083;
  wire popcount29_hn6m_core_087;
  wire popcount29_hn6m_core_088;
  wire popcount29_hn6m_core_090;
  wire popcount29_hn6m_core_091;
  wire popcount29_hn6m_core_093_not;
  wire popcount29_hn6m_core_094;
  wire popcount29_hn6m_core_095;
  wire popcount29_hn6m_core_096;
  wire popcount29_hn6m_core_097;
  wire popcount29_hn6m_core_098;
  wire popcount29_hn6m_core_099;
  wire popcount29_hn6m_core_101;
  wire popcount29_hn6m_core_102;
  wire popcount29_hn6m_core_103;
  wire popcount29_hn6m_core_104;
  wire popcount29_hn6m_core_105;
  wire popcount29_hn6m_core_106;
  wire popcount29_hn6m_core_107;
  wire popcount29_hn6m_core_108;
  wire popcount29_hn6m_core_110;
  wire popcount29_hn6m_core_112;
  wire popcount29_hn6m_core_113;
  wire popcount29_hn6m_core_114;
  wire popcount29_hn6m_core_115;
  wire popcount29_hn6m_core_116;
  wire popcount29_hn6m_core_117;
  wire popcount29_hn6m_core_118;
  wire popcount29_hn6m_core_119;
  wire popcount29_hn6m_core_120;
  wire popcount29_hn6m_core_121;
  wire popcount29_hn6m_core_122;
  wire popcount29_hn6m_core_125;
  wire popcount29_hn6m_core_126;
  wire popcount29_hn6m_core_127;
  wire popcount29_hn6m_core_128;
  wire popcount29_hn6m_core_129;
  wire popcount29_hn6m_core_130;
  wire popcount29_hn6m_core_132;
  wire popcount29_hn6m_core_133;
  wire popcount29_hn6m_core_134;
  wire popcount29_hn6m_core_135;
  wire popcount29_hn6m_core_138;
  wire popcount29_hn6m_core_139;
  wire popcount29_hn6m_core_140;
  wire popcount29_hn6m_core_141;
  wire popcount29_hn6m_core_142;
  wire popcount29_hn6m_core_145;
  wire popcount29_hn6m_core_147;
  wire popcount29_hn6m_core_148;
  wire popcount29_hn6m_core_149;
  wire popcount29_hn6m_core_151;
  wire popcount29_hn6m_core_152;
  wire popcount29_hn6m_core_155;
  wire popcount29_hn6m_core_156;
  wire popcount29_hn6m_core_158;
  wire popcount29_hn6m_core_159;
  wire popcount29_hn6m_core_160;
  wire popcount29_hn6m_core_162;
  wire popcount29_hn6m_core_164;
  wire popcount29_hn6m_core_165;
  wire popcount29_hn6m_core_170;
  wire popcount29_hn6m_core_174;
  wire popcount29_hn6m_core_175;
  wire popcount29_hn6m_core_176;
  wire popcount29_hn6m_core_177;
  wire popcount29_hn6m_core_181_not;
  wire popcount29_hn6m_core_183;
  wire popcount29_hn6m_core_184;
  wire popcount29_hn6m_core_186;
  wire popcount29_hn6m_core_188;
  wire popcount29_hn6m_core_189;
  wire popcount29_hn6m_core_190;
  wire popcount29_hn6m_core_193;
  wire popcount29_hn6m_core_194;
  wire popcount29_hn6m_core_195;
  wire popcount29_hn6m_core_198;
  wire popcount29_hn6m_core_200;
  wire popcount29_hn6m_core_201;
  wire popcount29_hn6m_core_202;
  wire popcount29_hn6m_core_204;
  wire popcount29_hn6m_core_206;

  assign popcount29_hn6m_core_031 = input_a[12] ^ input_a[25];
  assign popcount29_hn6m_core_032 = ~(input_a[13] ^ input_a[4]);
  assign popcount29_hn6m_core_033 = input_a[28] ^ input_a[21];
  assign popcount29_hn6m_core_037 = input_a[12] ^ input_a[19];
  assign popcount29_hn6m_core_038 = ~(input_a[27] & input_a[10]);
  assign popcount29_hn6m_core_039 = ~(input_a[13] & input_a[14]);
  assign popcount29_hn6m_core_042 = ~input_a[25];
  assign popcount29_hn6m_core_043 = input_a[11] | input_a[4];
  assign popcount29_hn6m_core_045 = ~(input_a[8] & input_a[21]);
  assign popcount29_hn6m_core_047 = ~(input_a[1] | input_a[2]);
  assign popcount29_hn6m_core_049 = input_a[14] | input_a[7];
  assign popcount29_hn6m_core_050 = input_a[25] & input_a[21];
  assign popcount29_hn6m_core_051 = input_a[11] & input_a[11];
  assign popcount29_hn6m_core_054 = input_a[11] | input_a[13];
  assign popcount29_hn6m_core_055 = ~(input_a[18] | input_a[4]);
  assign popcount29_hn6m_core_056 = ~input_a[23];
  assign popcount29_hn6m_core_057 = ~(input_a[16] & input_a[9]);
  assign popcount29_hn6m_core_058 = ~(input_a[28] & input_a[21]);
  assign popcount29_hn6m_core_059 = input_a[5] | input_a[21];
  assign popcount29_hn6m_core_061 = input_a[2] ^ input_a[12];
  assign popcount29_hn6m_core_062 = input_a[7] | input_a[1];
  assign popcount29_hn6m_core_064 = ~(input_a[12] & input_a[12]);
  assign popcount29_hn6m_core_067 = ~(input_a[23] ^ input_a[27]);
  assign popcount29_hn6m_core_068 = ~input_a[16];
  assign popcount29_hn6m_core_071 = ~(input_a[8] ^ input_a[7]);
  assign popcount29_hn6m_core_072 = ~(input_a[10] | input_a[24]);
  assign popcount29_hn6m_core_073 = input_a[13] | input_a[13];
  assign popcount29_hn6m_core_074 = input_a[14] & input_a[1];
  assign popcount29_hn6m_core_075 = ~(input_a[4] | input_a[28]);
  assign popcount29_hn6m_core_076 = ~(input_a[11] | input_a[10]);
  assign popcount29_hn6m_core_078 = input_a[6] | input_a[13];
  assign popcount29_hn6m_core_081 = input_a[0] & input_a[18];
  assign popcount29_hn6m_core_083 = input_a[15] & input_a[16];
  assign popcount29_hn6m_core_087 = input_a[7] | input_a[14];
  assign popcount29_hn6m_core_088 = input_a[19] | input_a[21];
  assign popcount29_hn6m_core_090 = input_a[5] & input_a[5];
  assign popcount29_hn6m_core_091 = ~(input_a[23] ^ input_a[27]);
  assign popcount29_hn6m_core_093_not = ~input_a[27];
  assign popcount29_hn6m_core_094 = ~(input_a[2] & input_a[4]);
  assign popcount29_hn6m_core_095 = ~input_a[6];
  assign popcount29_hn6m_core_096 = ~(input_a[24] ^ input_a[24]);
  assign popcount29_hn6m_core_097 = ~(input_a[8] ^ input_a[11]);
  assign popcount29_hn6m_core_098 = ~(input_a[11] | input_a[28]);
  assign popcount29_hn6m_core_099 = input_a[13] ^ input_a[23];
  assign popcount29_hn6m_core_101 = ~(input_a[16] & input_a[2]);
  assign popcount29_hn6m_core_102 = ~(input_a[20] | input_a[0]);
  assign popcount29_hn6m_core_103 = input_a[12] | input_a[11];
  assign popcount29_hn6m_core_104 = input_a[21] & input_a[25];
  assign popcount29_hn6m_core_105 = input_a[17] | input_a[11];
  assign popcount29_hn6m_core_106 = input_a[10] & input_a[16];
  assign popcount29_hn6m_core_107 = ~input_a[8];
  assign popcount29_hn6m_core_108 = ~(input_a[13] | input_a[19]);
  assign popcount29_hn6m_core_110 = ~(input_a[13] ^ input_a[15]);
  assign popcount29_hn6m_core_112 = input_a[2] & input_a[28];
  assign popcount29_hn6m_core_113 = ~(input_a[4] | input_a[18]);
  assign popcount29_hn6m_core_114 = ~input_a[28];
  assign popcount29_hn6m_core_115 = input_a[12] ^ input_a[28];
  assign popcount29_hn6m_core_116 = ~(input_a[7] & input_a[0]);
  assign popcount29_hn6m_core_117 = input_a[7] ^ input_a[13];
  assign popcount29_hn6m_core_118 = input_a[11] & input_a[6];
  assign popcount29_hn6m_core_119 = input_a[4] & input_a[28];
  assign popcount29_hn6m_core_120 = input_a[23] ^ input_a[12];
  assign popcount29_hn6m_core_121 = ~(input_a[6] | input_a[19]);
  assign popcount29_hn6m_core_122 = input_a[19] ^ input_a[1];
  assign popcount29_hn6m_core_125 = ~(input_a[15] ^ input_a[14]);
  assign popcount29_hn6m_core_126 = ~(input_a[5] | input_a[22]);
  assign popcount29_hn6m_core_127 = input_a[21] ^ input_a[8];
  assign popcount29_hn6m_core_128 = ~input_a[28];
  assign popcount29_hn6m_core_129 = ~(input_a[15] | input_a[6]);
  assign popcount29_hn6m_core_130 = ~(input_a[27] ^ input_a[0]);
  assign popcount29_hn6m_core_132 = input_a[15] ^ input_a[10];
  assign popcount29_hn6m_core_133 = ~(input_a[10] & input_a[10]);
  assign popcount29_hn6m_core_134 = ~(input_a[17] ^ input_a[27]);
  assign popcount29_hn6m_core_135 = ~(input_a[15] & input_a[5]);
  assign popcount29_hn6m_core_138 = ~(input_a[26] & input_a[27]);
  assign popcount29_hn6m_core_139 = input_a[24] & input_a[6];
  assign popcount29_hn6m_core_140 = ~input_a[25];
  assign popcount29_hn6m_core_141 = ~(input_a[13] & input_a[23]);
  assign popcount29_hn6m_core_142 = ~(input_a[5] & input_a[26]);
  assign popcount29_hn6m_core_145 = ~(input_a[19] | input_a[19]);
  assign popcount29_hn6m_core_147 = ~input_a[7];
  assign popcount29_hn6m_core_148 = ~(input_a[3] | input_a[20]);
  assign popcount29_hn6m_core_149 = ~input_a[20];
  assign popcount29_hn6m_core_151 = input_a[25] & input_a[22];
  assign popcount29_hn6m_core_152 = input_a[5] & input_a[8];
  assign popcount29_hn6m_core_155 = input_a[27] ^ input_a[11];
  assign popcount29_hn6m_core_156 = input_a[22] ^ input_a[25];
  assign popcount29_hn6m_core_158 = ~input_a[0];
  assign popcount29_hn6m_core_159 = input_a[27] ^ input_a[27];
  assign popcount29_hn6m_core_160 = ~(input_a[10] ^ input_a[27]);
  assign popcount29_hn6m_core_162 = ~(input_a[21] & input_a[26]);
  assign popcount29_hn6m_core_164 = ~input_a[26];
  assign popcount29_hn6m_core_165 = ~(input_a[7] & input_a[1]);
  assign popcount29_hn6m_core_170 = input_a[1] ^ input_a[2];
  assign popcount29_hn6m_core_174 = input_a[3] ^ input_a[1];
  assign popcount29_hn6m_core_175 = ~(input_a[8] ^ input_a[7]);
  assign popcount29_hn6m_core_176 = ~(input_a[17] | input_a[3]);
  assign popcount29_hn6m_core_177 = ~(input_a[0] | input_a[10]);
  assign popcount29_hn6m_core_181_not = ~input_a[12];
  assign popcount29_hn6m_core_183 = ~input_a[6];
  assign popcount29_hn6m_core_184 = input_a[14] | input_a[23];
  assign popcount29_hn6m_core_186 = ~input_a[0];
  assign popcount29_hn6m_core_188 = ~(input_a[17] ^ input_a[6]);
  assign popcount29_hn6m_core_189 = input_a[3] ^ input_a[15];
  assign popcount29_hn6m_core_190 = input_a[8] | input_a[1];
  assign popcount29_hn6m_core_193 = input_a[8] & input_a[11];
  assign popcount29_hn6m_core_194 = input_a[5] ^ input_a[11];
  assign popcount29_hn6m_core_195 = input_a[23] ^ input_a[0];
  assign popcount29_hn6m_core_198 = input_a[28] ^ input_a[4];
  assign popcount29_hn6m_core_200 = ~(input_a[15] ^ input_a[2]);
  assign popcount29_hn6m_core_201 = ~(input_a[10] | input_a[16]);
  assign popcount29_hn6m_core_202 = ~input_a[10];
  assign popcount29_hn6m_core_204 = ~input_a[1];
  assign popcount29_hn6m_core_206 = input_a[22] | input_a[14];

  assign popcount29_hn6m_out[0] = 1'b0;
  assign popcount29_hn6m_out[1] = input_a[17];
  assign popcount29_hn6m_out[2] = input_a[21];
  assign popcount29_hn6m_out[3] = 1'b0;
  assign popcount29_hn6m_out[4] = 1'b1;
endmodule