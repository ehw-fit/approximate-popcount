// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.8579
// WCE=49.0
// EP=0.973364%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount40_8d6x(input [39:0] input_a, output [5:0] popcount40_8d6x_out);
  wire popcount40_8d6x_core_043;
  wire popcount40_8d6x_core_044;
  wire popcount40_8d6x_core_045;
  wire popcount40_8d6x_core_047;
  wire popcount40_8d6x_core_050;
  wire popcount40_8d6x_core_051;
  wire popcount40_8d6x_core_053;
  wire popcount40_8d6x_core_054;
  wire popcount40_8d6x_core_056;
  wire popcount40_8d6x_core_057;
  wire popcount40_8d6x_core_058;
  wire popcount40_8d6x_core_060;
  wire popcount40_8d6x_core_061;
  wire popcount40_8d6x_core_063;
  wire popcount40_8d6x_core_064;
  wire popcount40_8d6x_core_065;
  wire popcount40_8d6x_core_066;
  wire popcount40_8d6x_core_067;
  wire popcount40_8d6x_core_069_not;
  wire popcount40_8d6x_core_070;
  wire popcount40_8d6x_core_072;
  wire popcount40_8d6x_core_073;
  wire popcount40_8d6x_core_075;
  wire popcount40_8d6x_core_076;
  wire popcount40_8d6x_core_077;
  wire popcount40_8d6x_core_079;
  wire popcount40_8d6x_core_080;
  wire popcount40_8d6x_core_081;
  wire popcount40_8d6x_core_082;
  wire popcount40_8d6x_core_084;
  wire popcount40_8d6x_core_085;
  wire popcount40_8d6x_core_086;
  wire popcount40_8d6x_core_088;
  wire popcount40_8d6x_core_089;
  wire popcount40_8d6x_core_090;
  wire popcount40_8d6x_core_091;
  wire popcount40_8d6x_core_092_not;
  wire popcount40_8d6x_core_094;
  wire popcount40_8d6x_core_095;
  wire popcount40_8d6x_core_098;
  wire popcount40_8d6x_core_100;
  wire popcount40_8d6x_core_101;
  wire popcount40_8d6x_core_102;
  wire popcount40_8d6x_core_103;
  wire popcount40_8d6x_core_106;
  wire popcount40_8d6x_core_107;
  wire popcount40_8d6x_core_108;
  wire popcount40_8d6x_core_109;
  wire popcount40_8d6x_core_110;
  wire popcount40_8d6x_core_111;
  wire popcount40_8d6x_core_113;
  wire popcount40_8d6x_core_115;
  wire popcount40_8d6x_core_117;
  wire popcount40_8d6x_core_119;
  wire popcount40_8d6x_core_120;
  wire popcount40_8d6x_core_121;
  wire popcount40_8d6x_core_122;
  wire popcount40_8d6x_core_124;
  wire popcount40_8d6x_core_125;
  wire popcount40_8d6x_core_126;
  wire popcount40_8d6x_core_129;
  wire popcount40_8d6x_core_130;
  wire popcount40_8d6x_core_132;
  wire popcount40_8d6x_core_136;
  wire popcount40_8d6x_core_137;
  wire popcount40_8d6x_core_139;
  wire popcount40_8d6x_core_140;
  wire popcount40_8d6x_core_143;
  wire popcount40_8d6x_core_145;
  wire popcount40_8d6x_core_146;
  wire popcount40_8d6x_core_147;
  wire popcount40_8d6x_core_148;
  wire popcount40_8d6x_core_150;
  wire popcount40_8d6x_core_151_not;
  wire popcount40_8d6x_core_153;
  wire popcount40_8d6x_core_155;
  wire popcount40_8d6x_core_156;
  wire popcount40_8d6x_core_157;
  wire popcount40_8d6x_core_158;
  wire popcount40_8d6x_core_159;
  wire popcount40_8d6x_core_160;
  wire popcount40_8d6x_core_161;
  wire popcount40_8d6x_core_162;
  wire popcount40_8d6x_core_163;
  wire popcount40_8d6x_core_164;
  wire popcount40_8d6x_core_165;
  wire popcount40_8d6x_core_166;
  wire popcount40_8d6x_core_167;
  wire popcount40_8d6x_core_168;
  wire popcount40_8d6x_core_169;
  wire popcount40_8d6x_core_173;
  wire popcount40_8d6x_core_175_not;
  wire popcount40_8d6x_core_176;
  wire popcount40_8d6x_core_177;
  wire popcount40_8d6x_core_178;
  wire popcount40_8d6x_core_179;
  wire popcount40_8d6x_core_180;
  wire popcount40_8d6x_core_181;
  wire popcount40_8d6x_core_182;
  wire popcount40_8d6x_core_183;
  wire popcount40_8d6x_core_185;
  wire popcount40_8d6x_core_186;
  wire popcount40_8d6x_core_187;
  wire popcount40_8d6x_core_190;
  wire popcount40_8d6x_core_191;
  wire popcount40_8d6x_core_192;
  wire popcount40_8d6x_core_195;
  wire popcount40_8d6x_core_196;
  wire popcount40_8d6x_core_197;
  wire popcount40_8d6x_core_198;
  wire popcount40_8d6x_core_199;
  wire popcount40_8d6x_core_200;
  wire popcount40_8d6x_core_201;
  wire popcount40_8d6x_core_202;
  wire popcount40_8d6x_core_203;
  wire popcount40_8d6x_core_204;
  wire popcount40_8d6x_core_205;
  wire popcount40_8d6x_core_207;
  wire popcount40_8d6x_core_208;
  wire popcount40_8d6x_core_209;
  wire popcount40_8d6x_core_210;
  wire popcount40_8d6x_core_211;
  wire popcount40_8d6x_core_212;
  wire popcount40_8d6x_core_215;
  wire popcount40_8d6x_core_217;
  wire popcount40_8d6x_core_218;
  wire popcount40_8d6x_core_220;
  wire popcount40_8d6x_core_225;
  wire popcount40_8d6x_core_226;
  wire popcount40_8d6x_core_227_not;
  wire popcount40_8d6x_core_228;
  wire popcount40_8d6x_core_229;
  wire popcount40_8d6x_core_230;
  wire popcount40_8d6x_core_231;
  wire popcount40_8d6x_core_233;
  wire popcount40_8d6x_core_234;
  wire popcount40_8d6x_core_235;
  wire popcount40_8d6x_core_236;
  wire popcount40_8d6x_core_237;
  wire popcount40_8d6x_core_239;
  wire popcount40_8d6x_core_240;
  wire popcount40_8d6x_core_241_not;
  wire popcount40_8d6x_core_242;
  wire popcount40_8d6x_core_244;
  wire popcount40_8d6x_core_246;
  wire popcount40_8d6x_core_247;
  wire popcount40_8d6x_core_249;
  wire popcount40_8d6x_core_251;
  wire popcount40_8d6x_core_252;
  wire popcount40_8d6x_core_253;
  wire popcount40_8d6x_core_255;
  wire popcount40_8d6x_core_258;
  wire popcount40_8d6x_core_259;
  wire popcount40_8d6x_core_261;
  wire popcount40_8d6x_core_262;
  wire popcount40_8d6x_core_265;
  wire popcount40_8d6x_core_268;
  wire popcount40_8d6x_core_269;
  wire popcount40_8d6x_core_271;
  wire popcount40_8d6x_core_272;
  wire popcount40_8d6x_core_274;
  wire popcount40_8d6x_core_276;
  wire popcount40_8d6x_core_277;
  wire popcount40_8d6x_core_279;
  wire popcount40_8d6x_core_280;
  wire popcount40_8d6x_core_281;
  wire popcount40_8d6x_core_282;
  wire popcount40_8d6x_core_284;
  wire popcount40_8d6x_core_287;
  wire popcount40_8d6x_core_288;
  wire popcount40_8d6x_core_289;
  wire popcount40_8d6x_core_290;
  wire popcount40_8d6x_core_291;
  wire popcount40_8d6x_core_293_not;
  wire popcount40_8d6x_core_295;
  wire popcount40_8d6x_core_297;
  wire popcount40_8d6x_core_299;
  wire popcount40_8d6x_core_300;
  wire popcount40_8d6x_core_302;
  wire popcount40_8d6x_core_304;
  wire popcount40_8d6x_core_305;
  wire popcount40_8d6x_core_306;
  wire popcount40_8d6x_core_309;
  wire popcount40_8d6x_core_310;
  wire popcount40_8d6x_core_311;
  wire popcount40_8d6x_core_312;
  wire popcount40_8d6x_core_313_not;
  wire popcount40_8d6x_core_314;
  wire popcount40_8d6x_core_315;

  assign popcount40_8d6x_core_043 = input_a[36] & input_a[37];
  assign popcount40_8d6x_core_044 = input_a[38] & input_a[2];
  assign popcount40_8d6x_core_045 = ~(input_a[12] ^ input_a[2]);
  assign popcount40_8d6x_core_047 = ~(input_a[32] & input_a[36]);
  assign popcount40_8d6x_core_050 = ~(input_a[4] ^ input_a[18]);
  assign popcount40_8d6x_core_051 = ~(input_a[8] ^ input_a[2]);
  assign popcount40_8d6x_core_053 = input_a[0] ^ input_a[10];
  assign popcount40_8d6x_core_054 = input_a[2] & input_a[26];
  assign popcount40_8d6x_core_056 = ~input_a[7];
  assign popcount40_8d6x_core_057 = input_a[8] | input_a[38];
  assign popcount40_8d6x_core_058 = input_a[4] | input_a[26];
  assign popcount40_8d6x_core_060 = input_a[35] | input_a[35];
  assign popcount40_8d6x_core_061 = ~(input_a[26] ^ input_a[38]);
  assign popcount40_8d6x_core_063 = ~(input_a[4] ^ input_a[39]);
  assign popcount40_8d6x_core_064 = input_a[26] | input_a[25];
  assign popcount40_8d6x_core_065 = ~input_a[22];
  assign popcount40_8d6x_core_066 = ~(input_a[22] & input_a[37]);
  assign popcount40_8d6x_core_067 = ~input_a[27];
  assign popcount40_8d6x_core_069_not = ~input_a[32];
  assign popcount40_8d6x_core_070 = input_a[4] & input_a[36];
  assign popcount40_8d6x_core_072 = ~(input_a[26] ^ input_a[16]);
  assign popcount40_8d6x_core_073 = input_a[18] ^ input_a[12];
  assign popcount40_8d6x_core_075 = input_a[4] | input_a[18];
  assign popcount40_8d6x_core_076 = ~(input_a[25] ^ input_a[0]);
  assign popcount40_8d6x_core_077 = input_a[34] ^ input_a[9];
  assign popcount40_8d6x_core_079 = ~(input_a[23] & input_a[36]);
  assign popcount40_8d6x_core_080 = ~(input_a[16] ^ input_a[0]);
  assign popcount40_8d6x_core_081 = input_a[12] & input_a[16];
  assign popcount40_8d6x_core_082 = ~(input_a[19] ^ input_a[17]);
  assign popcount40_8d6x_core_084 = ~(input_a[37] ^ input_a[26]);
  assign popcount40_8d6x_core_085 = input_a[0] | input_a[1];
  assign popcount40_8d6x_core_086 = ~input_a[31];
  assign popcount40_8d6x_core_088 = ~(input_a[23] ^ input_a[30]);
  assign popcount40_8d6x_core_089 = input_a[21] & input_a[18];
  assign popcount40_8d6x_core_090 = input_a[1] ^ input_a[25];
  assign popcount40_8d6x_core_091 = input_a[39] ^ input_a[12];
  assign popcount40_8d6x_core_092_not = ~input_a[27];
  assign popcount40_8d6x_core_094 = ~input_a[30];
  assign popcount40_8d6x_core_095 = ~(input_a[33] | input_a[28]);
  assign popcount40_8d6x_core_098 = ~(input_a[24] & input_a[9]);
  assign popcount40_8d6x_core_100 = input_a[39] ^ input_a[33];
  assign popcount40_8d6x_core_101 = ~(input_a[25] & input_a[16]);
  assign popcount40_8d6x_core_102 = input_a[7] ^ input_a[4];
  assign popcount40_8d6x_core_103 = ~(input_a[31] & input_a[7]);
  assign popcount40_8d6x_core_106 = ~(input_a[9] ^ input_a[6]);
  assign popcount40_8d6x_core_107 = ~input_a[22];
  assign popcount40_8d6x_core_108 = input_a[15] | input_a[6];
  assign popcount40_8d6x_core_109 = input_a[10] | input_a[1];
  assign popcount40_8d6x_core_110 = input_a[2] | input_a[34];
  assign popcount40_8d6x_core_111 = ~(input_a[5] ^ input_a[17]);
  assign popcount40_8d6x_core_113 = ~input_a[35];
  assign popcount40_8d6x_core_115 = ~(input_a[4] | input_a[3]);
  assign popcount40_8d6x_core_117 = ~input_a[33];
  assign popcount40_8d6x_core_119 = input_a[38] & input_a[3];
  assign popcount40_8d6x_core_120 = input_a[33] ^ input_a[18];
  assign popcount40_8d6x_core_121 = input_a[7] ^ input_a[0];
  assign popcount40_8d6x_core_122 = ~(input_a[35] ^ input_a[30]);
  assign popcount40_8d6x_core_124 = input_a[22] | input_a[35];
  assign popcount40_8d6x_core_125 = ~input_a[22];
  assign popcount40_8d6x_core_126 = ~input_a[3];
  assign popcount40_8d6x_core_129 = input_a[32] | input_a[31];
  assign popcount40_8d6x_core_130 = ~(input_a[26] & input_a[5]);
  assign popcount40_8d6x_core_132 = ~input_a[29];
  assign popcount40_8d6x_core_136 = input_a[39] ^ input_a[39];
  assign popcount40_8d6x_core_137 = input_a[15] & input_a[10];
  assign popcount40_8d6x_core_139 = input_a[38] & input_a[28];
  assign popcount40_8d6x_core_140 = ~input_a[31];
  assign popcount40_8d6x_core_143 = ~(input_a[1] | input_a[7]);
  assign popcount40_8d6x_core_145 = ~(input_a[20] & input_a[1]);
  assign popcount40_8d6x_core_146 = input_a[19] & input_a[36];
  assign popcount40_8d6x_core_147 = ~(input_a[27] & input_a[20]);
  assign popcount40_8d6x_core_148 = input_a[23] ^ input_a[9];
  assign popcount40_8d6x_core_150 = input_a[11] ^ input_a[36];
  assign popcount40_8d6x_core_151_not = ~input_a[5];
  assign popcount40_8d6x_core_153 = input_a[29] | input_a[18];
  assign popcount40_8d6x_core_155 = input_a[3] ^ input_a[33];
  assign popcount40_8d6x_core_156 = ~(input_a[16] & input_a[34]);
  assign popcount40_8d6x_core_157 = ~(input_a[39] ^ input_a[9]);
  assign popcount40_8d6x_core_158 = input_a[29] & input_a[13];
  assign popcount40_8d6x_core_159 = input_a[1] & input_a[25];
  assign popcount40_8d6x_core_160 = ~(input_a[33] | input_a[16]);
  assign popcount40_8d6x_core_161 = ~(input_a[6] & input_a[10]);
  assign popcount40_8d6x_core_162 = input_a[31] ^ input_a[32];
  assign popcount40_8d6x_core_163 = input_a[38] | input_a[20];
  assign popcount40_8d6x_core_164 = input_a[34] ^ input_a[22];
  assign popcount40_8d6x_core_165 = input_a[20] | input_a[39];
  assign popcount40_8d6x_core_166 = ~(input_a[21] ^ input_a[28]);
  assign popcount40_8d6x_core_167 = ~(input_a[1] | input_a[34]);
  assign popcount40_8d6x_core_168 = ~(input_a[12] | input_a[21]);
  assign popcount40_8d6x_core_169 = input_a[4] ^ input_a[37];
  assign popcount40_8d6x_core_173 = ~input_a[36];
  assign popcount40_8d6x_core_175_not = ~input_a[19];
  assign popcount40_8d6x_core_176 = ~(input_a[0] & input_a[32]);
  assign popcount40_8d6x_core_177 = ~(input_a[1] | input_a[22]);
  assign popcount40_8d6x_core_178 = ~input_a[25];
  assign popcount40_8d6x_core_179 = input_a[27] ^ input_a[8];
  assign popcount40_8d6x_core_180 = input_a[27] & input_a[21];
  assign popcount40_8d6x_core_181 = input_a[7] & input_a[6];
  assign popcount40_8d6x_core_182 = input_a[11] | input_a[2];
  assign popcount40_8d6x_core_183 = ~(input_a[3] & input_a[0]);
  assign popcount40_8d6x_core_185 = ~input_a[5];
  assign popcount40_8d6x_core_186 = input_a[3] | input_a[38];
  assign popcount40_8d6x_core_187 = input_a[29] | input_a[26];
  assign popcount40_8d6x_core_190 = input_a[11] | input_a[36];
  assign popcount40_8d6x_core_191 = input_a[8] | input_a[13];
  assign popcount40_8d6x_core_192 = input_a[8] ^ input_a[6];
  assign popcount40_8d6x_core_195 = ~input_a[19];
  assign popcount40_8d6x_core_196 = ~(input_a[21] & input_a[24]);
  assign popcount40_8d6x_core_197 = ~(input_a[31] & input_a[31]);
  assign popcount40_8d6x_core_198 = ~(input_a[17] | input_a[37]);
  assign popcount40_8d6x_core_199 = ~(input_a[11] | input_a[8]);
  assign popcount40_8d6x_core_200 = input_a[18] ^ input_a[32];
  assign popcount40_8d6x_core_201 = ~input_a[14];
  assign popcount40_8d6x_core_202 = ~(input_a[12] ^ input_a[24]);
  assign popcount40_8d6x_core_203 = ~(input_a[16] & input_a[37]);
  assign popcount40_8d6x_core_204 = ~input_a[22];
  assign popcount40_8d6x_core_205 = ~(input_a[8] & input_a[33]);
  assign popcount40_8d6x_core_207 = ~(input_a[31] | input_a[4]);
  assign popcount40_8d6x_core_208 = input_a[10] | input_a[2];
  assign popcount40_8d6x_core_209 = ~(input_a[21] ^ input_a[25]);
  assign popcount40_8d6x_core_210 = input_a[3] | input_a[36];
  assign popcount40_8d6x_core_211 = ~(input_a[14] | input_a[0]);
  assign popcount40_8d6x_core_212 = input_a[1] & input_a[11];
  assign popcount40_8d6x_core_215 = ~(input_a[9] | input_a[23]);
  assign popcount40_8d6x_core_217 = ~(input_a[26] | input_a[19]);
  assign popcount40_8d6x_core_218 = ~(input_a[36] & input_a[0]);
  assign popcount40_8d6x_core_220 = ~(input_a[1] & input_a[1]);
  assign popcount40_8d6x_core_225 = ~(input_a[20] ^ input_a[26]);
  assign popcount40_8d6x_core_226 = input_a[23] & input_a[4];
  assign popcount40_8d6x_core_227_not = ~input_a[8];
  assign popcount40_8d6x_core_228 = ~(input_a[27] & input_a[17]);
  assign popcount40_8d6x_core_229 = input_a[6] ^ input_a[20];
  assign popcount40_8d6x_core_230 = ~(input_a[19] & input_a[12]);
  assign popcount40_8d6x_core_231 = ~(input_a[15] ^ input_a[22]);
  assign popcount40_8d6x_core_233 = ~(input_a[33] & input_a[20]);
  assign popcount40_8d6x_core_234 = ~input_a[11];
  assign popcount40_8d6x_core_235 = ~(input_a[39] | input_a[6]);
  assign popcount40_8d6x_core_236 = input_a[16] & input_a[32];
  assign popcount40_8d6x_core_237 = ~(input_a[36] ^ input_a[16]);
  assign popcount40_8d6x_core_239 = input_a[25] ^ input_a[36];
  assign popcount40_8d6x_core_240 = input_a[15] ^ input_a[18];
  assign popcount40_8d6x_core_241_not = ~input_a[36];
  assign popcount40_8d6x_core_242 = ~(input_a[9] | input_a[7]);
  assign popcount40_8d6x_core_244 = input_a[27] & input_a[34];
  assign popcount40_8d6x_core_246 = input_a[38] | input_a[22];
  assign popcount40_8d6x_core_247 = ~(input_a[14] | input_a[33]);
  assign popcount40_8d6x_core_249 = ~(input_a[25] & input_a[26]);
  assign popcount40_8d6x_core_251 = ~(input_a[6] ^ input_a[21]);
  assign popcount40_8d6x_core_252 = ~(input_a[23] & input_a[20]);
  assign popcount40_8d6x_core_253 = ~(input_a[31] | input_a[13]);
  assign popcount40_8d6x_core_255 = ~(input_a[11] ^ input_a[21]);
  assign popcount40_8d6x_core_258 = ~input_a[26];
  assign popcount40_8d6x_core_259 = input_a[23] ^ input_a[7];
  assign popcount40_8d6x_core_261 = input_a[36] & input_a[8];
  assign popcount40_8d6x_core_262 = ~(input_a[27] & input_a[19]);
  assign popcount40_8d6x_core_265 = ~(input_a[35] ^ input_a[37]);
  assign popcount40_8d6x_core_268 = input_a[0] ^ input_a[15];
  assign popcount40_8d6x_core_269 = ~input_a[30];
  assign popcount40_8d6x_core_271 = ~(input_a[9] & input_a[13]);
  assign popcount40_8d6x_core_272 = ~(input_a[36] ^ input_a[8]);
  assign popcount40_8d6x_core_274 = input_a[37] ^ input_a[26];
  assign popcount40_8d6x_core_276 = ~(input_a[26] & input_a[28]);
  assign popcount40_8d6x_core_277 = ~(input_a[21] ^ input_a[2]);
  assign popcount40_8d6x_core_279 = ~(input_a[8] | input_a[2]);
  assign popcount40_8d6x_core_280 = ~(input_a[8] ^ input_a[28]);
  assign popcount40_8d6x_core_281 = ~(input_a[35] ^ input_a[17]);
  assign popcount40_8d6x_core_282 = ~input_a[33];
  assign popcount40_8d6x_core_284 = input_a[35] & input_a[39];
  assign popcount40_8d6x_core_287 = input_a[30] | input_a[19];
  assign popcount40_8d6x_core_288 = input_a[39] ^ input_a[15];
  assign popcount40_8d6x_core_289 = input_a[13] & input_a[37];
  assign popcount40_8d6x_core_290 = ~(input_a[39] & input_a[13]);
  assign popcount40_8d6x_core_291 = input_a[4] ^ input_a[10];
  assign popcount40_8d6x_core_293_not = ~input_a[9];
  assign popcount40_8d6x_core_295 = ~(input_a[16] | input_a[12]);
  assign popcount40_8d6x_core_297 = ~input_a[33];
  assign popcount40_8d6x_core_299 = ~input_a[15];
  assign popcount40_8d6x_core_300 = ~(input_a[31] | input_a[27]);
  assign popcount40_8d6x_core_302 = ~(input_a[19] ^ input_a[13]);
  assign popcount40_8d6x_core_304 = ~(input_a[2] | input_a[33]);
  assign popcount40_8d6x_core_305 = ~(input_a[30] ^ input_a[10]);
  assign popcount40_8d6x_core_306 = ~input_a[26];
  assign popcount40_8d6x_core_309 = ~(input_a[4] & input_a[6]);
  assign popcount40_8d6x_core_310 = ~(input_a[6] ^ input_a[19]);
  assign popcount40_8d6x_core_311 = input_a[16] | input_a[38];
  assign popcount40_8d6x_core_312 = input_a[15] ^ input_a[1];
  assign popcount40_8d6x_core_313_not = ~input_a[19];
  assign popcount40_8d6x_core_314 = input_a[16] | input_a[4];
  assign popcount40_8d6x_core_315 = input_a[29] ^ input_a[35];

  assign popcount40_8d6x_out[0] = input_a[7];
  assign popcount40_8d6x_out[1] = 1'b0;
  assign popcount40_8d6x_out[2] = input_a[23];
  assign popcount40_8d6x_out[3] = 1'b0;
  assign popcount40_8d6x_out[4] = input_a[32];
  assign popcount40_8d6x_out[5] = input_a[4];
endmodule