// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.5191
// WCE=17.0
// EP=0.876515%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount33_oce2(input [32:0] input_a, output [5:0] popcount33_oce2_out);
  wire popcount33_oce2_core_035;
  wire popcount33_oce2_core_036;
  wire popcount33_oce2_core_037;
  wire popcount33_oce2_core_040;
  wire popcount33_oce2_core_041;
  wire popcount33_oce2_core_042_not;
  wire popcount33_oce2_core_043;
  wire popcount33_oce2_core_045;
  wire popcount33_oce2_core_047;
  wire popcount33_oce2_core_050;
  wire popcount33_oce2_core_051;
  wire popcount33_oce2_core_052;
  wire popcount33_oce2_core_054;
  wire popcount33_oce2_core_055;
  wire popcount33_oce2_core_057;
  wire popcount33_oce2_core_058;
  wire popcount33_oce2_core_059;
  wire popcount33_oce2_core_060;
  wire popcount33_oce2_core_061;
  wire popcount33_oce2_core_062;
  wire popcount33_oce2_core_066;
  wire popcount33_oce2_core_068;
  wire popcount33_oce2_core_070;
  wire popcount33_oce2_core_071;
  wire popcount33_oce2_core_073;
  wire popcount33_oce2_core_075;
  wire popcount33_oce2_core_076;
  wire popcount33_oce2_core_080;
  wire popcount33_oce2_core_082;
  wire popcount33_oce2_core_083;
  wire popcount33_oce2_core_084;
  wire popcount33_oce2_core_085;
  wire popcount33_oce2_core_086;
  wire popcount33_oce2_core_087;
  wire popcount33_oce2_core_089;
  wire popcount33_oce2_core_091;
  wire popcount33_oce2_core_092;
  wire popcount33_oce2_core_093;
  wire popcount33_oce2_core_094;
  wire popcount33_oce2_core_096;
  wire popcount33_oce2_core_097;
  wire popcount33_oce2_core_098;
  wire popcount33_oce2_core_099;
  wire popcount33_oce2_core_100;
  wire popcount33_oce2_core_101;
  wire popcount33_oce2_core_102;
  wire popcount33_oce2_core_103;
  wire popcount33_oce2_core_104;
  wire popcount33_oce2_core_105;
  wire popcount33_oce2_core_106;
  wire popcount33_oce2_core_107;
  wire popcount33_oce2_core_108;
  wire popcount33_oce2_core_109;
  wire popcount33_oce2_core_110;
  wire popcount33_oce2_core_112;
  wire popcount33_oce2_core_113;
  wire popcount33_oce2_core_114;
  wire popcount33_oce2_core_115;
  wire popcount33_oce2_core_117;
  wire popcount33_oce2_core_118;
  wire popcount33_oce2_core_119;
  wire popcount33_oce2_core_121;
  wire popcount33_oce2_core_123;
  wire popcount33_oce2_core_125;
  wire popcount33_oce2_core_127;
  wire popcount33_oce2_core_129;
  wire popcount33_oce2_core_132;
  wire popcount33_oce2_core_133;
  wire popcount33_oce2_core_134;
  wire popcount33_oce2_core_135;
  wire popcount33_oce2_core_141;
  wire popcount33_oce2_core_142;
  wire popcount33_oce2_core_143;
  wire popcount33_oce2_core_144;
  wire popcount33_oce2_core_145;
  wire popcount33_oce2_core_146;
  wire popcount33_oce2_core_148;
  wire popcount33_oce2_core_149;
  wire popcount33_oce2_core_150;
  wire popcount33_oce2_core_151;
  wire popcount33_oce2_core_152;
  wire popcount33_oce2_core_154;
  wire popcount33_oce2_core_156;
  wire popcount33_oce2_core_158;
  wire popcount33_oce2_core_159;
  wire popcount33_oce2_core_163;
  wire popcount33_oce2_core_164;
  wire popcount33_oce2_core_165;
  wire popcount33_oce2_core_167;
  wire popcount33_oce2_core_171;
  wire popcount33_oce2_core_172;
  wire popcount33_oce2_core_173;
  wire popcount33_oce2_core_174;
  wire popcount33_oce2_core_176;
  wire popcount33_oce2_core_177;
  wire popcount33_oce2_core_178;
  wire popcount33_oce2_core_180;
  wire popcount33_oce2_core_181;
  wire popcount33_oce2_core_182;
  wire popcount33_oce2_core_183;
  wire popcount33_oce2_core_185;
  wire popcount33_oce2_core_186_not;
  wire popcount33_oce2_core_187;
  wire popcount33_oce2_core_189;
  wire popcount33_oce2_core_190;
  wire popcount33_oce2_core_191;
  wire popcount33_oce2_core_192;
  wire popcount33_oce2_core_193;
  wire popcount33_oce2_core_194;
  wire popcount33_oce2_core_196;
  wire popcount33_oce2_core_197;
  wire popcount33_oce2_core_198;
  wire popcount33_oce2_core_199;
  wire popcount33_oce2_core_202;
  wire popcount33_oce2_core_203;
  wire popcount33_oce2_core_205;
  wire popcount33_oce2_core_206;
  wire popcount33_oce2_core_210;
  wire popcount33_oce2_core_211;
  wire popcount33_oce2_core_213;
  wire popcount33_oce2_core_214_not;
  wire popcount33_oce2_core_215;
  wire popcount33_oce2_core_216;
  wire popcount33_oce2_core_217;
  wire popcount33_oce2_core_218;
  wire popcount33_oce2_core_220;
  wire popcount33_oce2_core_223_not;
  wire popcount33_oce2_core_224;
  wire popcount33_oce2_core_225;
  wire popcount33_oce2_core_227;
  wire popcount33_oce2_core_228;
  wire popcount33_oce2_core_229;
  wire popcount33_oce2_core_230;
  wire popcount33_oce2_core_231;
  wire popcount33_oce2_core_234;
  wire popcount33_oce2_core_235;
  wire popcount33_oce2_core_236;
  wire popcount33_oce2_core_237;

  assign popcount33_oce2_core_035 = input_a[4] ^ input_a[4];
  assign popcount33_oce2_core_036 = input_a[19] & input_a[2];
  assign popcount33_oce2_core_037 = input_a[2] ^ input_a[10];
  assign popcount33_oce2_core_040 = ~(input_a[22] | input_a[25]);
  assign popcount33_oce2_core_041 = input_a[27] | input_a[25];
  assign popcount33_oce2_core_042_not = ~input_a[3];
  assign popcount33_oce2_core_043 = input_a[20] | input_a[23];
  assign popcount33_oce2_core_045 = ~input_a[2];
  assign popcount33_oce2_core_047 = ~(input_a[14] ^ input_a[18]);
  assign popcount33_oce2_core_050 = input_a[30] ^ input_a[12];
  assign popcount33_oce2_core_051 = ~(input_a[6] & input_a[21]);
  assign popcount33_oce2_core_052 = input_a[17] ^ input_a[22];
  assign popcount33_oce2_core_054 = input_a[14] & input_a[12];
  assign popcount33_oce2_core_055 = input_a[5] ^ input_a[30];
  assign popcount33_oce2_core_057 = ~(input_a[21] & input_a[29]);
  assign popcount33_oce2_core_058 = input_a[11] ^ input_a[10];
  assign popcount33_oce2_core_059 = ~(input_a[26] | input_a[19]);
  assign popcount33_oce2_core_060 = input_a[19] | input_a[18];
  assign popcount33_oce2_core_061 = ~input_a[6];
  assign popcount33_oce2_core_062 = input_a[17] & input_a[28];
  assign popcount33_oce2_core_066 = input_a[11] & input_a[27];
  assign popcount33_oce2_core_068 = ~(input_a[23] & input_a[31]);
  assign popcount33_oce2_core_070 = ~(input_a[32] ^ input_a[6]);
  assign popcount33_oce2_core_071 = ~input_a[26];
  assign popcount33_oce2_core_073 = ~(input_a[21] | input_a[21]);
  assign popcount33_oce2_core_075 = input_a[32] | input_a[19];
  assign popcount33_oce2_core_076 = ~(input_a[8] & input_a[21]);
  assign popcount33_oce2_core_080 = ~(input_a[12] & input_a[25]);
  assign popcount33_oce2_core_082 = input_a[23] | input_a[6];
  assign popcount33_oce2_core_083 = input_a[15] & input_a[12];
  assign popcount33_oce2_core_084 = ~(input_a[31] & input_a[8]);
  assign popcount33_oce2_core_085 = input_a[4] ^ input_a[29];
  assign popcount33_oce2_core_086 = ~(input_a[13] ^ input_a[2]);
  assign popcount33_oce2_core_087 = ~(input_a[23] | input_a[32]);
  assign popcount33_oce2_core_089 = input_a[3] | input_a[21];
  assign popcount33_oce2_core_091 = ~(input_a[3] ^ input_a[32]);
  assign popcount33_oce2_core_092 = input_a[10] & input_a[1];
  assign popcount33_oce2_core_093 = input_a[4] & input_a[29];
  assign popcount33_oce2_core_094 = input_a[19] | input_a[17];
  assign popcount33_oce2_core_096 = input_a[26] & input_a[9];
  assign popcount33_oce2_core_097 = ~(input_a[25] & input_a[21]);
  assign popcount33_oce2_core_098 = input_a[28] ^ input_a[12];
  assign popcount33_oce2_core_099 = input_a[27] & input_a[21];
  assign popcount33_oce2_core_100 = ~input_a[19];
  assign popcount33_oce2_core_101 = ~(input_a[24] | input_a[20]);
  assign popcount33_oce2_core_102 = input_a[28] | input_a[6];
  assign popcount33_oce2_core_103 = ~(input_a[6] ^ input_a[7]);
  assign popcount33_oce2_core_104 = input_a[32] | input_a[14];
  assign popcount33_oce2_core_105 = input_a[7] | input_a[20];
  assign popcount33_oce2_core_106 = input_a[27] ^ input_a[30];
  assign popcount33_oce2_core_107 = ~(input_a[0] & input_a[3]);
  assign popcount33_oce2_core_108 = input_a[9] & input_a[2];
  assign popcount33_oce2_core_109 = input_a[15] & input_a[8];
  assign popcount33_oce2_core_110 = ~input_a[0];
  assign popcount33_oce2_core_112 = ~(input_a[29] | input_a[1]);
  assign popcount33_oce2_core_113 = input_a[22] | input_a[19];
  assign popcount33_oce2_core_114 = ~(input_a[23] & input_a[7]);
  assign popcount33_oce2_core_115 = ~(input_a[7] | input_a[22]);
  assign popcount33_oce2_core_117 = input_a[0] | input_a[4];
  assign popcount33_oce2_core_118 = ~input_a[23];
  assign popcount33_oce2_core_119 = ~input_a[26];
  assign popcount33_oce2_core_121 = input_a[5] ^ input_a[2];
  assign popcount33_oce2_core_123 = ~(input_a[0] | input_a[6]);
  assign popcount33_oce2_core_125 = ~(input_a[25] | input_a[24]);
  assign popcount33_oce2_core_127 = ~input_a[16];
  assign popcount33_oce2_core_129 = ~(input_a[1] | input_a[32]);
  assign popcount33_oce2_core_132 = ~(input_a[16] | input_a[23]);
  assign popcount33_oce2_core_133 = input_a[7] ^ input_a[12];
  assign popcount33_oce2_core_134 = ~(input_a[16] ^ input_a[19]);
  assign popcount33_oce2_core_135 = input_a[19] ^ input_a[29];
  assign popcount33_oce2_core_141 = ~(input_a[13] | input_a[26]);
  assign popcount33_oce2_core_142 = ~(input_a[29] & input_a[26]);
  assign popcount33_oce2_core_143 = ~(input_a[0] & input_a[5]);
  assign popcount33_oce2_core_144 = input_a[29] & input_a[12];
  assign popcount33_oce2_core_145 = ~input_a[4];
  assign popcount33_oce2_core_146 = ~(input_a[21] ^ input_a[1]);
  assign popcount33_oce2_core_148 = input_a[12] & input_a[25];
  assign popcount33_oce2_core_149 = input_a[12] ^ input_a[19];
  assign popcount33_oce2_core_150 = ~input_a[3];
  assign popcount33_oce2_core_151 = ~input_a[7];
  assign popcount33_oce2_core_152 = ~(input_a[28] | input_a[3]);
  assign popcount33_oce2_core_154 = ~(input_a[31] & input_a[27]);
  assign popcount33_oce2_core_156 = ~(input_a[11] | input_a[0]);
  assign popcount33_oce2_core_158 = input_a[27] | input_a[1];
  assign popcount33_oce2_core_159 = input_a[2] | input_a[29];
  assign popcount33_oce2_core_163 = ~(input_a[30] ^ input_a[10]);
  assign popcount33_oce2_core_164 = ~(input_a[13] ^ input_a[30]);
  assign popcount33_oce2_core_165 = ~(input_a[5] ^ input_a[31]);
  assign popcount33_oce2_core_167 = ~input_a[12];
  assign popcount33_oce2_core_171 = input_a[16] & input_a[25];
  assign popcount33_oce2_core_172 = input_a[22] & input_a[6];
  assign popcount33_oce2_core_173 = ~(input_a[12] & input_a[8]);
  assign popcount33_oce2_core_174 = input_a[4] ^ input_a[30];
  assign popcount33_oce2_core_176 = input_a[8] | input_a[1];
  assign popcount33_oce2_core_177 = ~(input_a[6] | input_a[27]);
  assign popcount33_oce2_core_178 = ~(input_a[17] | input_a[28]);
  assign popcount33_oce2_core_180 = ~input_a[30];
  assign popcount33_oce2_core_181 = input_a[24] | input_a[13];
  assign popcount33_oce2_core_182 = input_a[29] & input_a[6];
  assign popcount33_oce2_core_183 = ~(input_a[16] | input_a[13]);
  assign popcount33_oce2_core_185 = ~(input_a[2] & input_a[6]);
  assign popcount33_oce2_core_186_not = ~input_a[16];
  assign popcount33_oce2_core_187 = ~(input_a[18] | input_a[3]);
  assign popcount33_oce2_core_189 = input_a[30] | input_a[20];
  assign popcount33_oce2_core_190 = ~input_a[32];
  assign popcount33_oce2_core_191 = input_a[22] | input_a[24];
  assign popcount33_oce2_core_192 = input_a[31] ^ input_a[32];
  assign popcount33_oce2_core_193 = ~(input_a[25] ^ input_a[6]);
  assign popcount33_oce2_core_194 = input_a[28] | input_a[17];
  assign popcount33_oce2_core_196 = ~(input_a[1] | input_a[27]);
  assign popcount33_oce2_core_197 = input_a[2] | input_a[13];
  assign popcount33_oce2_core_198 = ~input_a[30];
  assign popcount33_oce2_core_199 = ~(input_a[27] ^ input_a[1]);
  assign popcount33_oce2_core_202 = input_a[22] | input_a[28];
  assign popcount33_oce2_core_203 = input_a[2] ^ input_a[32];
  assign popcount33_oce2_core_205 = ~(input_a[10] ^ input_a[27]);
  assign popcount33_oce2_core_206 = ~(input_a[0] | input_a[15]);
  assign popcount33_oce2_core_210 = ~input_a[3];
  assign popcount33_oce2_core_211 = ~(input_a[31] ^ input_a[1]);
  assign popcount33_oce2_core_213 = ~input_a[28];
  assign popcount33_oce2_core_214_not = ~input_a[11];
  assign popcount33_oce2_core_215 = ~(input_a[3] | input_a[18]);
  assign popcount33_oce2_core_216 = ~(input_a[15] | input_a[11]);
  assign popcount33_oce2_core_217 = ~input_a[31];
  assign popcount33_oce2_core_218 = ~input_a[1];
  assign popcount33_oce2_core_220 = ~(input_a[19] ^ input_a[8]);
  assign popcount33_oce2_core_223_not = ~input_a[6];
  assign popcount33_oce2_core_224 = ~(input_a[27] & input_a[18]);
  assign popcount33_oce2_core_225 = ~(input_a[19] & input_a[21]);
  assign popcount33_oce2_core_227 = ~(input_a[29] & input_a[19]);
  assign popcount33_oce2_core_228 = ~(input_a[9] ^ input_a[5]);
  assign popcount33_oce2_core_229 = ~input_a[28];
  assign popcount33_oce2_core_230 = input_a[20] | input_a[7];
  assign popcount33_oce2_core_231 = ~(input_a[7] & input_a[32]);
  assign popcount33_oce2_core_234 = ~(input_a[16] & input_a[9]);
  assign popcount33_oce2_core_235 = input_a[3] | input_a[2];
  assign popcount33_oce2_core_236 = ~(input_a[22] ^ input_a[5]);
  assign popcount33_oce2_core_237 = ~input_a[25];

  assign popcount33_oce2_out[0] = input_a[29];
  assign popcount33_oce2_out[1] = 1'b1;
  assign popcount33_oce2_out[2] = popcount33_oce2_core_229;
  assign popcount33_oce2_out[3] = popcount33_oce2_core_229;
  assign popcount33_oce2_out[4] = input_a[28];
  assign popcount33_oce2_out[5] = 1'b0;
endmodule