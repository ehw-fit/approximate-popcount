// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.56885
// WCE=6.0
// EP=0.810303%
// Printed PDK parameters:
//  Area=55256082.0
//  Delay=68428168.0
//  Power=3102600.0

module popcount28_fqia(input [27:0] input_a, output [4:0] popcount28_fqia_out);
  wire popcount28_fqia_core_030;
  wire popcount28_fqia_core_031;
  wire popcount28_fqia_core_033;
  wire popcount28_fqia_core_034;
  wire popcount28_fqia_core_036;
  wire popcount28_fqia_core_037;
  wire popcount28_fqia_core_038;
  wire popcount28_fqia_core_039;
  wire popcount28_fqia_core_040;
  wire popcount28_fqia_core_041;
  wire popcount28_fqia_core_042;
  wire popcount28_fqia_core_043;
  wire popcount28_fqia_core_044;
  wire popcount28_fqia_core_045;
  wire popcount28_fqia_core_047;
  wire popcount28_fqia_core_048;
  wire popcount28_fqia_core_049;
  wire popcount28_fqia_core_050;
  wire popcount28_fqia_core_051;
  wire popcount28_fqia_core_052;
  wire popcount28_fqia_core_053;
  wire popcount28_fqia_core_055;
  wire popcount28_fqia_core_056;
  wire popcount28_fqia_core_057;
  wire popcount28_fqia_core_058;
  wire popcount28_fqia_core_059;
  wire popcount28_fqia_core_060;
  wire popcount28_fqia_core_061;
  wire popcount28_fqia_core_063;
  wire popcount28_fqia_core_064;
  wire popcount28_fqia_core_066;
  wire popcount28_fqia_core_067;
  wire popcount28_fqia_core_068;
  wire popcount28_fqia_core_070;
  wire popcount28_fqia_core_071;
  wire popcount28_fqia_core_072;
  wire popcount28_fqia_core_073_not;
  wire popcount28_fqia_core_074;
  wire popcount28_fqia_core_075_not;
  wire popcount28_fqia_core_076;
  wire popcount28_fqia_core_077;
  wire popcount28_fqia_core_079;
  wire popcount28_fqia_core_080;
  wire popcount28_fqia_core_081;
  wire popcount28_fqia_core_082;
  wire popcount28_fqia_core_085;
  wire popcount28_fqia_core_086;
  wire popcount28_fqia_core_089;
  wire popcount28_fqia_core_090;
  wire popcount28_fqia_core_091;
  wire popcount28_fqia_core_092;
  wire popcount28_fqia_core_093;
  wire popcount28_fqia_core_094;
  wire popcount28_fqia_core_097;
  wire popcount28_fqia_core_098;
  wire popcount28_fqia_core_101_not;
  wire popcount28_fqia_core_105;
  wire popcount28_fqia_core_106;
  wire popcount28_fqia_core_107;
  wire popcount28_fqia_core_111;
  wire popcount28_fqia_core_112;
  wire popcount28_fqia_core_113;
  wire popcount28_fqia_core_114;
  wire popcount28_fqia_core_115;
  wire popcount28_fqia_core_116;
  wire popcount28_fqia_core_117;
  wire popcount28_fqia_core_118;
  wire popcount28_fqia_core_119;
  wire popcount28_fqia_core_122;
  wire popcount28_fqia_core_123;
  wire popcount28_fqia_core_124;
  wire popcount28_fqia_core_125;
  wire popcount28_fqia_core_126;
  wire popcount28_fqia_core_127;
  wire popcount28_fqia_core_128;
  wire popcount28_fqia_core_130;
  wire popcount28_fqia_core_131;
  wire popcount28_fqia_core_134;
  wire popcount28_fqia_core_135;
  wire popcount28_fqia_core_136;
  wire popcount28_fqia_core_137;
  wire popcount28_fqia_core_138;
  wire popcount28_fqia_core_139;
  wire popcount28_fqia_core_143;
  wire popcount28_fqia_core_144;
  wire popcount28_fqia_core_145;
  wire popcount28_fqia_core_148;
  wire popcount28_fqia_core_149;
  wire popcount28_fqia_core_151;
  wire popcount28_fqia_core_153;
  wire popcount28_fqia_core_154;
  wire popcount28_fqia_core_158;
  wire popcount28_fqia_core_160;
  wire popcount28_fqia_core_161;
  wire popcount28_fqia_core_163;
  wire popcount28_fqia_core_164;
  wire popcount28_fqia_core_165;
  wire popcount28_fqia_core_166;
  wire popcount28_fqia_core_167;
  wire popcount28_fqia_core_168;
  wire popcount28_fqia_core_169;
  wire popcount28_fqia_core_170;
  wire popcount28_fqia_core_171;
  wire popcount28_fqia_core_172;
  wire popcount28_fqia_core_173;
  wire popcount28_fqia_core_174;
  wire popcount28_fqia_core_177;
  wire popcount28_fqia_core_178;
  wire popcount28_fqia_core_180;
  wire popcount28_fqia_core_181;
  wire popcount28_fqia_core_182;
  wire popcount28_fqia_core_183;
  wire popcount28_fqia_core_184;
  wire popcount28_fqia_core_185;
  wire popcount28_fqia_core_186;
  wire popcount28_fqia_core_187;
  wire popcount28_fqia_core_188;
  wire popcount28_fqia_core_189;
  wire popcount28_fqia_core_190;
  wire popcount28_fqia_core_191;
  wire popcount28_fqia_core_192;
  wire popcount28_fqia_core_193;
  wire popcount28_fqia_core_194;
  wire popcount28_fqia_core_195;
  wire popcount28_fqia_core_196;
  wire popcount28_fqia_core_198;
  wire popcount28_fqia_core_199;
  wire popcount28_fqia_core_201;

  assign popcount28_fqia_core_030 = input_a[1] | input_a[2];
  assign popcount28_fqia_core_031 = input_a[1] & input_a[2];
  assign popcount28_fqia_core_033 = input_a[7] & popcount28_fqia_core_030;
  assign popcount28_fqia_core_034 = popcount28_fqia_core_031 | popcount28_fqia_core_033;
  assign popcount28_fqia_core_036 = input_a[3] ^ input_a[4];
  assign popcount28_fqia_core_037 = input_a[3] & input_a[4];
  assign popcount28_fqia_core_038 = input_a[5] ^ input_a[6];
  assign popcount28_fqia_core_039 = input_a[5] & input_a[6];
  assign popcount28_fqia_core_040 = popcount28_fqia_core_036 ^ popcount28_fqia_core_038;
  assign popcount28_fqia_core_041 = popcount28_fqia_core_036 & popcount28_fqia_core_038;
  assign popcount28_fqia_core_042 = popcount28_fqia_core_037 ^ popcount28_fqia_core_039;
  assign popcount28_fqia_core_043 = popcount28_fqia_core_037 & popcount28_fqia_core_039;
  assign popcount28_fqia_core_044 = popcount28_fqia_core_042 | popcount28_fqia_core_041;
  assign popcount28_fqia_core_045 = ~(input_a[12] & input_a[15]);
  assign popcount28_fqia_core_047 = input_a[14] ^ input_a[15];
  assign popcount28_fqia_core_048 = input_a[9] & popcount28_fqia_core_040;
  assign popcount28_fqia_core_049 = popcount28_fqia_core_034 ^ popcount28_fqia_core_044;
  assign popcount28_fqia_core_050 = popcount28_fqia_core_034 & popcount28_fqia_core_044;
  assign popcount28_fqia_core_051 = popcount28_fqia_core_049 ^ popcount28_fqia_core_048;
  assign popcount28_fqia_core_052 = popcount28_fqia_core_049 & popcount28_fqia_core_048;
  assign popcount28_fqia_core_053 = popcount28_fqia_core_050 | popcount28_fqia_core_052;
  assign popcount28_fqia_core_055 = ~(input_a[11] | input_a[17]);
  assign popcount28_fqia_core_056 = popcount28_fqia_core_043 | popcount28_fqia_core_053;
  assign popcount28_fqia_core_057 = ~input_a[21];
  assign popcount28_fqia_core_058 = ~(input_a[11] | input_a[25]);
  assign popcount28_fqia_core_059 = input_a[13] ^ input_a[20];
  assign popcount28_fqia_core_060 = ~input_a[16];
  assign popcount28_fqia_core_061 = ~input_a[18];
  assign popcount28_fqia_core_063 = input_a[3] & input_a[8];
  assign popcount28_fqia_core_064 = input_a[18] | input_a[1];
  assign popcount28_fqia_core_066 = input_a[17] ^ input_a[2];
  assign popcount28_fqia_core_067 = input_a[20] & input_a[27];
  assign popcount28_fqia_core_068 = input_a[12] & input_a[18];
  assign popcount28_fqia_core_070 = ~(input_a[5] ^ input_a[25]);
  assign popcount28_fqia_core_071 = input_a[22] & input_a[15];
  assign popcount28_fqia_core_072 = input_a[3] | input_a[6];
  assign popcount28_fqia_core_073_not = ~input_a[22];
  assign popcount28_fqia_core_074 = ~(input_a[3] ^ input_a[12]);
  assign popcount28_fqia_core_075_not = ~input_a[21];
  assign popcount28_fqia_core_076 = ~(input_a[20] ^ input_a[13]);
  assign popcount28_fqia_core_077 = ~(input_a[14] | input_a[6]);
  assign popcount28_fqia_core_079 = input_a[25] & input_a[11];
  assign popcount28_fqia_core_080 = input_a[0] | input_a[27];
  assign popcount28_fqia_core_081 = input_a[9] | input_a[8];
  assign popcount28_fqia_core_082 = input_a[15] | input_a[16];
  assign popcount28_fqia_core_085 = input_a[5] ^ input_a[25];
  assign popcount28_fqia_core_086 = input_a[26] | input_a[5];
  assign popcount28_fqia_core_089 = ~input_a[16];
  assign popcount28_fqia_core_090 = popcount28_fqia_core_051 ^ popcount28_fqia_core_080;
  assign popcount28_fqia_core_091 = popcount28_fqia_core_051 & popcount28_fqia_core_080;
  assign popcount28_fqia_core_092 = popcount28_fqia_core_090 ^ input_a[25];
  assign popcount28_fqia_core_093 = popcount28_fqia_core_090 & input_a[25];
  assign popcount28_fqia_core_094 = popcount28_fqia_core_091 | popcount28_fqia_core_093;
  assign popcount28_fqia_core_097 = popcount28_fqia_core_056 ^ popcount28_fqia_core_094;
  assign popcount28_fqia_core_098 = popcount28_fqia_core_056 & popcount28_fqia_core_094;
  assign popcount28_fqia_core_101_not = ~input_a[3];
  assign popcount28_fqia_core_105 = input_a[13] ^ input_a[25];
  assign popcount28_fqia_core_106 = input_a[23] & input_a[8];
  assign popcount28_fqia_core_107 = ~(input_a[15] | input_a[16]);
  assign popcount28_fqia_core_111 = input_a[17] ^ input_a[18];
  assign popcount28_fqia_core_112 = input_a[17] & input_a[18];
  assign popcount28_fqia_core_113 = input_a[19] ^ input_a[20];
  assign popcount28_fqia_core_114 = input_a[19] & input_a[20];
  assign popcount28_fqia_core_115 = popcount28_fqia_core_111 ^ popcount28_fqia_core_113;
  assign popcount28_fqia_core_116 = popcount28_fqia_core_111 & popcount28_fqia_core_113;
  assign popcount28_fqia_core_117 = popcount28_fqia_core_112 ^ popcount28_fqia_core_114;
  assign popcount28_fqia_core_118 = popcount28_fqia_core_112 & popcount28_fqia_core_114;
  assign popcount28_fqia_core_119 = popcount28_fqia_core_117 | popcount28_fqia_core_116;
  assign popcount28_fqia_core_122 = input_a[14] ^ popcount28_fqia_core_115;
  assign popcount28_fqia_core_123 = input_a[14] & popcount28_fqia_core_115;
  assign popcount28_fqia_core_124 = popcount28_fqia_core_106 ^ popcount28_fqia_core_119;
  assign popcount28_fqia_core_125 = popcount28_fqia_core_106 & popcount28_fqia_core_119;
  assign popcount28_fqia_core_126 = popcount28_fqia_core_124 ^ popcount28_fqia_core_123;
  assign popcount28_fqia_core_127 = popcount28_fqia_core_124 & popcount28_fqia_core_123;
  assign popcount28_fqia_core_128 = popcount28_fqia_core_125 | popcount28_fqia_core_127;
  assign popcount28_fqia_core_130 = input_a[0] & input_a[20];
  assign popcount28_fqia_core_131 = popcount28_fqia_core_118 | popcount28_fqia_core_128;
  assign popcount28_fqia_core_134 = ~(input_a[26] | input_a[5]);
  assign popcount28_fqia_core_135 = input_a[22] & input_a[21];
  assign popcount28_fqia_core_136 = input_a[24] | input_a[12];
  assign popcount28_fqia_core_137 = input_a[15] & input_a[12];
  assign popcount28_fqia_core_138 = popcount28_fqia_core_135 | popcount28_fqia_core_137;
  assign popcount28_fqia_core_139 = input_a[12] | input_a[25];
  assign popcount28_fqia_core_143 = ~(input_a[10] ^ input_a[20]);
  assign popcount28_fqia_core_144 = ~(input_a[17] ^ input_a[8]);
  assign popcount28_fqia_core_145 = ~(input_a[18] | input_a[3]);
  assign popcount28_fqia_core_148 = input_a[21] & input_a[24];
  assign popcount28_fqia_core_149 = input_a[25] & input_a[18];
  assign popcount28_fqia_core_151 = input_a[25] ^ input_a[14];
  assign popcount28_fqia_core_153 = popcount28_fqia_core_138 ^ input_a[16];
  assign popcount28_fqia_core_154 = popcount28_fqia_core_138 & input_a[16];
  assign popcount28_fqia_core_158 = input_a[11] | input_a[10];
  assign popcount28_fqia_core_160 = popcount28_fqia_core_158 ^ popcount28_fqia_core_154;
  assign popcount28_fqia_core_161 = popcount28_fqia_core_158 & popcount28_fqia_core_154;
  assign popcount28_fqia_core_163 = popcount28_fqia_core_122 ^ input_a[26];
  assign popcount28_fqia_core_164 = popcount28_fqia_core_122 & input_a[26];
  assign popcount28_fqia_core_165 = popcount28_fqia_core_126 ^ popcount28_fqia_core_153;
  assign popcount28_fqia_core_166 = popcount28_fqia_core_126 & popcount28_fqia_core_153;
  assign popcount28_fqia_core_167 = popcount28_fqia_core_165 ^ popcount28_fqia_core_164;
  assign popcount28_fqia_core_168 = popcount28_fqia_core_165 & popcount28_fqia_core_164;
  assign popcount28_fqia_core_169 = popcount28_fqia_core_166 | popcount28_fqia_core_168;
  assign popcount28_fqia_core_170 = popcount28_fqia_core_131 ^ popcount28_fqia_core_160;
  assign popcount28_fqia_core_171 = popcount28_fqia_core_131 & popcount28_fqia_core_160;
  assign popcount28_fqia_core_172 = popcount28_fqia_core_170 ^ popcount28_fqia_core_169;
  assign popcount28_fqia_core_173 = popcount28_fqia_core_170 & popcount28_fqia_core_169;
  assign popcount28_fqia_core_174 = popcount28_fqia_core_171 | popcount28_fqia_core_173;
  assign popcount28_fqia_core_177 = popcount28_fqia_core_161 ^ popcount28_fqia_core_174;
  assign popcount28_fqia_core_178 = popcount28_fqia_core_161 & popcount28_fqia_core_174;
  assign popcount28_fqia_core_180 = input_a[23] ^ input_a[12];
  assign popcount28_fqia_core_181 = input_a[24] & popcount28_fqia_core_163;
  assign popcount28_fqia_core_182 = popcount28_fqia_core_092 ^ popcount28_fqia_core_167;
  assign popcount28_fqia_core_183 = popcount28_fqia_core_092 & popcount28_fqia_core_167;
  assign popcount28_fqia_core_184 = popcount28_fqia_core_182 ^ popcount28_fqia_core_181;
  assign popcount28_fqia_core_185 = popcount28_fqia_core_182 & popcount28_fqia_core_181;
  assign popcount28_fqia_core_186 = popcount28_fqia_core_183 | popcount28_fqia_core_185;
  assign popcount28_fqia_core_187 = popcount28_fqia_core_097 ^ popcount28_fqia_core_172;
  assign popcount28_fqia_core_188 = popcount28_fqia_core_097 & popcount28_fqia_core_172;
  assign popcount28_fqia_core_189 = popcount28_fqia_core_187 ^ popcount28_fqia_core_186;
  assign popcount28_fqia_core_190 = popcount28_fqia_core_187 & popcount28_fqia_core_186;
  assign popcount28_fqia_core_191 = popcount28_fqia_core_188 | popcount28_fqia_core_190;
  assign popcount28_fqia_core_192 = popcount28_fqia_core_098 ^ popcount28_fqia_core_177;
  assign popcount28_fqia_core_193 = popcount28_fqia_core_098 & popcount28_fqia_core_177;
  assign popcount28_fqia_core_194 = popcount28_fqia_core_192 ^ popcount28_fqia_core_191;
  assign popcount28_fqia_core_195 = popcount28_fqia_core_192 & popcount28_fqia_core_191;
  assign popcount28_fqia_core_196 = popcount28_fqia_core_193 | popcount28_fqia_core_195;
  assign popcount28_fqia_core_198 = input_a[20] | input_a[3];
  assign popcount28_fqia_core_199 = popcount28_fqia_core_178 | popcount28_fqia_core_196;
  assign popcount28_fqia_core_201 = input_a[25] | input_a[4];

  assign popcount28_fqia_out[0] = input_a[13];
  assign popcount28_fqia_out[1] = popcount28_fqia_core_184;
  assign popcount28_fqia_out[2] = popcount28_fqia_core_189;
  assign popcount28_fqia_out[3] = popcount28_fqia_core_194;
  assign popcount28_fqia_out[4] = popcount28_fqia_core_199;
endmodule