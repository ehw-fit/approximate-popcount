// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.23047
// WCE=5.0
// EP=0.753906%
// Printed PDK parameters:
//  Area=37279120.0
//  Delay=58922736.0
//  Power=1615800.0

module popcount25_3f06(input [24:0] input_a, output [4:0] popcount25_3f06_out);
  wire popcount25_3f06_core_027;
  wire popcount25_3f06_core_028;
  wire popcount25_3f06_core_029;
  wire popcount25_3f06_core_032;
  wire popcount25_3f06_core_033;
  wire popcount25_3f06_core_034;
  wire popcount25_3f06_core_035;
  wire popcount25_3f06_core_037;
  wire popcount25_3f06_core_038;
  wire popcount25_3f06_core_039;
  wire popcount25_3f06_core_040;
  wire popcount25_3f06_core_041;
  wire popcount25_3f06_core_042;
  wire popcount25_3f06_core_043;
  wire popcount25_3f06_core_044;
  wire popcount25_3f06_core_045;
  wire popcount25_3f06_core_049;
  wire popcount25_3f06_core_051;
  wire popcount25_3f06_core_052;
  wire popcount25_3f06_core_054;
  wire popcount25_3f06_core_055;
  wire popcount25_3f06_core_057;
  wire popcount25_3f06_core_058;
  wire popcount25_3f06_core_059;
  wire popcount25_3f06_core_060;
  wire popcount25_3f06_core_061;
  wire popcount25_3f06_core_062;
  wire popcount25_3f06_core_063;
  wire popcount25_3f06_core_065;
  wire popcount25_3f06_core_066;
  wire popcount25_3f06_core_076;
  wire popcount25_3f06_core_077;
  wire popcount25_3f06_core_078;
  wire popcount25_3f06_core_079;
  wire popcount25_3f06_core_080;
  wire popcount25_3f06_core_081;
  wire popcount25_3f06_core_082;
  wire popcount25_3f06_core_083;
  wire popcount25_3f06_core_084;
  wire popcount25_3f06_core_085;
  wire popcount25_3f06_core_086;
  wire popcount25_3f06_core_090;
  wire popcount25_3f06_core_092;
  wire popcount25_3f06_core_094;
  wire popcount25_3f06_core_095;
  wire popcount25_3f06_core_097;
  wire popcount25_3f06_core_098;
  wire popcount25_3f06_core_099;
  wire popcount25_3f06_core_100;
  wire popcount25_3f06_core_101;
  wire popcount25_3f06_core_102;
  wire popcount25_3f06_core_103;
  wire popcount25_3f06_core_104;
  wire popcount25_3f06_core_105;
  wire popcount25_3f06_core_106;
  wire popcount25_3f06_core_107;
  wire popcount25_3f06_core_112;
  wire popcount25_3f06_core_114;
  wire popcount25_3f06_core_115;
  wire popcount25_3f06_core_121;
  wire popcount25_3f06_core_122_not;
  wire popcount25_3f06_core_123;
  wire popcount25_3f06_core_125;
  wire popcount25_3f06_core_126;
  wire popcount25_3f06_core_127;
  wire popcount25_3f06_core_128;
  wire popcount25_3f06_core_131;
  wire popcount25_3f06_core_132;
  wire popcount25_3f06_core_133;
  wire popcount25_3f06_core_134;
  wire popcount25_3f06_core_135_not;
  wire popcount25_3f06_core_141;
  wire popcount25_3f06_core_145;
  wire popcount25_3f06_core_146;
  wire popcount25_3f06_core_147;
  wire popcount25_3f06_core_148;
  wire popcount25_3f06_core_149;
  wire popcount25_3f06_core_150;
  wire popcount25_3f06_core_151;
  wire popcount25_3f06_core_152;
  wire popcount25_3f06_core_153;
  wire popcount25_3f06_core_154;
  wire popcount25_3f06_core_155;
  wire popcount25_3f06_core_156;
  wire popcount25_3f06_core_158;
  wire popcount25_3f06_core_161;
  wire popcount25_3f06_core_164;
  wire popcount25_3f06_core_166;
  wire popcount25_3f06_core_168;
  wire popcount25_3f06_core_169;
  wire popcount25_3f06_core_170;
  wire popcount25_3f06_core_171;
  wire popcount25_3f06_core_172;
  wire popcount25_3f06_core_173;
  wire popcount25_3f06_core_174;
  wire popcount25_3f06_core_175;
  wire popcount25_3f06_core_176;
  wire popcount25_3f06_core_177;
  wire popcount25_3f06_core_178;
  wire popcount25_3f06_core_180;
  wire popcount25_3f06_core_181_not;

  assign popcount25_3f06_core_027 = ~(input_a[3] | input_a[22]);
  assign popcount25_3f06_core_028 = input_a[1] & input_a[2];
  assign popcount25_3f06_core_029 = ~(input_a[23] & input_a[12]);
  assign popcount25_3f06_core_032 = ~(input_a[16] & input_a[15]);
  assign popcount25_3f06_core_033 = ~input_a[5];
  assign popcount25_3f06_core_034 = input_a[4] & input_a[5];
  assign popcount25_3f06_core_035 = ~(input_a[3] & popcount25_3f06_core_033);
  assign popcount25_3f06_core_037 = popcount25_3f06_core_034 | input_a[3];
  assign popcount25_3f06_core_038 = ~(input_a[16] ^ input_a[1]);
  assign popcount25_3f06_core_039 = input_a[0] ^ popcount25_3f06_core_035;
  assign popcount25_3f06_core_040 = input_a[0] & popcount25_3f06_core_035;
  assign popcount25_3f06_core_041 = popcount25_3f06_core_028 ^ popcount25_3f06_core_037;
  assign popcount25_3f06_core_042 = popcount25_3f06_core_028 & popcount25_3f06_core_037;
  assign popcount25_3f06_core_043 = popcount25_3f06_core_041 ^ popcount25_3f06_core_040;
  assign popcount25_3f06_core_044 = popcount25_3f06_core_041 & popcount25_3f06_core_040;
  assign popcount25_3f06_core_045 = popcount25_3f06_core_042 | popcount25_3f06_core_044;
  assign popcount25_3f06_core_049 = ~(input_a[7] & input_a[6]);
  assign popcount25_3f06_core_051 = input_a[7] | input_a[8];
  assign popcount25_3f06_core_052 = input_a[7] & input_a[8];
  assign popcount25_3f06_core_054 = input_a[6] & popcount25_3f06_core_051;
  assign popcount25_3f06_core_055 = popcount25_3f06_core_052 | popcount25_3f06_core_054;
  assign popcount25_3f06_core_057 = input_a[10] | input_a[11];
  assign popcount25_3f06_core_058 = input_a[10] & input_a[11];
  assign popcount25_3f06_core_059 = input_a[11] | input_a[19];
  assign popcount25_3f06_core_060 = input_a[9] & popcount25_3f06_core_057;
  assign popcount25_3f06_core_061 = popcount25_3f06_core_058 | popcount25_3f06_core_060;
  assign popcount25_3f06_core_062 = ~(input_a[1] | input_a[1]);
  assign popcount25_3f06_core_063 = input_a[6] & input_a[15];
  assign popcount25_3f06_core_065 = popcount25_3f06_core_055 ^ popcount25_3f06_core_061;
  assign popcount25_3f06_core_066 = popcount25_3f06_core_055 & popcount25_3f06_core_061;
  assign popcount25_3f06_core_076 = popcount25_3f06_core_039 & input_a[20];
  assign popcount25_3f06_core_077 = popcount25_3f06_core_043 ^ popcount25_3f06_core_065;
  assign popcount25_3f06_core_078 = popcount25_3f06_core_043 & popcount25_3f06_core_065;
  assign popcount25_3f06_core_079 = popcount25_3f06_core_077 ^ popcount25_3f06_core_076;
  assign popcount25_3f06_core_080 = popcount25_3f06_core_077 & popcount25_3f06_core_076;
  assign popcount25_3f06_core_081 = popcount25_3f06_core_078 | popcount25_3f06_core_080;
  assign popcount25_3f06_core_082 = popcount25_3f06_core_045 ^ popcount25_3f06_core_066;
  assign popcount25_3f06_core_083 = popcount25_3f06_core_045 & popcount25_3f06_core_066;
  assign popcount25_3f06_core_084 = popcount25_3f06_core_082 ^ popcount25_3f06_core_081;
  assign popcount25_3f06_core_085 = popcount25_3f06_core_082 & popcount25_3f06_core_081;
  assign popcount25_3f06_core_086 = popcount25_3f06_core_083 | popcount25_3f06_core_085;
  assign popcount25_3f06_core_090 = input_a[8] | input_a[7];
  assign popcount25_3f06_core_092 = ~input_a[11];
  assign popcount25_3f06_core_094 = ~(input_a[22] | input_a[21]);
  assign popcount25_3f06_core_095 = input_a[12] & input_a[14];
  assign popcount25_3f06_core_097 = input_a[5] & input_a[13];
  assign popcount25_3f06_core_098 = input_a[16] | input_a[17];
  assign popcount25_3f06_core_099 = input_a[16] & input_a[17];
  assign popcount25_3f06_core_100 = input_a[15] ^ input_a[6];
  assign popcount25_3f06_core_101 = input_a[15] & popcount25_3f06_core_098;
  assign popcount25_3f06_core_102 = popcount25_3f06_core_099 | popcount25_3f06_core_101;
  assign popcount25_3f06_core_103 = ~(input_a[16] ^ input_a[5]);
  assign popcount25_3f06_core_104 = input_a[1] | input_a[24];
  assign popcount25_3f06_core_105 = input_a[4] & input_a[9];
  assign popcount25_3f06_core_106 = popcount25_3f06_core_095 ^ popcount25_3f06_core_102;
  assign popcount25_3f06_core_107 = popcount25_3f06_core_095 & popcount25_3f06_core_102;
  assign popcount25_3f06_core_112 = ~(input_a[11] ^ input_a[11]);
  assign popcount25_3f06_core_114 = ~input_a[7];
  assign popcount25_3f06_core_115 = input_a[14] ^ input_a[17];
  assign popcount25_3f06_core_121 = input_a[24] ^ input_a[1];
  assign popcount25_3f06_core_122_not = ~input_a[16];
  assign popcount25_3f06_core_123 = input_a[21] & input_a[22];
  assign popcount25_3f06_core_125 = input_a[23] & input_a[24];
  assign popcount25_3f06_core_126 = input_a[8] | input_a[8];
  assign popcount25_3f06_core_127 = input_a[17] ^ input_a[15];
  assign popcount25_3f06_core_128 = popcount25_3f06_core_123 | popcount25_3f06_core_125;
  assign popcount25_3f06_core_131 = input_a[7] | input_a[22];
  assign popcount25_3f06_core_132 = ~(input_a[6] ^ input_a[4]);
  assign popcount25_3f06_core_133 = input_a[18] | input_a[7];
  assign popcount25_3f06_core_134 = input_a[10] | input_a[0];
  assign popcount25_3f06_core_135_not = ~popcount25_3f06_core_128;
  assign popcount25_3f06_core_141 = ~(input_a[22] & input_a[2]);
  assign popcount25_3f06_core_145 = ~input_a[4];
  assign popcount25_3f06_core_146 = input_a[19] & input_a[18];
  assign popcount25_3f06_core_147 = popcount25_3f06_core_106 ^ popcount25_3f06_core_135_not;
  assign popcount25_3f06_core_148 = popcount25_3f06_core_106 & popcount25_3f06_core_135_not;
  assign popcount25_3f06_core_149 = popcount25_3f06_core_147 ^ popcount25_3f06_core_146;
  assign popcount25_3f06_core_150 = popcount25_3f06_core_147 & popcount25_3f06_core_146;
  assign popcount25_3f06_core_151 = popcount25_3f06_core_148 | popcount25_3f06_core_150;
  assign popcount25_3f06_core_152 = popcount25_3f06_core_107 ^ popcount25_3f06_core_128;
  assign popcount25_3f06_core_153 = popcount25_3f06_core_107 & popcount25_3f06_core_128;
  assign popcount25_3f06_core_154 = popcount25_3f06_core_152 ^ popcount25_3f06_core_151;
  assign popcount25_3f06_core_155 = popcount25_3f06_core_152 & popcount25_3f06_core_151;
  assign popcount25_3f06_core_156 = popcount25_3f06_core_153 | popcount25_3f06_core_155;
  assign popcount25_3f06_core_158 = ~(input_a[20] ^ input_a[23]);
  assign popcount25_3f06_core_161 = ~(input_a[5] & input_a[20]);
  assign popcount25_3f06_core_164 = popcount25_3f06_core_079 ^ popcount25_3f06_core_149;
  assign popcount25_3f06_core_166 = ~popcount25_3f06_core_164;
  assign popcount25_3f06_core_168 = popcount25_3f06_core_079 | popcount25_3f06_core_164;
  assign popcount25_3f06_core_169 = popcount25_3f06_core_084 ^ popcount25_3f06_core_154;
  assign popcount25_3f06_core_170 = popcount25_3f06_core_084 & popcount25_3f06_core_154;
  assign popcount25_3f06_core_171 = popcount25_3f06_core_169 ^ popcount25_3f06_core_168;
  assign popcount25_3f06_core_172 = popcount25_3f06_core_169 & popcount25_3f06_core_168;
  assign popcount25_3f06_core_173 = popcount25_3f06_core_170 | popcount25_3f06_core_172;
  assign popcount25_3f06_core_174 = popcount25_3f06_core_086 ^ popcount25_3f06_core_156;
  assign popcount25_3f06_core_175 = popcount25_3f06_core_086 & popcount25_3f06_core_156;
  assign popcount25_3f06_core_176 = popcount25_3f06_core_174 ^ popcount25_3f06_core_173;
  assign popcount25_3f06_core_177 = popcount25_3f06_core_174 & popcount25_3f06_core_173;
  assign popcount25_3f06_core_178 = popcount25_3f06_core_175 | popcount25_3f06_core_177;
  assign popcount25_3f06_core_180 = input_a[24] ^ input_a[6];
  assign popcount25_3f06_core_181_not = ~input_a[1];

  assign popcount25_3f06_out[0] = input_a[13];
  assign popcount25_3f06_out[1] = popcount25_3f06_core_166;
  assign popcount25_3f06_out[2] = popcount25_3f06_core_171;
  assign popcount25_3f06_out[3] = popcount25_3f06_core_176;
  assign popcount25_3f06_out[4] = popcount25_3f06_core_178;
endmodule