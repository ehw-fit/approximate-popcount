// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.15146
// WCE=11.0
// EP=0.857946%
// Printed PDK parameters:
//  Area=2300720.0
//  Delay=10025376.0
//  Power=119680.0

module popcount22_n1n6(input [21:0] input_a, output [4:0] popcount22_n1n6_out);
  wire popcount22_n1n6_core_026;
  wire popcount22_n1n6_core_027;
  wire popcount22_n1n6_core_028;
  wire popcount22_n1n6_core_030;
  wire popcount22_n1n6_core_031;
  wire popcount22_n1n6_core_032;
  wire popcount22_n1n6_core_035;
  wire popcount22_n1n6_core_036;
  wire popcount22_n1n6_core_038;
  wire popcount22_n1n6_core_040;
  wire popcount22_n1n6_core_042;
  wire popcount22_n1n6_core_043;
  wire popcount22_n1n6_core_044;
  wire popcount22_n1n6_core_045;
  wire popcount22_n1n6_core_046;
  wire popcount22_n1n6_core_047;
  wire popcount22_n1n6_core_048;
  wire popcount22_n1n6_core_051;
  wire popcount22_n1n6_core_054;
  wire popcount22_n1n6_core_055;
  wire popcount22_n1n6_core_058;
  wire popcount22_n1n6_core_059;
  wire popcount22_n1n6_core_060;
  wire popcount22_n1n6_core_062;
  wire popcount22_n1n6_core_064;
  wire popcount22_n1n6_core_065;
  wire popcount22_n1n6_core_066;
  wire popcount22_n1n6_core_068;
  wire popcount22_n1n6_core_069;
  wire popcount22_n1n6_core_070;
  wire popcount22_n1n6_core_071;
  wire popcount22_n1n6_core_072;
  wire popcount22_n1n6_core_074;
  wire popcount22_n1n6_core_076_not;
  wire popcount22_n1n6_core_077;
  wire popcount22_n1n6_core_078;
  wire popcount22_n1n6_core_079;
  wire popcount22_n1n6_core_080;
  wire popcount22_n1n6_core_081;
  wire popcount22_n1n6_core_082;
  wire popcount22_n1n6_core_083_not;
  wire popcount22_n1n6_core_084;
  wire popcount22_n1n6_core_085;
  wire popcount22_n1n6_core_086;
  wire popcount22_n1n6_core_087;
  wire popcount22_n1n6_core_088;
  wire popcount22_n1n6_core_089;
  wire popcount22_n1n6_core_090;
  wire popcount22_n1n6_core_092;
  wire popcount22_n1n6_core_094;
  wire popcount22_n1n6_core_095;
  wire popcount22_n1n6_core_098;
  wire popcount22_n1n6_core_099;
  wire popcount22_n1n6_core_101;
  wire popcount22_n1n6_core_102;
  wire popcount22_n1n6_core_104;
  wire popcount22_n1n6_core_105;
  wire popcount22_n1n6_core_107;
  wire popcount22_n1n6_core_108;
  wire popcount22_n1n6_core_109;
  wire popcount22_n1n6_core_110;
  wire popcount22_n1n6_core_111;
  wire popcount22_n1n6_core_112;
  wire popcount22_n1n6_core_116;
  wire popcount22_n1n6_core_117;
  wire popcount22_n1n6_core_119;
  wire popcount22_n1n6_core_120;
  wire popcount22_n1n6_core_121;
  wire popcount22_n1n6_core_124;
  wire popcount22_n1n6_core_127_not;
  wire popcount22_n1n6_core_128_not;
  wire popcount22_n1n6_core_129;
  wire popcount22_n1n6_core_130;
  wire popcount22_n1n6_core_131;
  wire popcount22_n1n6_core_132;
  wire popcount22_n1n6_core_134;
  wire popcount22_n1n6_core_135;
  wire popcount22_n1n6_core_136;
  wire popcount22_n1n6_core_137;
  wire popcount22_n1n6_core_139;
  wire popcount22_n1n6_core_140;
  wire popcount22_n1n6_core_144_not;
  wire popcount22_n1n6_core_147;
  wire popcount22_n1n6_core_149;
  wire popcount22_n1n6_core_153;
  wire popcount22_n1n6_core_154;
  wire popcount22_n1n6_core_155;
  wire popcount22_n1n6_core_157;
  wire popcount22_n1n6_core_158;
  wire popcount22_n1n6_core_161;

  assign popcount22_n1n6_core_026 = ~(input_a[12] | input_a[20]);
  assign popcount22_n1n6_core_027 = input_a[4] ^ input_a[12];
  assign popcount22_n1n6_core_028 = ~input_a[9];
  assign popcount22_n1n6_core_030 = ~(input_a[20] & input_a[14]);
  assign popcount22_n1n6_core_031 = input_a[3] & input_a[10];
  assign popcount22_n1n6_core_032 = input_a[10] & input_a[17];
  assign popcount22_n1n6_core_035 = ~input_a[16];
  assign popcount22_n1n6_core_036 = ~(input_a[12] | input_a[18]);
  assign popcount22_n1n6_core_038 = ~(input_a[16] & input_a[6]);
  assign popcount22_n1n6_core_040 = ~(input_a[10] ^ input_a[11]);
  assign popcount22_n1n6_core_042 = input_a[1] & input_a[5];
  assign popcount22_n1n6_core_043 = ~input_a[11];
  assign popcount22_n1n6_core_044 = ~(input_a[10] & input_a[1]);
  assign popcount22_n1n6_core_045 = ~(input_a[10] | input_a[5]);
  assign popcount22_n1n6_core_046 = ~(input_a[20] ^ input_a[12]);
  assign popcount22_n1n6_core_047 = ~(input_a[0] | input_a[19]);
  assign popcount22_n1n6_core_048 = input_a[8] & input_a[13];
  assign popcount22_n1n6_core_051 = ~(input_a[5] ^ input_a[6]);
  assign popcount22_n1n6_core_054 = ~(input_a[10] & input_a[4]);
  assign popcount22_n1n6_core_055 = ~input_a[19];
  assign popcount22_n1n6_core_058 = input_a[7] ^ input_a[7];
  assign popcount22_n1n6_core_059 = ~(input_a[7] & input_a[12]);
  assign popcount22_n1n6_core_060 = ~input_a[7];
  assign popcount22_n1n6_core_062 = input_a[2] & input_a[1];
  assign popcount22_n1n6_core_064 = ~(input_a[7] | input_a[17]);
  assign popcount22_n1n6_core_065 = input_a[13] ^ input_a[0];
  assign popcount22_n1n6_core_066 = ~input_a[1];
  assign popcount22_n1n6_core_068 = ~(input_a[21] | input_a[8]);
  assign popcount22_n1n6_core_069 = ~(input_a[14] ^ input_a[20]);
  assign popcount22_n1n6_core_070 = input_a[15] ^ input_a[11];
  assign popcount22_n1n6_core_071 = ~input_a[6];
  assign popcount22_n1n6_core_072 = ~(popcount22_n1n6_core_031 & popcount22_n1n6_core_062);
  assign popcount22_n1n6_core_074 = popcount22_n1n6_core_072 ^ input_a[12];
  assign popcount22_n1n6_core_076_not = ~input_a[5];
  assign popcount22_n1n6_core_077 = ~input_a[3];
  assign popcount22_n1n6_core_078 = input_a[19] & input_a[18];
  assign popcount22_n1n6_core_079 = ~input_a[14];
  assign popcount22_n1n6_core_080 = input_a[15] & input_a[8];
  assign popcount22_n1n6_core_081 = ~(input_a[12] & input_a[21]);
  assign popcount22_n1n6_core_082 = ~(input_a[14] | input_a[1]);
  assign popcount22_n1n6_core_083_not = ~input_a[11];
  assign popcount22_n1n6_core_084 = ~(input_a[2] | input_a[21]);
  assign popcount22_n1n6_core_085 = input_a[14] ^ input_a[1];
  assign popcount22_n1n6_core_086 = input_a[20] & input_a[8];
  assign popcount22_n1n6_core_087 = input_a[5] & input_a[14];
  assign popcount22_n1n6_core_088 = ~input_a[12];
  assign popcount22_n1n6_core_089 = input_a[8] ^ input_a[14];
  assign popcount22_n1n6_core_090 = ~input_a[12];
  assign popcount22_n1n6_core_092 = ~(input_a[9] | input_a[14]);
  assign popcount22_n1n6_core_094 = ~(input_a[5] | input_a[2]);
  assign popcount22_n1n6_core_095 = input_a[12] & input_a[15];
  assign popcount22_n1n6_core_098 = ~(input_a[0] | input_a[2]);
  assign popcount22_n1n6_core_099 = ~input_a[12];
  assign popcount22_n1n6_core_101 = input_a[9] & input_a[15];
  assign popcount22_n1n6_core_102 = ~(input_a[3] ^ input_a[12]);
  assign popcount22_n1n6_core_104 = ~(input_a[5] ^ input_a[17]);
  assign popcount22_n1n6_core_105 = ~(input_a[16] & input_a[3]);
  assign popcount22_n1n6_core_107 = input_a[0] ^ input_a[11];
  assign popcount22_n1n6_core_108 = ~input_a[2];
  assign popcount22_n1n6_core_109 = ~(input_a[12] & input_a[6]);
  assign popcount22_n1n6_core_110 = input_a[20] ^ input_a[6];
  assign popcount22_n1n6_core_111 = ~(input_a[1] & input_a[8]);
  assign popcount22_n1n6_core_112 = ~input_a[18];
  assign popcount22_n1n6_core_116 = input_a[20] & input_a[4];
  assign popcount22_n1n6_core_117 = ~(input_a[6] & input_a[14]);
  assign popcount22_n1n6_core_119 = ~(input_a[0] | input_a[14]);
  assign popcount22_n1n6_core_120 = ~(input_a[0] | input_a[7]);
  assign popcount22_n1n6_core_121 = ~input_a[9];
  assign popcount22_n1n6_core_124 = ~(input_a[21] | input_a[7]);
  assign popcount22_n1n6_core_127_not = ~input_a[12];
  assign popcount22_n1n6_core_128_not = ~input_a[21];
  assign popcount22_n1n6_core_129 = input_a[16] | input_a[14];
  assign popcount22_n1n6_core_130 = ~(input_a[6] | input_a[11]);
  assign popcount22_n1n6_core_131 = input_a[12] | input_a[4];
  assign popcount22_n1n6_core_132 = input_a[4] | input_a[15];
  assign popcount22_n1n6_core_134 = input_a[17] ^ input_a[14];
  assign popcount22_n1n6_core_135 = ~input_a[14];
  assign popcount22_n1n6_core_136 = input_a[15] | input_a[9];
  assign popcount22_n1n6_core_137 = input_a[16] ^ input_a[20];
  assign popcount22_n1n6_core_139 = ~(input_a[14] & input_a[17]);
  assign popcount22_n1n6_core_140 = ~(input_a[1] ^ input_a[13]);
  assign popcount22_n1n6_core_144_not = ~input_a[18];
  assign popcount22_n1n6_core_147 = ~popcount22_n1n6_core_074;
  assign popcount22_n1n6_core_149 = input_a[0] ^ input_a[17];
  assign popcount22_n1n6_core_153 = ~input_a[2];
  assign popcount22_n1n6_core_154 = ~(input_a[12] & popcount22_n1n6_core_074);
  assign popcount22_n1n6_core_155 = input_a[12] & popcount22_n1n6_core_074;
  assign popcount22_n1n6_core_157 = ~(input_a[8] ^ input_a[3]);
  assign popcount22_n1n6_core_158 = ~input_a[1];
  assign popcount22_n1n6_core_161 = ~(input_a[14] | input_a[21]);

  assign popcount22_n1n6_out[0] = input_a[9];
  assign popcount22_n1n6_out[1] = 1'b0;
  assign popcount22_n1n6_out[2] = popcount22_n1n6_core_147;
  assign popcount22_n1n6_out[3] = popcount22_n1n6_core_154;
  assign popcount22_n1n6_out[4] = popcount22_n1n6_core_155;
endmodule