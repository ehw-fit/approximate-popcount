// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.61443
// WCE=11.0
// EP=0.887348%
// Printed PDK parameters:
//  Area=17486038.0
//  Delay=38683108.0
//  Power=582210.0

module popcount22_ujfe(input [21:0] input_a, output [4:0] popcount22_ujfe_out);
  wire popcount22_ujfe_core_024;
  wire popcount22_ujfe_core_026;
  wire popcount22_ujfe_core_027;
  wire popcount22_ujfe_core_029;
  wire popcount22_ujfe_core_030;
  wire popcount22_ujfe_core_031;
  wire popcount22_ujfe_core_033;
  wire popcount22_ujfe_core_036;
  wire popcount22_ujfe_core_037;
  wire popcount22_ujfe_core_039;
  wire popcount22_ujfe_core_041;
  wire popcount22_ujfe_core_042;
  wire popcount22_ujfe_core_043;
  wire popcount22_ujfe_core_044;
  wire popcount22_ujfe_core_046_not;
  wire popcount22_ujfe_core_047;
  wire popcount22_ujfe_core_048;
  wire popcount22_ujfe_core_049;
  wire popcount22_ujfe_core_051;
  wire popcount22_ujfe_core_052;
  wire popcount22_ujfe_core_053;
  wire popcount22_ujfe_core_054;
  wire popcount22_ujfe_core_055;
  wire popcount22_ujfe_core_056;
  wire popcount22_ujfe_core_057;
  wire popcount22_ujfe_core_059;
  wire popcount22_ujfe_core_060;
  wire popcount22_ujfe_core_062;
  wire popcount22_ujfe_core_063;
  wire popcount22_ujfe_core_064;
  wire popcount22_ujfe_core_065;
  wire popcount22_ujfe_core_066;
  wire popcount22_ujfe_core_067;
  wire popcount22_ujfe_core_068;
  wire popcount22_ujfe_core_069;
  wire popcount22_ujfe_core_070;
  wire popcount22_ujfe_core_072;
  wire popcount22_ujfe_core_075;
  wire popcount22_ujfe_core_081;
  wire popcount22_ujfe_core_083;
  wire popcount22_ujfe_core_084;
  wire popcount22_ujfe_core_085;
  wire popcount22_ujfe_core_090;
  wire popcount22_ujfe_core_091;
  wire popcount22_ujfe_core_092;
  wire popcount22_ujfe_core_093;
  wire popcount22_ujfe_core_094;
  wire popcount22_ujfe_core_095;
  wire popcount22_ujfe_core_096;
  wire popcount22_ujfe_core_098;
  wire popcount22_ujfe_core_101;
  wire popcount22_ujfe_core_102;
  wire popcount22_ujfe_core_103;
  wire popcount22_ujfe_core_104;
  wire popcount22_ujfe_core_107;
  wire popcount22_ujfe_core_108;
  wire popcount22_ujfe_core_109;
  wire popcount22_ujfe_core_111;
  wire popcount22_ujfe_core_112;
  wire popcount22_ujfe_core_115;
  wire popcount22_ujfe_core_116;
  wire popcount22_ujfe_core_119;
  wire popcount22_ujfe_core_121;
  wire popcount22_ujfe_core_122;
  wire popcount22_ujfe_core_123;
  wire popcount22_ujfe_core_124;
  wire popcount22_ujfe_core_125;
  wire popcount22_ujfe_core_126;
  wire popcount22_ujfe_core_127;
  wire popcount22_ujfe_core_128;
  wire popcount22_ujfe_core_129;
  wire popcount22_ujfe_core_130;
  wire popcount22_ujfe_core_131;
  wire popcount22_ujfe_core_132;
  wire popcount22_ujfe_core_133;
  wire popcount22_ujfe_core_134;
  wire popcount22_ujfe_core_141;
  wire popcount22_ujfe_core_142;
  wire popcount22_ujfe_core_143;
  wire popcount22_ujfe_core_144;
  wire popcount22_ujfe_core_145;
  wire popcount22_ujfe_core_146;
  wire popcount22_ujfe_core_147_not;
  wire popcount22_ujfe_core_150;
  wire popcount22_ujfe_core_152;
  wire popcount22_ujfe_core_153;
  wire popcount22_ujfe_core_154;
  wire popcount22_ujfe_core_155;
  wire popcount22_ujfe_core_156;
  wire popcount22_ujfe_core_158;
  wire popcount22_ujfe_core_159;
  wire popcount22_ujfe_core_161;

  assign popcount22_ujfe_core_024 = ~(input_a[11] ^ input_a[19]);
  assign popcount22_ujfe_core_026 = input_a[15] & input_a[21];
  assign popcount22_ujfe_core_027 = input_a[16] & input_a[0];
  assign popcount22_ujfe_core_029 = input_a[12] & input_a[15];
  assign popcount22_ujfe_core_030 = popcount22_ujfe_core_027 | popcount22_ujfe_core_029;
  assign popcount22_ujfe_core_031 = popcount22_ujfe_core_027 & popcount22_ujfe_core_029;
  assign popcount22_ujfe_core_033 = input_a[13] & input_a[19];
  assign popcount22_ujfe_core_036 = ~(input_a[14] & input_a[5]);
  assign popcount22_ujfe_core_037 = popcount22_ujfe_core_030 & popcount22_ujfe_core_033;
  assign popcount22_ujfe_core_039 = popcount22_ujfe_core_031 | popcount22_ujfe_core_037;
  assign popcount22_ujfe_core_041 = ~(input_a[17] & input_a[20]);
  assign popcount22_ujfe_core_042 = ~(input_a[11] & input_a[10]);
  assign popcount22_ujfe_core_043 = input_a[10] & input_a[2];
  assign popcount22_ujfe_core_044 = input_a[13] ^ input_a[3];
  assign popcount22_ujfe_core_046_not = ~input_a[17];
  assign popcount22_ujfe_core_047 = ~(input_a[1] ^ input_a[5]);
  assign popcount22_ujfe_core_048 = ~(input_a[11] ^ input_a[4]);
  assign popcount22_ujfe_core_049 = ~(input_a[0] ^ input_a[8]);
  assign popcount22_ujfe_core_051 = ~(input_a[14] ^ input_a[7]);
  assign popcount22_ujfe_core_052 = ~input_a[20];
  assign popcount22_ujfe_core_053 = input_a[9] & input_a[17];
  assign popcount22_ujfe_core_054 = input_a[9] | input_a[21];
  assign popcount22_ujfe_core_055 = ~input_a[3];
  assign popcount22_ujfe_core_056 = ~(input_a[14] ^ input_a[8]);
  assign popcount22_ujfe_core_057 = input_a[10] & input_a[4];
  assign popcount22_ujfe_core_059 = ~(input_a[6] & input_a[4]);
  assign popcount22_ujfe_core_060 = input_a[18] | input_a[4];
  assign popcount22_ujfe_core_062 = input_a[21] & input_a[2];
  assign popcount22_ujfe_core_063 = ~input_a[3];
  assign popcount22_ujfe_core_064 = ~(input_a[13] ^ input_a[18]);
  assign popcount22_ujfe_core_065 = input_a[8] ^ input_a[2];
  assign popcount22_ujfe_core_066 = ~input_a[1];
  assign popcount22_ujfe_core_067 = ~(input_a[20] & input_a[4]);
  assign popcount22_ujfe_core_068 = input_a[19] ^ input_a[21];
  assign popcount22_ujfe_core_069 = ~(input_a[8] ^ input_a[17]);
  assign popcount22_ujfe_core_070 = input_a[14] & input_a[16];
  assign popcount22_ujfe_core_072 = ~(input_a[16] | input_a[15]);
  assign popcount22_ujfe_core_075 = input_a[6] ^ input_a[2];
  assign popcount22_ujfe_core_081 = input_a[15] & input_a[3];
  assign popcount22_ujfe_core_083 = input_a[18] & input_a[20];
  assign popcount22_ujfe_core_084 = ~(input_a[0] ^ input_a[19]);
  assign popcount22_ujfe_core_085 = input_a[2] & input_a[7];
  assign popcount22_ujfe_core_090 = ~input_a[20];
  assign popcount22_ujfe_core_091 = input_a[17] & input_a[3];
  assign popcount22_ujfe_core_092 = popcount22_ujfe_core_083 ^ popcount22_ujfe_core_085;
  assign popcount22_ujfe_core_093 = popcount22_ujfe_core_083 & popcount22_ujfe_core_085;
  assign popcount22_ujfe_core_094 = popcount22_ujfe_core_092 ^ popcount22_ujfe_core_091;
  assign popcount22_ujfe_core_095 = popcount22_ujfe_core_092 & popcount22_ujfe_core_091;
  assign popcount22_ujfe_core_096 = popcount22_ujfe_core_093 | popcount22_ujfe_core_095;
  assign popcount22_ujfe_core_098 = input_a[12] | input_a[17];
  assign popcount22_ujfe_core_101 = input_a[12] & input_a[16];
  assign popcount22_ujfe_core_102 = ~(input_a[9] & input_a[5]);
  assign popcount22_ujfe_core_103 = ~(input_a[14] | input_a[5]);
  assign popcount22_ujfe_core_104 = ~input_a[6];
  assign popcount22_ujfe_core_107 = input_a[20] | input_a[5];
  assign popcount22_ujfe_core_108 = ~(input_a[17] | input_a[10]);
  assign popcount22_ujfe_core_109 = input_a[14] ^ input_a[8];
  assign popcount22_ujfe_core_111 = input_a[19] & input_a[0];
  assign popcount22_ujfe_core_112 = input_a[1] & input_a[14];
  assign popcount22_ujfe_core_115 = input_a[8] ^ popcount22_ujfe_core_112;
  assign popcount22_ujfe_core_116 = input_a[8] & popcount22_ujfe_core_112;
  assign popcount22_ujfe_core_119 = ~(input_a[9] ^ input_a[16]);
  assign popcount22_ujfe_core_121 = ~(input_a[0] ^ input_a[8]);
  assign popcount22_ujfe_core_122 = input_a[13] & input_a[21];
  assign popcount22_ujfe_core_123 = input_a[10] | input_a[12];
  assign popcount22_ujfe_core_124 = input_a[21] & input_a[11];
  assign popcount22_ujfe_core_125 = popcount22_ujfe_core_094 | popcount22_ujfe_core_115;
  assign popcount22_ujfe_core_126 = popcount22_ujfe_core_094 & popcount22_ujfe_core_115;
  assign popcount22_ujfe_core_127 = input_a[18] | input_a[4];
  assign popcount22_ujfe_core_128 = popcount22_ujfe_core_125 & popcount22_ujfe_core_124;
  assign popcount22_ujfe_core_129 = popcount22_ujfe_core_126 | popcount22_ujfe_core_128;
  assign popcount22_ujfe_core_130 = popcount22_ujfe_core_096 ^ popcount22_ujfe_core_116;
  assign popcount22_ujfe_core_131 = popcount22_ujfe_core_096 & popcount22_ujfe_core_116;
  assign popcount22_ujfe_core_132 = popcount22_ujfe_core_130 ^ popcount22_ujfe_core_129;
  assign popcount22_ujfe_core_133 = popcount22_ujfe_core_130 & popcount22_ujfe_core_129;
  assign popcount22_ujfe_core_134 = popcount22_ujfe_core_131 | popcount22_ujfe_core_133;
  assign popcount22_ujfe_core_141 = ~(input_a[2] | input_a[18]);
  assign popcount22_ujfe_core_142 = ~(input_a[6] & input_a[4]);
  assign popcount22_ujfe_core_143 = input_a[21] ^ input_a[19];
  assign popcount22_ujfe_core_144 = ~(input_a[13] | input_a[9]);
  assign popcount22_ujfe_core_145 = ~popcount22_ujfe_core_142;
  assign popcount22_ujfe_core_146 = input_a[15] | input_a[7];
  assign popcount22_ujfe_core_147_not = ~input_a[17];
  assign popcount22_ujfe_core_150 = ~(input_a[8] & input_a[3]);
  assign popcount22_ujfe_core_152 = popcount22_ujfe_core_039 ^ popcount22_ujfe_core_134;
  assign popcount22_ujfe_core_153 = popcount22_ujfe_core_039 & popcount22_ujfe_core_134;
  assign popcount22_ujfe_core_154 = popcount22_ujfe_core_152 ^ popcount22_ujfe_core_132;
  assign popcount22_ujfe_core_155 = popcount22_ujfe_core_152 & popcount22_ujfe_core_132;
  assign popcount22_ujfe_core_156 = popcount22_ujfe_core_153 | popcount22_ujfe_core_155;
  assign popcount22_ujfe_core_158 = ~input_a[16];
  assign popcount22_ujfe_core_159 = input_a[13] & input_a[9];
  assign popcount22_ujfe_core_161 = input_a[16] & input_a[5];

  assign popcount22_ujfe_out[0] = input_a[5];
  assign popcount22_ujfe_out[1] = popcount22_ujfe_core_142;
  assign popcount22_ujfe_out[2] = popcount22_ujfe_core_145;
  assign popcount22_ujfe_out[3] = popcount22_ujfe_core_154;
  assign popcount22_ujfe_out[4] = popcount22_ujfe_core_156;
endmodule