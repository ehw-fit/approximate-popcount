// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5004
// WCE=43.0
// EP=0.999746%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount47_31yb(input [46:0] input_a, output [5:0] popcount47_31yb_out);
  wire popcount47_31yb_core_049;
  wire popcount47_31yb_core_050;
  wire popcount47_31yb_core_051;
  wire popcount47_31yb_core_053;
  wire popcount47_31yb_core_054;
  wire popcount47_31yb_core_055;
  wire popcount47_31yb_core_056;
  wire popcount47_31yb_core_059;
  wire popcount47_31yb_core_060;
  wire popcount47_31yb_core_061;
  wire popcount47_31yb_core_062;
  wire popcount47_31yb_core_063;
  wire popcount47_31yb_core_064;
  wire popcount47_31yb_core_066;
  wire popcount47_31yb_core_068;
  wire popcount47_31yb_core_069;
  wire popcount47_31yb_core_070;
  wire popcount47_31yb_core_071;
  wire popcount47_31yb_core_072;
  wire popcount47_31yb_core_073;
  wire popcount47_31yb_core_076;
  wire popcount47_31yb_core_077;
  wire popcount47_31yb_core_078;
  wire popcount47_31yb_core_079;
  wire popcount47_31yb_core_080;
  wire popcount47_31yb_core_081;
  wire popcount47_31yb_core_083;
  wire popcount47_31yb_core_085;
  wire popcount47_31yb_core_086;
  wire popcount47_31yb_core_087;
  wire popcount47_31yb_core_089;
  wire popcount47_31yb_core_090;
  wire popcount47_31yb_core_092;
  wire popcount47_31yb_core_094;
  wire popcount47_31yb_core_095;
  wire popcount47_31yb_core_096;
  wire popcount47_31yb_core_097;
  wire popcount47_31yb_core_099;
  wire popcount47_31yb_core_100;
  wire popcount47_31yb_core_101;
  wire popcount47_31yb_core_103;
  wire popcount47_31yb_core_105;
  wire popcount47_31yb_core_107;
  wire popcount47_31yb_core_109;
  wire popcount47_31yb_core_110_not;
  wire popcount47_31yb_core_114;
  wire popcount47_31yb_core_115;
  wire popcount47_31yb_core_116;
  wire popcount47_31yb_core_117;
  wire popcount47_31yb_core_120;
  wire popcount47_31yb_core_121;
  wire popcount47_31yb_core_123;
  wire popcount47_31yb_core_124;
  wire popcount47_31yb_core_125;
  wire popcount47_31yb_core_128;
  wire popcount47_31yb_core_129;
  wire popcount47_31yb_core_130;
  wire popcount47_31yb_core_131;
  wire popcount47_31yb_core_132;
  wire popcount47_31yb_core_133;
  wire popcount47_31yb_core_136;
  wire popcount47_31yb_core_137;
  wire popcount47_31yb_core_138;
  wire popcount47_31yb_core_139;
  wire popcount47_31yb_core_140;
  wire popcount47_31yb_core_141;
  wire popcount47_31yb_core_142;
  wire popcount47_31yb_core_143;
  wire popcount47_31yb_core_144;
  wire popcount47_31yb_core_146;
  wire popcount47_31yb_core_147;
  wire popcount47_31yb_core_148;
  wire popcount47_31yb_core_149;
  wire popcount47_31yb_core_150;
  wire popcount47_31yb_core_152;
  wire popcount47_31yb_core_153;
  wire popcount47_31yb_core_154;
  wire popcount47_31yb_core_155;
  wire popcount47_31yb_core_158;
  wire popcount47_31yb_core_159;
  wire popcount47_31yb_core_161;
  wire popcount47_31yb_core_162;
  wire popcount47_31yb_core_163;
  wire popcount47_31yb_core_164;
  wire popcount47_31yb_core_167;
  wire popcount47_31yb_core_168;
  wire popcount47_31yb_core_169;
  wire popcount47_31yb_core_170;
  wire popcount47_31yb_core_172;
  wire popcount47_31yb_core_173;
  wire popcount47_31yb_core_174;
  wire popcount47_31yb_core_175;
  wire popcount47_31yb_core_179;
  wire popcount47_31yb_core_181;
  wire popcount47_31yb_core_184;
  wire popcount47_31yb_core_185;
  wire popcount47_31yb_core_186;
  wire popcount47_31yb_core_188;
  wire popcount47_31yb_core_189;
  wire popcount47_31yb_core_190;
  wire popcount47_31yb_core_191;
  wire popcount47_31yb_core_192;
  wire popcount47_31yb_core_193;
  wire popcount47_31yb_core_194;
  wire popcount47_31yb_core_197;
  wire popcount47_31yb_core_198;
  wire popcount47_31yb_core_200;
  wire popcount47_31yb_core_202;
  wire popcount47_31yb_core_205;
  wire popcount47_31yb_core_206;
  wire popcount47_31yb_core_207;
  wire popcount47_31yb_core_208;
  wire popcount47_31yb_core_209;
  wire popcount47_31yb_core_210;
  wire popcount47_31yb_core_211;
  wire popcount47_31yb_core_212;
  wire popcount47_31yb_core_215;
  wire popcount47_31yb_core_216;
  wire popcount47_31yb_core_217;
  wire popcount47_31yb_core_218_not;
  wire popcount47_31yb_core_219;
  wire popcount47_31yb_core_220;
  wire popcount47_31yb_core_221;
  wire popcount47_31yb_core_223;
  wire popcount47_31yb_core_225;
  wire popcount47_31yb_core_226;
  wire popcount47_31yb_core_229;
  wire popcount47_31yb_core_231;
  wire popcount47_31yb_core_232;
  wire popcount47_31yb_core_233;
  wire popcount47_31yb_core_234;
  wire popcount47_31yb_core_235;
  wire popcount47_31yb_core_238;
  wire popcount47_31yb_core_240;
  wire popcount47_31yb_core_242;
  wire popcount47_31yb_core_243;
  wire popcount47_31yb_core_244;
  wire popcount47_31yb_core_245;
  wire popcount47_31yb_core_247;
  wire popcount47_31yb_core_248;
  wire popcount47_31yb_core_249;
  wire popcount47_31yb_core_250;
  wire popcount47_31yb_core_254;
  wire popcount47_31yb_core_257;
  wire popcount47_31yb_core_258;
  wire popcount47_31yb_core_259;
  wire popcount47_31yb_core_260;
  wire popcount47_31yb_core_263;
  wire popcount47_31yb_core_264;
  wire popcount47_31yb_core_266;
  wire popcount47_31yb_core_267;
  wire popcount47_31yb_core_268;
  wire popcount47_31yb_core_269;
  wire popcount47_31yb_core_270;
  wire popcount47_31yb_core_271;
  wire popcount47_31yb_core_272;
  wire popcount47_31yb_core_273;
  wire popcount47_31yb_core_274;
  wire popcount47_31yb_core_275;
  wire popcount47_31yb_core_276;
  wire popcount47_31yb_core_280;
  wire popcount47_31yb_core_281;
  wire popcount47_31yb_core_282;
  wire popcount47_31yb_core_283;
  wire popcount47_31yb_core_284;
  wire popcount47_31yb_core_286;
  wire popcount47_31yb_core_288;
  wire popcount47_31yb_core_289;
  wire popcount47_31yb_core_291;
  wire popcount47_31yb_core_292;
  wire popcount47_31yb_core_293;
  wire popcount47_31yb_core_294;
  wire popcount47_31yb_core_295;
  wire popcount47_31yb_core_296;
  wire popcount47_31yb_core_301;
  wire popcount47_31yb_core_302;
  wire popcount47_31yb_core_303;
  wire popcount47_31yb_core_304;
  wire popcount47_31yb_core_305;
  wire popcount47_31yb_core_312;
  wire popcount47_31yb_core_313;
  wire popcount47_31yb_core_317;
  wire popcount47_31yb_core_318;
  wire popcount47_31yb_core_320;
  wire popcount47_31yb_core_321;
  wire popcount47_31yb_core_322;
  wire popcount47_31yb_core_323;
  wire popcount47_31yb_core_324;
  wire popcount47_31yb_core_326;
  wire popcount47_31yb_core_327;
  wire popcount47_31yb_core_328;
  wire popcount47_31yb_core_330;
  wire popcount47_31yb_core_331;
  wire popcount47_31yb_core_332;
  wire popcount47_31yb_core_333;
  wire popcount47_31yb_core_334;
  wire popcount47_31yb_core_335;
  wire popcount47_31yb_core_336_not;
  wire popcount47_31yb_core_337;
  wire popcount47_31yb_core_338;
  wire popcount47_31yb_core_340;
  wire popcount47_31yb_core_341;
  wire popcount47_31yb_core_347;
  wire popcount47_31yb_core_349;
  wire popcount47_31yb_core_350;
  wire popcount47_31yb_core_352;
  wire popcount47_31yb_core_353;
  wire popcount47_31yb_core_354;
  wire popcount47_31yb_core_355;
  wire popcount47_31yb_core_356;
  wire popcount47_31yb_core_357;
  wire popcount47_31yb_core_358;
  wire popcount47_31yb_core_359;
  wire popcount47_31yb_core_360;
  wire popcount47_31yb_core_361;
  wire popcount47_31yb_core_362;
  wire popcount47_31yb_core_363;
  wire popcount47_31yb_core_364;
  wire popcount47_31yb_core_365;
  wire popcount47_31yb_core_366;
  wire popcount47_31yb_core_368;
  wire popcount47_31yb_core_369;
  wire popcount47_31yb_core_370;
  wire popcount47_31yb_core_372;

  assign popcount47_31yb_core_049 = ~(input_a[44] ^ input_a[46]);
  assign popcount47_31yb_core_050 = input_a[2] ^ input_a[14];
  assign popcount47_31yb_core_051 = input_a[13] | input_a[36];
  assign popcount47_31yb_core_053 = input_a[39] ^ input_a[33];
  assign popcount47_31yb_core_054 = ~input_a[16];
  assign popcount47_31yb_core_055 = ~(input_a[11] | input_a[9]);
  assign popcount47_31yb_core_056 = input_a[11] & input_a[14];
  assign popcount47_31yb_core_059 = ~(input_a[17] & input_a[41]);
  assign popcount47_31yb_core_060 = input_a[19] & input_a[34];
  assign popcount47_31yb_core_061 = input_a[45] ^ input_a[25];
  assign popcount47_31yb_core_062 = input_a[23] ^ input_a[20];
  assign popcount47_31yb_core_063 = ~(input_a[40] | input_a[6]);
  assign popcount47_31yb_core_064 = ~input_a[17];
  assign popcount47_31yb_core_066 = ~(input_a[14] ^ input_a[46]);
  assign popcount47_31yb_core_068 = ~(input_a[23] & input_a[12]);
  assign popcount47_31yb_core_069 = ~(input_a[21] ^ input_a[8]);
  assign popcount47_31yb_core_070 = ~input_a[6];
  assign popcount47_31yb_core_071 = input_a[33] & input_a[4];
  assign popcount47_31yb_core_072 = input_a[40] & input_a[10];
  assign popcount47_31yb_core_073 = input_a[3] & input_a[31];
  assign popcount47_31yb_core_076 = ~(input_a[31] ^ input_a[7]);
  assign popcount47_31yb_core_077 = input_a[15] | input_a[17];
  assign popcount47_31yb_core_078 = ~input_a[30];
  assign popcount47_31yb_core_079 = input_a[8] ^ input_a[38];
  assign popcount47_31yb_core_080 = input_a[3] | input_a[2];
  assign popcount47_31yb_core_081 = ~(input_a[0] ^ input_a[42]);
  assign popcount47_31yb_core_083 = input_a[39] ^ input_a[31];
  assign popcount47_31yb_core_085 = ~input_a[12];
  assign popcount47_31yb_core_086 = input_a[20] ^ input_a[9];
  assign popcount47_31yb_core_087 = input_a[46] | input_a[22];
  assign popcount47_31yb_core_089 = ~(input_a[8] ^ input_a[14]);
  assign popcount47_31yb_core_090 = ~(input_a[34] & input_a[22]);
  assign popcount47_31yb_core_092 = ~(input_a[2] ^ input_a[46]);
  assign popcount47_31yb_core_094 = input_a[7] | input_a[1];
  assign popcount47_31yb_core_095 = input_a[20] | input_a[3];
  assign popcount47_31yb_core_096 = input_a[22] | input_a[33];
  assign popcount47_31yb_core_097 = ~(input_a[34] | input_a[32]);
  assign popcount47_31yb_core_099 = input_a[10] | input_a[7];
  assign popcount47_31yb_core_100 = input_a[22] | input_a[28];
  assign popcount47_31yb_core_101 = ~(input_a[24] | input_a[12]);
  assign popcount47_31yb_core_103 = ~(input_a[9] ^ input_a[6]);
  assign popcount47_31yb_core_105 = ~input_a[34];
  assign popcount47_31yb_core_107 = ~(input_a[20] | input_a[44]);
  assign popcount47_31yb_core_109 = input_a[36] ^ input_a[27];
  assign popcount47_31yb_core_110_not = ~input_a[2];
  assign popcount47_31yb_core_114 = ~(input_a[39] ^ input_a[40]);
  assign popcount47_31yb_core_115 = ~input_a[9];
  assign popcount47_31yb_core_116 = ~(input_a[14] & input_a[13]);
  assign popcount47_31yb_core_117 = ~(input_a[29] ^ input_a[21]);
  assign popcount47_31yb_core_120 = ~input_a[8];
  assign popcount47_31yb_core_121 = ~input_a[44];
  assign popcount47_31yb_core_123 = ~(input_a[8] | input_a[38]);
  assign popcount47_31yb_core_124 = input_a[23] | input_a[42];
  assign popcount47_31yb_core_125 = input_a[6] | input_a[44];
  assign popcount47_31yb_core_128 = ~(input_a[28] ^ input_a[10]);
  assign popcount47_31yb_core_129 = ~input_a[34];
  assign popcount47_31yb_core_130 = input_a[31] & input_a[25];
  assign popcount47_31yb_core_131 = ~(input_a[22] & input_a[4]);
  assign popcount47_31yb_core_132 = input_a[22] | input_a[10];
  assign popcount47_31yb_core_133 = ~(input_a[38] ^ input_a[29]);
  assign popcount47_31yb_core_136 = ~input_a[20];
  assign popcount47_31yb_core_137 = input_a[29] | input_a[21];
  assign popcount47_31yb_core_138 = input_a[39] & input_a[23];
  assign popcount47_31yb_core_139 = input_a[4] ^ input_a[36];
  assign popcount47_31yb_core_140 = input_a[30] ^ input_a[45];
  assign popcount47_31yb_core_141 = ~(input_a[8] | input_a[36]);
  assign popcount47_31yb_core_142 = ~(input_a[31] | input_a[21]);
  assign popcount47_31yb_core_143 = ~(input_a[26] & input_a[17]);
  assign popcount47_31yb_core_144 = input_a[36] & input_a[39];
  assign popcount47_31yb_core_146 = input_a[24] ^ input_a[36];
  assign popcount47_31yb_core_147 = ~input_a[46];
  assign popcount47_31yb_core_148 = ~(input_a[31] & input_a[46]);
  assign popcount47_31yb_core_149 = ~(input_a[12] ^ input_a[31]);
  assign popcount47_31yb_core_150 = ~input_a[35];
  assign popcount47_31yb_core_152 = ~(input_a[44] | input_a[36]);
  assign popcount47_31yb_core_153 = ~input_a[40];
  assign popcount47_31yb_core_154 = ~input_a[39];
  assign popcount47_31yb_core_155 = input_a[21] | input_a[28];
  assign popcount47_31yb_core_158 = ~(input_a[18] ^ input_a[13]);
  assign popcount47_31yb_core_159 = ~(input_a[6] ^ input_a[18]);
  assign popcount47_31yb_core_161 = input_a[7] | input_a[18];
  assign popcount47_31yb_core_162 = input_a[23] & input_a[4];
  assign popcount47_31yb_core_163 = ~(input_a[15] & input_a[41]);
  assign popcount47_31yb_core_164 = ~(input_a[28] & input_a[15]);
  assign popcount47_31yb_core_167 = ~(input_a[32] ^ input_a[0]);
  assign popcount47_31yb_core_168 = input_a[4] | input_a[35];
  assign popcount47_31yb_core_169 = ~(input_a[4] | input_a[0]);
  assign popcount47_31yb_core_170 = ~(input_a[4] ^ input_a[41]);
  assign popcount47_31yb_core_172 = ~(input_a[16] | input_a[9]);
  assign popcount47_31yb_core_173 = ~input_a[21];
  assign popcount47_31yb_core_174 = input_a[3] | input_a[6];
  assign popcount47_31yb_core_175 = ~(input_a[7] ^ input_a[38]);
  assign popcount47_31yb_core_179 = input_a[15] & input_a[8];
  assign popcount47_31yb_core_181 = ~(input_a[43] & input_a[39]);
  assign popcount47_31yb_core_184 = ~(input_a[8] | input_a[8]);
  assign popcount47_31yb_core_185 = ~(input_a[28] | input_a[45]);
  assign popcount47_31yb_core_186 = input_a[3] & input_a[42];
  assign popcount47_31yb_core_188 = input_a[30] ^ input_a[40];
  assign popcount47_31yb_core_189 = ~(input_a[1] | input_a[3]);
  assign popcount47_31yb_core_190 = ~(input_a[34] ^ input_a[5]);
  assign popcount47_31yb_core_191 = ~input_a[38];
  assign popcount47_31yb_core_192 = input_a[36] | input_a[28];
  assign popcount47_31yb_core_193 = input_a[31] | input_a[15];
  assign popcount47_31yb_core_194 = input_a[4] | input_a[21];
  assign popcount47_31yb_core_197 = input_a[29] ^ input_a[3];
  assign popcount47_31yb_core_198 = input_a[22] ^ input_a[19];
  assign popcount47_31yb_core_200 = input_a[6] ^ input_a[0];
  assign popcount47_31yb_core_202 = ~(input_a[40] ^ input_a[25]);
  assign popcount47_31yb_core_205 = ~(input_a[29] | input_a[4]);
  assign popcount47_31yb_core_206 = input_a[4] & input_a[36];
  assign popcount47_31yb_core_207 = input_a[42] | input_a[16];
  assign popcount47_31yb_core_208 = input_a[41] | input_a[12];
  assign popcount47_31yb_core_209 = ~(input_a[42] ^ input_a[4]);
  assign popcount47_31yb_core_210 = ~(input_a[4] & input_a[9]);
  assign popcount47_31yb_core_211 = ~input_a[6];
  assign popcount47_31yb_core_212 = ~input_a[3];
  assign popcount47_31yb_core_215 = ~input_a[43];
  assign popcount47_31yb_core_216 = ~(input_a[18] | input_a[12]);
  assign popcount47_31yb_core_217 = ~(input_a[43] | input_a[19]);
  assign popcount47_31yb_core_218_not = ~input_a[23];
  assign popcount47_31yb_core_219 = ~(input_a[11] | input_a[18]);
  assign popcount47_31yb_core_220 = ~(input_a[8] | input_a[19]);
  assign popcount47_31yb_core_221 = input_a[7] ^ input_a[13];
  assign popcount47_31yb_core_223 = input_a[13] | input_a[43];
  assign popcount47_31yb_core_225 = ~input_a[27];
  assign popcount47_31yb_core_226 = ~input_a[46];
  assign popcount47_31yb_core_229 = input_a[22] | input_a[42];
  assign popcount47_31yb_core_231 = input_a[12] & input_a[14];
  assign popcount47_31yb_core_232 = ~(input_a[16] | input_a[43]);
  assign popcount47_31yb_core_233 = input_a[14] | input_a[0];
  assign popcount47_31yb_core_234 = input_a[14] | input_a[39];
  assign popcount47_31yb_core_235 = ~(input_a[37] | input_a[14]);
  assign popcount47_31yb_core_238 = ~input_a[29];
  assign popcount47_31yb_core_240 = ~(input_a[23] & input_a[23]);
  assign popcount47_31yb_core_242 = input_a[41] ^ input_a[14];
  assign popcount47_31yb_core_243 = input_a[19] & input_a[14];
  assign popcount47_31yb_core_244 = ~input_a[15];
  assign popcount47_31yb_core_245 = ~(input_a[20] ^ input_a[12]);
  assign popcount47_31yb_core_247 = ~(input_a[35] ^ input_a[33]);
  assign popcount47_31yb_core_248 = ~input_a[16];
  assign popcount47_31yb_core_249 = input_a[3] | input_a[7];
  assign popcount47_31yb_core_250 = ~input_a[16];
  assign popcount47_31yb_core_254 = input_a[12] & input_a[21];
  assign popcount47_31yb_core_257 = input_a[6] ^ input_a[28];
  assign popcount47_31yb_core_258 = input_a[2] | input_a[34];
  assign popcount47_31yb_core_259 = input_a[44] ^ input_a[23];
  assign popcount47_31yb_core_260 = ~(input_a[13] ^ input_a[36]);
  assign popcount47_31yb_core_263 = input_a[33] & input_a[0];
  assign popcount47_31yb_core_264 = input_a[31] | input_a[9];
  assign popcount47_31yb_core_266 = ~(input_a[24] ^ input_a[11]);
  assign popcount47_31yb_core_267 = ~(input_a[16] ^ input_a[10]);
  assign popcount47_31yb_core_268 = ~(input_a[34] ^ input_a[24]);
  assign popcount47_31yb_core_269 = ~input_a[16];
  assign popcount47_31yb_core_270 = ~(input_a[8] ^ input_a[30]);
  assign popcount47_31yb_core_271 = ~(input_a[25] | input_a[14]);
  assign popcount47_31yb_core_272 = ~(input_a[38] | input_a[46]);
  assign popcount47_31yb_core_273 = ~input_a[31];
  assign popcount47_31yb_core_274 = ~(input_a[7] ^ input_a[45]);
  assign popcount47_31yb_core_275 = input_a[37] & input_a[44];
  assign popcount47_31yb_core_276 = ~input_a[40];
  assign popcount47_31yb_core_280 = ~(input_a[14] & input_a[34]);
  assign popcount47_31yb_core_281 = input_a[21] & input_a[22];
  assign popcount47_31yb_core_282 = input_a[41] | input_a[34];
  assign popcount47_31yb_core_283 = ~input_a[6];
  assign popcount47_31yb_core_284 = input_a[21] | input_a[33];
  assign popcount47_31yb_core_286 = ~(input_a[20] ^ input_a[19]);
  assign popcount47_31yb_core_288 = input_a[5] ^ input_a[5];
  assign popcount47_31yb_core_289 = ~(input_a[36] | input_a[10]);
  assign popcount47_31yb_core_291 = input_a[22] ^ input_a[16];
  assign popcount47_31yb_core_292 = ~input_a[22];
  assign popcount47_31yb_core_293 = input_a[39] | input_a[15];
  assign popcount47_31yb_core_294 = input_a[43] | input_a[3];
  assign popcount47_31yb_core_295 = input_a[27] & input_a[19];
  assign popcount47_31yb_core_296 = ~(input_a[18] | input_a[20]);
  assign popcount47_31yb_core_301 = input_a[8] | input_a[13];
  assign popcount47_31yb_core_302 = ~(input_a[17] | input_a[9]);
  assign popcount47_31yb_core_303 = ~(input_a[21] ^ input_a[7]);
  assign popcount47_31yb_core_304 = ~input_a[46];
  assign popcount47_31yb_core_305 = ~(input_a[15] & input_a[44]);
  assign popcount47_31yb_core_312 = ~(input_a[39] & input_a[3]);
  assign popcount47_31yb_core_313 = input_a[27] ^ input_a[11];
  assign popcount47_31yb_core_317 = ~(input_a[12] | input_a[13]);
  assign popcount47_31yb_core_318 = ~input_a[17];
  assign popcount47_31yb_core_320 = input_a[0] & input_a[5];
  assign popcount47_31yb_core_321 = input_a[29] ^ input_a[29];
  assign popcount47_31yb_core_322 = input_a[27] ^ input_a[32];
  assign popcount47_31yb_core_323 = ~(input_a[24] ^ input_a[25]);
  assign popcount47_31yb_core_324 = ~(input_a[3] ^ input_a[10]);
  assign popcount47_31yb_core_326 = input_a[5] ^ input_a[12];
  assign popcount47_31yb_core_327 = input_a[27] ^ input_a[2];
  assign popcount47_31yb_core_328 = ~(input_a[27] & input_a[26]);
  assign popcount47_31yb_core_330 = ~(input_a[7] ^ input_a[23]);
  assign popcount47_31yb_core_331 = ~(input_a[10] | input_a[19]);
  assign popcount47_31yb_core_332 = ~(input_a[35] | input_a[44]);
  assign popcount47_31yb_core_333 = ~(input_a[25] | input_a[16]);
  assign popcount47_31yb_core_334 = ~(input_a[32] & input_a[4]);
  assign popcount47_31yb_core_335 = input_a[4] ^ input_a[32];
  assign popcount47_31yb_core_336_not = ~input_a[35];
  assign popcount47_31yb_core_337 = ~input_a[25];
  assign popcount47_31yb_core_338 = ~(input_a[34] ^ input_a[45]);
  assign popcount47_31yb_core_340 = input_a[19] | input_a[21];
  assign popcount47_31yb_core_341 = ~(input_a[28] | input_a[17]);
  assign popcount47_31yb_core_347 = ~(input_a[14] & input_a[25]);
  assign popcount47_31yb_core_349 = input_a[23] & input_a[41];
  assign popcount47_31yb_core_350 = ~(input_a[14] | input_a[1]);
  assign popcount47_31yb_core_352 = ~(input_a[45] | input_a[40]);
  assign popcount47_31yb_core_353 = input_a[35] | input_a[2];
  assign popcount47_31yb_core_354 = ~(input_a[37] & input_a[39]);
  assign popcount47_31yb_core_355 = input_a[6] ^ input_a[32];
  assign popcount47_31yb_core_356 = ~input_a[28];
  assign popcount47_31yb_core_357 = ~(input_a[22] ^ input_a[38]);
  assign popcount47_31yb_core_358 = ~input_a[14];
  assign popcount47_31yb_core_359 = input_a[23] & input_a[14];
  assign popcount47_31yb_core_360 = ~(input_a[19] ^ input_a[11]);
  assign popcount47_31yb_core_361 = ~(input_a[7] & input_a[35]);
  assign popcount47_31yb_core_362 = ~(input_a[29] & input_a[27]);
  assign popcount47_31yb_core_363 = ~(input_a[37] | input_a[28]);
  assign popcount47_31yb_core_364 = ~(input_a[22] ^ input_a[33]);
  assign popcount47_31yb_core_365 = ~(input_a[40] & input_a[43]);
  assign popcount47_31yb_core_366 = input_a[44] & input_a[23];
  assign popcount47_31yb_core_368 = ~(input_a[32] | input_a[38]);
  assign popcount47_31yb_core_369 = ~input_a[0];
  assign popcount47_31yb_core_370 = ~input_a[34];
  assign popcount47_31yb_core_372 = ~input_a[22];

  assign popcount47_31yb_out[0] = input_a[15];
  assign popcount47_31yb_out[1] = 1'b0;
  assign popcount47_31yb_out[2] = input_a[39];
  assign popcount47_31yb_out[3] = input_a[37];
  assign popcount47_31yb_out[4] = 1'b0;
  assign popcount47_31yb_out[5] = input_a[13];
endmodule