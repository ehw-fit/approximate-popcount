// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.90772
// WCE=24.0
// EP=0.929838%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_j1nz(input [34:0] input_a, output [5:0] popcount35_j1nz_out);
  wire popcount35_j1nz_core_037;
  wire popcount35_j1nz_core_038;
  wire popcount35_j1nz_core_039;
  wire popcount35_j1nz_core_040;
  wire popcount35_j1nz_core_041;
  wire popcount35_j1nz_core_043;
  wire popcount35_j1nz_core_044;
  wire popcount35_j1nz_core_045;
  wire popcount35_j1nz_core_046;
  wire popcount35_j1nz_core_047;
  wire popcount35_j1nz_core_048;
  wire popcount35_j1nz_core_049;
  wire popcount35_j1nz_core_052;
  wire popcount35_j1nz_core_053;
  wire popcount35_j1nz_core_054;
  wire popcount35_j1nz_core_055;
  wire popcount35_j1nz_core_056;
  wire popcount35_j1nz_core_057;
  wire popcount35_j1nz_core_061;
  wire popcount35_j1nz_core_063;
  wire popcount35_j1nz_core_064;
  wire popcount35_j1nz_core_066;
  wire popcount35_j1nz_core_067;
  wire popcount35_j1nz_core_069;
  wire popcount35_j1nz_core_070;
  wire popcount35_j1nz_core_072;
  wire popcount35_j1nz_core_076;
  wire popcount35_j1nz_core_077;
  wire popcount35_j1nz_core_079_not;
  wire popcount35_j1nz_core_080;
  wire popcount35_j1nz_core_081;
  wire popcount35_j1nz_core_082;
  wire popcount35_j1nz_core_083;
  wire popcount35_j1nz_core_084;
  wire popcount35_j1nz_core_085;
  wire popcount35_j1nz_core_090;
  wire popcount35_j1nz_core_093;
  wire popcount35_j1nz_core_097;
  wire popcount35_j1nz_core_102;
  wire popcount35_j1nz_core_105;
  wire popcount35_j1nz_core_108;
  wire popcount35_j1nz_core_109;
  wire popcount35_j1nz_core_110;
  wire popcount35_j1nz_core_111;
  wire popcount35_j1nz_core_112;
  wire popcount35_j1nz_core_115;
  wire popcount35_j1nz_core_116;
  wire popcount35_j1nz_core_120;
  wire popcount35_j1nz_core_123_not;
  wire popcount35_j1nz_core_125;
  wire popcount35_j1nz_core_126;
  wire popcount35_j1nz_core_128;
  wire popcount35_j1nz_core_129;
  wire popcount35_j1nz_core_131;
  wire popcount35_j1nz_core_132;
  wire popcount35_j1nz_core_134;
  wire popcount35_j1nz_core_137;
  wire popcount35_j1nz_core_138;
  wire popcount35_j1nz_core_143;
  wire popcount35_j1nz_core_145;
  wire popcount35_j1nz_core_146;
  wire popcount35_j1nz_core_147;
  wire popcount35_j1nz_core_150;
  wire popcount35_j1nz_core_151;
  wire popcount35_j1nz_core_152;
  wire popcount35_j1nz_core_153;
  wire popcount35_j1nz_core_155;
  wire popcount35_j1nz_core_159;
  wire popcount35_j1nz_core_160;
  wire popcount35_j1nz_core_161;
  wire popcount35_j1nz_core_162;
  wire popcount35_j1nz_core_163;
  wire popcount35_j1nz_core_166;
  wire popcount35_j1nz_core_169;
  wire popcount35_j1nz_core_170;
  wire popcount35_j1nz_core_171;
  wire popcount35_j1nz_core_172;
  wire popcount35_j1nz_core_173;
  wire popcount35_j1nz_core_174;
  wire popcount35_j1nz_core_176;
  wire popcount35_j1nz_core_177;
  wire popcount35_j1nz_core_179;
  wire popcount35_j1nz_core_183;
  wire popcount35_j1nz_core_184;
  wire popcount35_j1nz_core_185;
  wire popcount35_j1nz_core_186;
  wire popcount35_j1nz_core_187;
  wire popcount35_j1nz_core_189;
  wire popcount35_j1nz_core_190;
  wire popcount35_j1nz_core_193;
  wire popcount35_j1nz_core_195;
  wire popcount35_j1nz_core_196;
  wire popcount35_j1nz_core_197;
  wire popcount35_j1nz_core_198;
  wire popcount35_j1nz_core_200;
  wire popcount35_j1nz_core_201_not;
  wire popcount35_j1nz_core_202;
  wire popcount35_j1nz_core_204;
  wire popcount35_j1nz_core_205;
  wire popcount35_j1nz_core_206;
  wire popcount35_j1nz_core_208;
  wire popcount35_j1nz_core_209;
  wire popcount35_j1nz_core_214;
  wire popcount35_j1nz_core_217;
  wire popcount35_j1nz_core_218;
  wire popcount35_j1nz_core_220;
  wire popcount35_j1nz_core_221;
  wire popcount35_j1nz_core_223;
  wire popcount35_j1nz_core_224;
  wire popcount35_j1nz_core_227;
  wire popcount35_j1nz_core_229;
  wire popcount35_j1nz_core_230;
  wire popcount35_j1nz_core_231;
  wire popcount35_j1nz_core_233;
  wire popcount35_j1nz_core_234;
  wire popcount35_j1nz_core_235;
  wire popcount35_j1nz_core_237;
  wire popcount35_j1nz_core_238;
  wire popcount35_j1nz_core_240;
  wire popcount35_j1nz_core_242;
  wire popcount35_j1nz_core_243;
  wire popcount35_j1nz_core_245;
  wire popcount35_j1nz_core_246;
  wire popcount35_j1nz_core_247;
  wire popcount35_j1nz_core_249;
  wire popcount35_j1nz_core_250;
  wire popcount35_j1nz_core_252;
  wire popcount35_j1nz_core_254;
  wire popcount35_j1nz_core_255;
  wire popcount35_j1nz_core_256;
  wire popcount35_j1nz_core_257;
  wire popcount35_j1nz_core_259;
  wire popcount35_j1nz_core_260;
  wire popcount35_j1nz_core_261;
  wire popcount35_j1nz_core_262;
  wire popcount35_j1nz_core_263;
  wire popcount35_j1nz_core_264;

  assign popcount35_j1nz_core_037 = ~(input_a[5] | input_a[2]);
  assign popcount35_j1nz_core_038 = ~(input_a[16] ^ input_a[25]);
  assign popcount35_j1nz_core_039 = input_a[31] | input_a[21];
  assign popcount35_j1nz_core_040 = input_a[22] | input_a[32];
  assign popcount35_j1nz_core_041 = ~(input_a[18] | input_a[14]);
  assign popcount35_j1nz_core_043 = input_a[22] | input_a[23];
  assign popcount35_j1nz_core_044 = ~(input_a[34] ^ input_a[30]);
  assign popcount35_j1nz_core_045 = ~(input_a[30] & input_a[4]);
  assign popcount35_j1nz_core_046 = ~(input_a[14] & input_a[31]);
  assign popcount35_j1nz_core_047 = ~input_a[9];
  assign popcount35_j1nz_core_048 = input_a[1] & input_a[21];
  assign popcount35_j1nz_core_049 = input_a[33] & input_a[16];
  assign popcount35_j1nz_core_052 = input_a[2] & input_a[20];
  assign popcount35_j1nz_core_053 = input_a[17] | input_a[28];
  assign popcount35_j1nz_core_054 = input_a[24] & input_a[32];
  assign popcount35_j1nz_core_055 = ~(input_a[33] ^ input_a[1]);
  assign popcount35_j1nz_core_056 = ~(input_a[10] ^ input_a[25]);
  assign popcount35_j1nz_core_057 = ~(input_a[22] & input_a[14]);
  assign popcount35_j1nz_core_061 = ~(input_a[23] ^ input_a[17]);
  assign popcount35_j1nz_core_063 = input_a[30] | input_a[22];
  assign popcount35_j1nz_core_064 = ~(input_a[32] & input_a[21]);
  assign popcount35_j1nz_core_066 = ~input_a[26];
  assign popcount35_j1nz_core_067 = input_a[19] & input_a[6];
  assign popcount35_j1nz_core_069 = ~(input_a[16] ^ input_a[27]);
  assign popcount35_j1nz_core_070 = ~input_a[7];
  assign popcount35_j1nz_core_072 = input_a[21] | input_a[26];
  assign popcount35_j1nz_core_076 = ~(input_a[9] ^ input_a[2]);
  assign popcount35_j1nz_core_077 = ~(input_a[26] | input_a[6]);
  assign popcount35_j1nz_core_079_not = ~input_a[31];
  assign popcount35_j1nz_core_080 = ~input_a[30];
  assign popcount35_j1nz_core_081 = input_a[19] | input_a[20];
  assign popcount35_j1nz_core_082 = ~(input_a[3] & input_a[27]);
  assign popcount35_j1nz_core_083 = input_a[15] | input_a[7];
  assign popcount35_j1nz_core_084 = input_a[19] & input_a[7];
  assign popcount35_j1nz_core_085 = ~(input_a[1] | input_a[12]);
  assign popcount35_j1nz_core_090 = ~(input_a[24] | input_a[9]);
  assign popcount35_j1nz_core_093 = ~(input_a[13] & input_a[22]);
  assign popcount35_j1nz_core_097 = ~(input_a[32] | input_a[14]);
  assign popcount35_j1nz_core_102 = input_a[21] | input_a[28];
  assign popcount35_j1nz_core_105 = ~input_a[15];
  assign popcount35_j1nz_core_108 = input_a[8] ^ input_a[17];
  assign popcount35_j1nz_core_109 = ~(input_a[9] & input_a[6]);
  assign popcount35_j1nz_core_110 = input_a[14] & input_a[12];
  assign popcount35_j1nz_core_111 = input_a[28] | input_a[16];
  assign popcount35_j1nz_core_112 = input_a[8] & input_a[26];
  assign popcount35_j1nz_core_115 = input_a[9] | input_a[0];
  assign popcount35_j1nz_core_116 = ~(input_a[26] ^ input_a[13]);
  assign popcount35_j1nz_core_120 = ~input_a[25];
  assign popcount35_j1nz_core_123_not = ~input_a[31];
  assign popcount35_j1nz_core_125 = ~(input_a[26] & input_a[1]);
  assign popcount35_j1nz_core_126 = input_a[13] ^ input_a[32];
  assign popcount35_j1nz_core_128 = input_a[13] ^ input_a[4];
  assign popcount35_j1nz_core_129 = ~(input_a[23] | input_a[24]);
  assign popcount35_j1nz_core_131 = ~(input_a[29] & input_a[20]);
  assign popcount35_j1nz_core_132 = ~input_a[5];
  assign popcount35_j1nz_core_134 = input_a[14] ^ input_a[29];
  assign popcount35_j1nz_core_137 = input_a[24] ^ input_a[28];
  assign popcount35_j1nz_core_138 = input_a[12] & input_a[15];
  assign popcount35_j1nz_core_143 = ~(input_a[31] & input_a[34]);
  assign popcount35_j1nz_core_145 = ~input_a[12];
  assign popcount35_j1nz_core_146 = input_a[31] & input_a[5];
  assign popcount35_j1nz_core_147 = ~(input_a[0] & input_a[0]);
  assign popcount35_j1nz_core_150 = input_a[22] ^ input_a[25];
  assign popcount35_j1nz_core_151 = ~input_a[31];
  assign popcount35_j1nz_core_152 = ~(input_a[14] | input_a[32]);
  assign popcount35_j1nz_core_153 = input_a[17] | input_a[2];
  assign popcount35_j1nz_core_155 = input_a[15] | input_a[1];
  assign popcount35_j1nz_core_159 = input_a[34] | input_a[1];
  assign popcount35_j1nz_core_160 = ~(input_a[27] & input_a[0]);
  assign popcount35_j1nz_core_161 = ~input_a[25];
  assign popcount35_j1nz_core_162 = ~input_a[6];
  assign popcount35_j1nz_core_163 = input_a[8] | input_a[24];
  assign popcount35_j1nz_core_166 = ~(input_a[26] ^ input_a[25]);
  assign popcount35_j1nz_core_169 = ~(input_a[26] & input_a[3]);
  assign popcount35_j1nz_core_170 = ~(input_a[24] & input_a[6]);
  assign popcount35_j1nz_core_171 = input_a[7] | input_a[31];
  assign popcount35_j1nz_core_172 = ~(input_a[14] | input_a[28]);
  assign popcount35_j1nz_core_173 = input_a[19] ^ input_a[30];
  assign popcount35_j1nz_core_174 = ~input_a[31];
  assign popcount35_j1nz_core_176 = input_a[29] | input_a[27];
  assign popcount35_j1nz_core_177 = ~(input_a[21] ^ input_a[5]);
  assign popcount35_j1nz_core_179 = ~input_a[3];
  assign popcount35_j1nz_core_183 = ~(input_a[21] & input_a[26]);
  assign popcount35_j1nz_core_184 = ~input_a[1];
  assign popcount35_j1nz_core_185 = ~(input_a[22] & input_a[34]);
  assign popcount35_j1nz_core_186 = ~(input_a[6] & input_a[7]);
  assign popcount35_j1nz_core_187 = ~(input_a[23] ^ input_a[18]);
  assign popcount35_j1nz_core_189 = input_a[28] ^ input_a[3];
  assign popcount35_j1nz_core_190 = ~input_a[13];
  assign popcount35_j1nz_core_193 = input_a[5] ^ input_a[4];
  assign popcount35_j1nz_core_195 = ~input_a[32];
  assign popcount35_j1nz_core_196 = ~input_a[19];
  assign popcount35_j1nz_core_197 = ~input_a[28];
  assign popcount35_j1nz_core_198 = input_a[31] & input_a[7];
  assign popcount35_j1nz_core_200 = ~(input_a[32] | input_a[13]);
  assign popcount35_j1nz_core_201_not = ~input_a[7];
  assign popcount35_j1nz_core_202 = input_a[31] | input_a[0];
  assign popcount35_j1nz_core_204 = ~input_a[10];
  assign popcount35_j1nz_core_205 = input_a[19] & input_a[23];
  assign popcount35_j1nz_core_206 = ~(input_a[3] ^ input_a[33]);
  assign popcount35_j1nz_core_208 = ~input_a[9];
  assign popcount35_j1nz_core_209 = input_a[30] | input_a[30];
  assign popcount35_j1nz_core_214 = ~(input_a[15] & input_a[30]);
  assign popcount35_j1nz_core_217 = input_a[1] | input_a[20];
  assign popcount35_j1nz_core_218 = input_a[12] | input_a[21];
  assign popcount35_j1nz_core_220 = ~(input_a[28] | input_a[33]);
  assign popcount35_j1nz_core_221 = ~input_a[4];
  assign popcount35_j1nz_core_223 = input_a[34] | input_a[10];
  assign popcount35_j1nz_core_224 = input_a[10] | input_a[3];
  assign popcount35_j1nz_core_227 = input_a[11] ^ input_a[9];
  assign popcount35_j1nz_core_229 = input_a[4] ^ input_a[1];
  assign popcount35_j1nz_core_230 = input_a[2] ^ input_a[10];
  assign popcount35_j1nz_core_231 = ~(input_a[20] & input_a[15]);
  assign popcount35_j1nz_core_233 = input_a[33] & input_a[12];
  assign popcount35_j1nz_core_234 = ~input_a[33];
  assign popcount35_j1nz_core_235 = ~(input_a[26] ^ input_a[0]);
  assign popcount35_j1nz_core_237 = ~(input_a[27] ^ input_a[26]);
  assign popcount35_j1nz_core_238 = ~input_a[7];
  assign popcount35_j1nz_core_240 = ~input_a[22];
  assign popcount35_j1nz_core_242 = ~(input_a[7] & input_a[29]);
  assign popcount35_j1nz_core_243 = input_a[34] & input_a[27];
  assign popcount35_j1nz_core_245 = input_a[29] ^ input_a[17];
  assign popcount35_j1nz_core_246 = ~(input_a[25] | input_a[31]);
  assign popcount35_j1nz_core_247 = ~(input_a[5] ^ input_a[27]);
  assign popcount35_j1nz_core_249 = ~(input_a[3] ^ input_a[20]);
  assign popcount35_j1nz_core_250 = ~(input_a[25] & input_a[31]);
  assign popcount35_j1nz_core_252 = input_a[16] ^ input_a[1];
  assign popcount35_j1nz_core_254 = input_a[4] ^ input_a[18];
  assign popcount35_j1nz_core_255 = ~input_a[6];
  assign popcount35_j1nz_core_256 = ~(input_a[6] & input_a[31]);
  assign popcount35_j1nz_core_257 = ~input_a[19];
  assign popcount35_j1nz_core_259 = input_a[3] ^ input_a[1];
  assign popcount35_j1nz_core_260 = input_a[16] ^ input_a[10];
  assign popcount35_j1nz_core_261 = ~(input_a[16] | input_a[28]);
  assign popcount35_j1nz_core_262 = input_a[21] & input_a[1];
  assign popcount35_j1nz_core_263 = ~(input_a[6] & input_a[32]);
  assign popcount35_j1nz_core_264 = ~(input_a[11] ^ input_a[14]);

  assign popcount35_j1nz_out[0] = input_a[10];
  assign popcount35_j1nz_out[1] = input_a[23];
  assign popcount35_j1nz_out[2] = 1'b0;
  assign popcount35_j1nz_out[3] = input_a[16];
  assign popcount35_j1nz_out[4] = 1'b1;
  assign popcount35_j1nz_out[5] = 1'b0;
endmodule