// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.8044
// WCE=28.0
// EP=0.959077%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_1ht9(input [34:0] input_a, output [5:0] popcount35_1ht9_out);
  wire popcount35_1ht9_core_037;
  wire popcount35_1ht9_core_039;
  wire popcount35_1ht9_core_041;
  wire popcount35_1ht9_core_042;
  wire popcount35_1ht9_core_043;
  wire popcount35_1ht9_core_044;
  wire popcount35_1ht9_core_045;
  wire popcount35_1ht9_core_046;
  wire popcount35_1ht9_core_047;
  wire popcount35_1ht9_core_048;
  wire popcount35_1ht9_core_050;
  wire popcount35_1ht9_core_051;
  wire popcount35_1ht9_core_052;
  wire popcount35_1ht9_core_053;
  wire popcount35_1ht9_core_055;
  wire popcount35_1ht9_core_057;
  wire popcount35_1ht9_core_058;
  wire popcount35_1ht9_core_061;
  wire popcount35_1ht9_core_062;
  wire popcount35_1ht9_core_066;
  wire popcount35_1ht9_core_067;
  wire popcount35_1ht9_core_068;
  wire popcount35_1ht9_core_069;
  wire popcount35_1ht9_core_070;
  wire popcount35_1ht9_core_071;
  wire popcount35_1ht9_core_072;
  wire popcount35_1ht9_core_073;
  wire popcount35_1ht9_core_074;
  wire popcount35_1ht9_core_075;
  wire popcount35_1ht9_core_076;
  wire popcount35_1ht9_core_077;
  wire popcount35_1ht9_core_081;
  wire popcount35_1ht9_core_082;
  wire popcount35_1ht9_core_084;
  wire popcount35_1ht9_core_085;
  wire popcount35_1ht9_core_086;
  wire popcount35_1ht9_core_089;
  wire popcount35_1ht9_core_090;
  wire popcount35_1ht9_core_091;
  wire popcount35_1ht9_core_092;
  wire popcount35_1ht9_core_094;
  wire popcount35_1ht9_core_097;
  wire popcount35_1ht9_core_099;
  wire popcount35_1ht9_core_100;
  wire popcount35_1ht9_core_101;
  wire popcount35_1ht9_core_102;
  wire popcount35_1ht9_core_103;
  wire popcount35_1ht9_core_106;
  wire popcount35_1ht9_core_107;
  wire popcount35_1ht9_core_108;
  wire popcount35_1ht9_core_110;
  wire popcount35_1ht9_core_112;
  wire popcount35_1ht9_core_113;
  wire popcount35_1ht9_core_114;
  wire popcount35_1ht9_core_115;
  wire popcount35_1ht9_core_117;
  wire popcount35_1ht9_core_118;
  wire popcount35_1ht9_core_119;
  wire popcount35_1ht9_core_120;
  wire popcount35_1ht9_core_123;
  wire popcount35_1ht9_core_124;
  wire popcount35_1ht9_core_125;
  wire popcount35_1ht9_core_126;
  wire popcount35_1ht9_core_127;
  wire popcount35_1ht9_core_128;
  wire popcount35_1ht9_core_130;
  wire popcount35_1ht9_core_131;
  wire popcount35_1ht9_core_133;
  wire popcount35_1ht9_core_134;
  wire popcount35_1ht9_core_135;
  wire popcount35_1ht9_core_136;
  wire popcount35_1ht9_core_137;
  wire popcount35_1ht9_core_138;
  wire popcount35_1ht9_core_140;
  wire popcount35_1ht9_core_141;
  wire popcount35_1ht9_core_142;
  wire popcount35_1ht9_core_146;
  wire popcount35_1ht9_core_147;
  wire popcount35_1ht9_core_148;
  wire popcount35_1ht9_core_150;
  wire popcount35_1ht9_core_151;
  wire popcount35_1ht9_core_152;
  wire popcount35_1ht9_core_153;
  wire popcount35_1ht9_core_154;
  wire popcount35_1ht9_core_157;
  wire popcount35_1ht9_core_158;
  wire popcount35_1ht9_core_159;
  wire popcount35_1ht9_core_162;
  wire popcount35_1ht9_core_165;
  wire popcount35_1ht9_core_166;
  wire popcount35_1ht9_core_167;
  wire popcount35_1ht9_core_169;
  wire popcount35_1ht9_core_170;
  wire popcount35_1ht9_core_172;
  wire popcount35_1ht9_core_173;
  wire popcount35_1ht9_core_175;
  wire popcount35_1ht9_core_176;
  wire popcount35_1ht9_core_178;
  wire popcount35_1ht9_core_179_not;
  wire popcount35_1ht9_core_180;
  wire popcount35_1ht9_core_181;
  wire popcount35_1ht9_core_183;
  wire popcount35_1ht9_core_186;
  wire popcount35_1ht9_core_187;
  wire popcount35_1ht9_core_190;
  wire popcount35_1ht9_core_191;
  wire popcount35_1ht9_core_192;
  wire popcount35_1ht9_core_197;
  wire popcount35_1ht9_core_200;
  wire popcount35_1ht9_core_201;
  wire popcount35_1ht9_core_202;
  wire popcount35_1ht9_core_203;
  wire popcount35_1ht9_core_204;
  wire popcount35_1ht9_core_207;
  wire popcount35_1ht9_core_208;
  wire popcount35_1ht9_core_209;
  wire popcount35_1ht9_core_212;
  wire popcount35_1ht9_core_215;
  wire popcount35_1ht9_core_216;
  wire popcount35_1ht9_core_219;
  wire popcount35_1ht9_core_220;
  wire popcount35_1ht9_core_223;
  wire popcount35_1ht9_core_224;
  wire popcount35_1ht9_core_225;
  wire popcount35_1ht9_core_226;
  wire popcount35_1ht9_core_227;
  wire popcount35_1ht9_core_231;
  wire popcount35_1ht9_core_233;
  wire popcount35_1ht9_core_235;
  wire popcount35_1ht9_core_236;
  wire popcount35_1ht9_core_237;
  wire popcount35_1ht9_core_238;
  wire popcount35_1ht9_core_239;
  wire popcount35_1ht9_core_240;
  wire popcount35_1ht9_core_242;
  wire popcount35_1ht9_core_243;
  wire popcount35_1ht9_core_244;
  wire popcount35_1ht9_core_246;
  wire popcount35_1ht9_core_249;
  wire popcount35_1ht9_core_250;
  wire popcount35_1ht9_core_251;
  wire popcount35_1ht9_core_252;
  wire popcount35_1ht9_core_253;
  wire popcount35_1ht9_core_254;
  wire popcount35_1ht9_core_257;
  wire popcount35_1ht9_core_258;
  wire popcount35_1ht9_core_259;
  wire popcount35_1ht9_core_260;
  wire popcount35_1ht9_core_264;

  assign popcount35_1ht9_core_037 = ~(input_a[5] | input_a[32]);
  assign popcount35_1ht9_core_039 = ~(input_a[2] | input_a[25]);
  assign popcount35_1ht9_core_041 = input_a[5] & input_a[32];
  assign popcount35_1ht9_core_042 = ~(input_a[11] | input_a[11]);
  assign popcount35_1ht9_core_043 = input_a[3] | input_a[18];
  assign popcount35_1ht9_core_044 = ~input_a[25];
  assign popcount35_1ht9_core_045 = ~input_a[5];
  assign popcount35_1ht9_core_046 = ~(input_a[25] ^ input_a[27]);
  assign popcount35_1ht9_core_047 = input_a[29] ^ input_a[2];
  assign popcount35_1ht9_core_048 = input_a[0] | input_a[13];
  assign popcount35_1ht9_core_050 = input_a[22] ^ input_a[12];
  assign popcount35_1ht9_core_051 = input_a[29] ^ input_a[17];
  assign popcount35_1ht9_core_052 = input_a[16] ^ input_a[26];
  assign popcount35_1ht9_core_053 = ~(input_a[2] ^ input_a[10]);
  assign popcount35_1ht9_core_055 = input_a[21] & input_a[17];
  assign popcount35_1ht9_core_057 = input_a[9] | input_a[10];
  assign popcount35_1ht9_core_058 = input_a[13] & input_a[11];
  assign popcount35_1ht9_core_061 = input_a[32] ^ input_a[7];
  assign popcount35_1ht9_core_062 = input_a[18] | input_a[22];
  assign popcount35_1ht9_core_066 = ~input_a[12];
  assign popcount35_1ht9_core_067 = ~(input_a[12] & input_a[13]);
  assign popcount35_1ht9_core_068 = input_a[24] | input_a[2];
  assign popcount35_1ht9_core_069 = input_a[5] & input_a[19];
  assign popcount35_1ht9_core_070 = input_a[1] ^ input_a[8];
  assign popcount35_1ht9_core_071 = ~(input_a[27] ^ input_a[8]);
  assign popcount35_1ht9_core_072 = ~input_a[13];
  assign popcount35_1ht9_core_073 = ~(input_a[23] & input_a[33]);
  assign popcount35_1ht9_core_074 = input_a[1] ^ input_a[32];
  assign popcount35_1ht9_core_075 = input_a[24] ^ input_a[11];
  assign popcount35_1ht9_core_076 = input_a[20] & input_a[15];
  assign popcount35_1ht9_core_077 = input_a[31] ^ input_a[32];
  assign popcount35_1ht9_core_081 = input_a[22] ^ input_a[8];
  assign popcount35_1ht9_core_082 = ~(input_a[18] ^ input_a[19]);
  assign popcount35_1ht9_core_084 = input_a[33] | input_a[11];
  assign popcount35_1ht9_core_085 = input_a[9] | input_a[1];
  assign popcount35_1ht9_core_086 = input_a[20] & input_a[6];
  assign popcount35_1ht9_core_089 = input_a[4] & input_a[33];
  assign popcount35_1ht9_core_090 = input_a[0] ^ input_a[13];
  assign popcount35_1ht9_core_091 = ~(input_a[16] ^ input_a[1]);
  assign popcount35_1ht9_core_092 = input_a[2] | input_a[3];
  assign popcount35_1ht9_core_094 = ~(input_a[19] & input_a[31]);
  assign popcount35_1ht9_core_097 = ~(input_a[22] | input_a[9]);
  assign popcount35_1ht9_core_099 = ~input_a[21];
  assign popcount35_1ht9_core_100 = ~(input_a[7] ^ input_a[5]);
  assign popcount35_1ht9_core_101 = ~input_a[9];
  assign popcount35_1ht9_core_102 = input_a[8] ^ input_a[15];
  assign popcount35_1ht9_core_103 = ~(input_a[4] | input_a[18]);
  assign popcount35_1ht9_core_106 = ~input_a[17];
  assign popcount35_1ht9_core_107 = input_a[30] ^ input_a[33];
  assign popcount35_1ht9_core_108 = input_a[11] | input_a[6];
  assign popcount35_1ht9_core_110 = ~(input_a[13] ^ input_a[29]);
  assign popcount35_1ht9_core_112 = input_a[27] & input_a[29];
  assign popcount35_1ht9_core_113 = input_a[31] ^ input_a[29];
  assign popcount35_1ht9_core_114 = input_a[29] & input_a[5];
  assign popcount35_1ht9_core_115 = ~(input_a[32] & input_a[4]);
  assign popcount35_1ht9_core_117 = ~(input_a[16] | input_a[27]);
  assign popcount35_1ht9_core_118 = ~(input_a[23] & input_a[33]);
  assign popcount35_1ht9_core_119 = ~(input_a[13] & input_a[0]);
  assign popcount35_1ht9_core_120 = input_a[8] | input_a[23];
  assign popcount35_1ht9_core_123 = ~(input_a[23] ^ input_a[4]);
  assign popcount35_1ht9_core_124 = input_a[17] | input_a[33];
  assign popcount35_1ht9_core_125 = ~(input_a[6] & input_a[15]);
  assign popcount35_1ht9_core_126 = ~(input_a[21] ^ input_a[22]);
  assign popcount35_1ht9_core_127 = ~input_a[10];
  assign popcount35_1ht9_core_128 = ~(input_a[18] ^ input_a[19]);
  assign popcount35_1ht9_core_130 = input_a[21] | input_a[17];
  assign popcount35_1ht9_core_131 = ~(input_a[28] & input_a[1]);
  assign popcount35_1ht9_core_133 = input_a[9] | input_a[32];
  assign popcount35_1ht9_core_134 = input_a[6] ^ input_a[25];
  assign popcount35_1ht9_core_135 = ~(input_a[0] ^ input_a[32]);
  assign popcount35_1ht9_core_136 = ~(input_a[29] ^ input_a[9]);
  assign popcount35_1ht9_core_137 = input_a[11] ^ input_a[25];
  assign popcount35_1ht9_core_138 = ~(input_a[18] ^ input_a[9]);
  assign popcount35_1ht9_core_140 = input_a[10] ^ input_a[22];
  assign popcount35_1ht9_core_141 = ~(input_a[26] & input_a[32]);
  assign popcount35_1ht9_core_142 = ~(input_a[26] ^ input_a[24]);
  assign popcount35_1ht9_core_146 = input_a[12] ^ input_a[29];
  assign popcount35_1ht9_core_147 = ~(input_a[33] ^ input_a[10]);
  assign popcount35_1ht9_core_148 = ~(input_a[23] ^ input_a[4]);
  assign popcount35_1ht9_core_150 = ~(input_a[32] | input_a[23]);
  assign popcount35_1ht9_core_151 = ~(input_a[26] ^ input_a[22]);
  assign popcount35_1ht9_core_152 = input_a[2] & input_a[9];
  assign popcount35_1ht9_core_153 = ~(input_a[34] & input_a[34]);
  assign popcount35_1ht9_core_154 = input_a[5] ^ input_a[18];
  assign popcount35_1ht9_core_157 = ~input_a[13];
  assign popcount35_1ht9_core_158 = ~(input_a[25] ^ input_a[4]);
  assign popcount35_1ht9_core_159 = ~(input_a[26] & input_a[2]);
  assign popcount35_1ht9_core_162 = ~(input_a[22] & input_a[31]);
  assign popcount35_1ht9_core_165 = ~input_a[12];
  assign popcount35_1ht9_core_166 = input_a[31] ^ input_a[21];
  assign popcount35_1ht9_core_167 = ~input_a[13];
  assign popcount35_1ht9_core_169 = ~(input_a[34] | input_a[6]);
  assign popcount35_1ht9_core_170 = input_a[9] & input_a[31];
  assign popcount35_1ht9_core_172 = input_a[6] ^ input_a[23];
  assign popcount35_1ht9_core_173 = ~input_a[2];
  assign popcount35_1ht9_core_175 = ~input_a[24];
  assign popcount35_1ht9_core_176 = ~(input_a[13] | input_a[8]);
  assign popcount35_1ht9_core_178 = ~input_a[11];
  assign popcount35_1ht9_core_179_not = ~input_a[21];
  assign popcount35_1ht9_core_180 = input_a[18] & input_a[11];
  assign popcount35_1ht9_core_181 = input_a[21] ^ input_a[4];
  assign popcount35_1ht9_core_183 = ~(input_a[32] & input_a[30]);
  assign popcount35_1ht9_core_186 = ~(input_a[24] ^ input_a[27]);
  assign popcount35_1ht9_core_187 = ~(input_a[10] ^ input_a[26]);
  assign popcount35_1ht9_core_190 = ~input_a[4];
  assign popcount35_1ht9_core_191 = ~(input_a[14] | input_a[34]);
  assign popcount35_1ht9_core_192 = ~(input_a[30] & input_a[21]);
  assign popcount35_1ht9_core_197 = input_a[1] | input_a[2];
  assign popcount35_1ht9_core_200 = ~(input_a[10] ^ input_a[6]);
  assign popcount35_1ht9_core_201 = ~(input_a[0] & input_a[27]);
  assign popcount35_1ht9_core_202 = input_a[4] ^ input_a[33];
  assign popcount35_1ht9_core_203 = input_a[14] & input_a[11];
  assign popcount35_1ht9_core_204 = ~(input_a[12] | input_a[23]);
  assign popcount35_1ht9_core_207 = ~(input_a[25] & input_a[27]);
  assign popcount35_1ht9_core_208 = ~(input_a[26] & input_a[20]);
  assign popcount35_1ht9_core_209 = input_a[28] | input_a[13];
  assign popcount35_1ht9_core_212 = ~(input_a[19] & input_a[4]);
  assign popcount35_1ht9_core_215 = ~(input_a[27] & input_a[7]);
  assign popcount35_1ht9_core_216 = input_a[27] ^ input_a[6];
  assign popcount35_1ht9_core_219 = input_a[31] ^ input_a[26];
  assign popcount35_1ht9_core_220 = input_a[18] ^ input_a[0];
  assign popcount35_1ht9_core_223 = input_a[13] | input_a[0];
  assign popcount35_1ht9_core_224 = input_a[21] | input_a[32];
  assign popcount35_1ht9_core_225 = input_a[33] | input_a[12];
  assign popcount35_1ht9_core_226 = ~(input_a[7] | input_a[5]);
  assign popcount35_1ht9_core_227 = ~input_a[17];
  assign popcount35_1ht9_core_231 = ~(input_a[4] ^ input_a[34]);
  assign popcount35_1ht9_core_233 = input_a[10] & input_a[13];
  assign popcount35_1ht9_core_235 = ~(input_a[10] | input_a[15]);
  assign popcount35_1ht9_core_236 = input_a[0] & input_a[5];
  assign popcount35_1ht9_core_237 = input_a[3] ^ input_a[6];
  assign popcount35_1ht9_core_238 = ~(input_a[4] ^ input_a[9]);
  assign popcount35_1ht9_core_239 = ~(input_a[21] & input_a[1]);
  assign popcount35_1ht9_core_240 = ~(input_a[2] ^ input_a[13]);
  assign popcount35_1ht9_core_242 = input_a[5] & input_a[5];
  assign popcount35_1ht9_core_243 = input_a[18] ^ input_a[21];
  assign popcount35_1ht9_core_244 = ~(input_a[10] ^ input_a[22]);
  assign popcount35_1ht9_core_246 = input_a[3] ^ input_a[28];
  assign popcount35_1ht9_core_249 = ~(input_a[6] ^ input_a[13]);
  assign popcount35_1ht9_core_250 = ~input_a[1];
  assign popcount35_1ht9_core_251 = ~(input_a[19] ^ input_a[9]);
  assign popcount35_1ht9_core_252 = input_a[24] | input_a[4];
  assign popcount35_1ht9_core_253 = input_a[22] & input_a[3];
  assign popcount35_1ht9_core_254 = ~(input_a[0] & input_a[23]);
  assign popcount35_1ht9_core_257 = ~(input_a[11] & input_a[23]);
  assign popcount35_1ht9_core_258 = ~input_a[25];
  assign popcount35_1ht9_core_259 = input_a[31] & input_a[20];
  assign popcount35_1ht9_core_260 = ~(input_a[10] ^ input_a[7]);
  assign popcount35_1ht9_core_264 = input_a[32] ^ input_a[31];

  assign popcount35_1ht9_out[0] = 1'b1;
  assign popcount35_1ht9_out[1] = input_a[28];
  assign popcount35_1ht9_out[2] = input_a[27];
  assign popcount35_1ht9_out[3] = input_a[9];
  assign popcount35_1ht9_out[4] = 1'b1;
  assign popcount35_1ht9_out[5] = 1'b0;
endmodule