// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.1759
// WCE=17.0
// EP=0.914479%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_95lk(input [21:0] input_a, output [4:0] popcount22_95lk_out);
  wire popcount22_95lk_core_025;
  wire popcount22_95lk_core_026;
  wire popcount22_95lk_core_027;
  wire popcount22_95lk_core_028;
  wire popcount22_95lk_core_029;
  wire popcount22_95lk_core_031;
  wire popcount22_95lk_core_032;
  wire popcount22_95lk_core_034;
  wire popcount22_95lk_core_035;
  wire popcount22_95lk_core_037;
  wire popcount22_95lk_core_040;
  wire popcount22_95lk_core_041;
  wire popcount22_95lk_core_043;
  wire popcount22_95lk_core_045;
  wire popcount22_95lk_core_046;
  wire popcount22_95lk_core_047;
  wire popcount22_95lk_core_049;
  wire popcount22_95lk_core_052;
  wire popcount22_95lk_core_053;
  wire popcount22_95lk_core_054;
  wire popcount22_95lk_core_057;
  wire popcount22_95lk_core_058;
  wire popcount22_95lk_core_062;
  wire popcount22_95lk_core_066_not;
  wire popcount22_95lk_core_067;
  wire popcount22_95lk_core_068;
  wire popcount22_95lk_core_070;
  wire popcount22_95lk_core_072;
  wire popcount22_95lk_core_075;
  wire popcount22_95lk_core_076;
  wire popcount22_95lk_core_077;
  wire popcount22_95lk_core_080;
  wire popcount22_95lk_core_081;
  wire popcount22_95lk_core_086;
  wire popcount22_95lk_core_089;
  wire popcount22_95lk_core_090;
  wire popcount22_95lk_core_091;
  wire popcount22_95lk_core_092;
  wire popcount22_95lk_core_093;
  wire popcount22_95lk_core_097;
  wire popcount22_95lk_core_098;
  wire popcount22_95lk_core_099;
  wire popcount22_95lk_core_100;
  wire popcount22_95lk_core_101;
  wire popcount22_95lk_core_103;
  wire popcount22_95lk_core_105;
  wire popcount22_95lk_core_107;
  wire popcount22_95lk_core_110;
  wire popcount22_95lk_core_113_not;
  wire popcount22_95lk_core_114;
  wire popcount22_95lk_core_116;
  wire popcount22_95lk_core_119;
  wire popcount22_95lk_core_121;
  wire popcount22_95lk_core_122;
  wire popcount22_95lk_core_123;
  wire popcount22_95lk_core_124;
  wire popcount22_95lk_core_125;
  wire popcount22_95lk_core_126;
  wire popcount22_95lk_core_129;
  wire popcount22_95lk_core_130;
  wire popcount22_95lk_core_132;
  wire popcount22_95lk_core_136;
  wire popcount22_95lk_core_138;
  wire popcount22_95lk_core_139;
  wire popcount22_95lk_core_143;
  wire popcount22_95lk_core_144_not;
  wire popcount22_95lk_core_145;
  wire popcount22_95lk_core_146;
  wire popcount22_95lk_core_147;
  wire popcount22_95lk_core_149;
  wire popcount22_95lk_core_151;
  wire popcount22_95lk_core_153;
  wire popcount22_95lk_core_155;
  wire popcount22_95lk_core_156;
  wire popcount22_95lk_core_157;
  wire popcount22_95lk_core_161;

  assign popcount22_95lk_core_025 = ~(input_a[20] & input_a[5]);
  assign popcount22_95lk_core_026 = input_a[6] | input_a[12];
  assign popcount22_95lk_core_027 = ~(input_a[18] | input_a[10]);
  assign popcount22_95lk_core_028 = ~(input_a[2] | input_a[21]);
  assign popcount22_95lk_core_029 = input_a[2] | input_a[2];
  assign popcount22_95lk_core_031 = ~(input_a[21] & input_a[17]);
  assign popcount22_95lk_core_032 = ~(input_a[13] | input_a[19]);
  assign popcount22_95lk_core_034 = input_a[19] ^ input_a[12];
  assign popcount22_95lk_core_035 = ~(input_a[0] & input_a[20]);
  assign popcount22_95lk_core_037 = input_a[8] ^ input_a[15];
  assign popcount22_95lk_core_040 = ~(input_a[14] & input_a[7]);
  assign popcount22_95lk_core_041 = input_a[16] | input_a[14];
  assign popcount22_95lk_core_043 = ~(input_a[0] | input_a[6]);
  assign popcount22_95lk_core_045 = input_a[1] ^ input_a[3];
  assign popcount22_95lk_core_046 = ~input_a[16];
  assign popcount22_95lk_core_047 = ~(input_a[14] | input_a[19]);
  assign popcount22_95lk_core_049 = ~input_a[19];
  assign popcount22_95lk_core_052 = input_a[13] ^ input_a[17];
  assign popcount22_95lk_core_053 = input_a[9] | input_a[21];
  assign popcount22_95lk_core_054 = ~(input_a[12] & input_a[6]);
  assign popcount22_95lk_core_057 = ~(input_a[10] & input_a[9]);
  assign popcount22_95lk_core_058 = input_a[0] | input_a[2];
  assign popcount22_95lk_core_062 = ~input_a[2];
  assign popcount22_95lk_core_066_not = ~input_a[1];
  assign popcount22_95lk_core_067 = input_a[8] | input_a[12];
  assign popcount22_95lk_core_068 = ~(input_a[10] | input_a[12]);
  assign popcount22_95lk_core_070 = input_a[8] ^ input_a[4];
  assign popcount22_95lk_core_072 = input_a[8] & input_a[0];
  assign popcount22_95lk_core_075 = input_a[13] & input_a[4];
  assign popcount22_95lk_core_076 = input_a[21] ^ input_a[1];
  assign popcount22_95lk_core_077 = input_a[10] | input_a[0];
  assign popcount22_95lk_core_080 = input_a[18] | input_a[14];
  assign popcount22_95lk_core_081 = ~(input_a[5] & input_a[21]);
  assign popcount22_95lk_core_086 = input_a[15] ^ input_a[12];
  assign popcount22_95lk_core_089 = input_a[4] | input_a[7];
  assign popcount22_95lk_core_090 = ~input_a[0];
  assign popcount22_95lk_core_091 = input_a[3] ^ input_a[1];
  assign popcount22_95lk_core_092 = ~(input_a[21] ^ input_a[9]);
  assign popcount22_95lk_core_093 = ~(input_a[7] ^ input_a[6]);
  assign popcount22_95lk_core_097 = input_a[16] | input_a[13];
  assign popcount22_95lk_core_098 = input_a[19] ^ input_a[16];
  assign popcount22_95lk_core_099 = ~(input_a[5] & input_a[21]);
  assign popcount22_95lk_core_100 = ~(input_a[7] ^ input_a[8]);
  assign popcount22_95lk_core_101 = input_a[3] & input_a[13];
  assign popcount22_95lk_core_103 = input_a[20] ^ input_a[6];
  assign popcount22_95lk_core_105 = ~(input_a[9] | input_a[8]);
  assign popcount22_95lk_core_107 = ~(input_a[6] | input_a[13]);
  assign popcount22_95lk_core_110 = ~(input_a[8] | input_a[21]);
  assign popcount22_95lk_core_113_not = ~input_a[14];
  assign popcount22_95lk_core_114 = input_a[0] | input_a[0];
  assign popcount22_95lk_core_116 = input_a[20] | input_a[7];
  assign popcount22_95lk_core_119 = ~(input_a[6] ^ input_a[6]);
  assign popcount22_95lk_core_121 = ~input_a[17];
  assign popcount22_95lk_core_122 = ~input_a[11];
  assign popcount22_95lk_core_123 = input_a[10] ^ input_a[15];
  assign popcount22_95lk_core_124 = ~input_a[21];
  assign popcount22_95lk_core_125 = ~(input_a[9] | input_a[20]);
  assign popcount22_95lk_core_126 = ~(input_a[5] ^ input_a[9]);
  assign popcount22_95lk_core_129 = ~(input_a[8] ^ input_a[3]);
  assign popcount22_95lk_core_130 = ~input_a[10];
  assign popcount22_95lk_core_132 = input_a[3] & input_a[10];
  assign popcount22_95lk_core_136 = input_a[16] ^ input_a[10];
  assign popcount22_95lk_core_138 = ~(input_a[2] ^ input_a[11]);
  assign popcount22_95lk_core_139 = input_a[15] ^ input_a[13];
  assign popcount22_95lk_core_143 = input_a[7] | input_a[16];
  assign popcount22_95lk_core_144_not = ~input_a[12];
  assign popcount22_95lk_core_145 = input_a[5] | input_a[5];
  assign popcount22_95lk_core_146 = ~(input_a[5] | input_a[17]);
  assign popcount22_95lk_core_147 = input_a[20] ^ input_a[11];
  assign popcount22_95lk_core_149 = input_a[4] & input_a[9];
  assign popcount22_95lk_core_151 = ~(input_a[3] | input_a[20]);
  assign popcount22_95lk_core_153 = ~(input_a[13] ^ input_a[2]);
  assign popcount22_95lk_core_155 = ~(input_a[12] & input_a[15]);
  assign popcount22_95lk_core_156 = input_a[4] | input_a[17];
  assign popcount22_95lk_core_157 = ~(input_a[18] | input_a[12]);
  assign popcount22_95lk_core_161 = ~(input_a[8] ^ input_a[21]);

  assign popcount22_95lk_out[0] = 1'b0;
  assign popcount22_95lk_out[1] = 1'b0;
  assign popcount22_95lk_out[2] = 1'b1;
  assign popcount22_95lk_out[3] = input_a[2];
  assign popcount22_95lk_out[4] = 1'b0;
endmodule