// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.16352
// WCE=18.0
// EP=0.948785%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_zzpw(input [26:0] input_a, output [4:0] popcount27_zzpw_out);
  wire popcount27_zzpw_core_029;
  wire popcount27_zzpw_core_030;
  wire popcount27_zzpw_core_032;
  wire popcount27_zzpw_core_033;
  wire popcount27_zzpw_core_036;
  wire popcount27_zzpw_core_037;
  wire popcount27_zzpw_core_038;
  wire popcount27_zzpw_core_040;
  wire popcount27_zzpw_core_042;
  wire popcount27_zzpw_core_043;
  wire popcount27_zzpw_core_044;
  wire popcount27_zzpw_core_046;
  wire popcount27_zzpw_core_049;
  wire popcount27_zzpw_core_050;
  wire popcount27_zzpw_core_051;
  wire popcount27_zzpw_core_052;
  wire popcount27_zzpw_core_055;
  wire popcount27_zzpw_core_056;
  wire popcount27_zzpw_core_058;
  wire popcount27_zzpw_core_061;
  wire popcount27_zzpw_core_062;
  wire popcount27_zzpw_core_064;
  wire popcount27_zzpw_core_066;
  wire popcount27_zzpw_core_067;
  wire popcount27_zzpw_core_068;
  wire popcount27_zzpw_core_069;
  wire popcount27_zzpw_core_070;
  wire popcount27_zzpw_core_073;
  wire popcount27_zzpw_core_074;
  wire popcount27_zzpw_core_075;
  wire popcount27_zzpw_core_076;
  wire popcount27_zzpw_core_077;
  wire popcount27_zzpw_core_078;
  wire popcount27_zzpw_core_081;
  wire popcount27_zzpw_core_082;
  wire popcount27_zzpw_core_086;
  wire popcount27_zzpw_core_088;
  wire popcount27_zzpw_core_089_not;
  wire popcount27_zzpw_core_090;
  wire popcount27_zzpw_core_091;
  wire popcount27_zzpw_core_093;
  wire popcount27_zzpw_core_094;
  wire popcount27_zzpw_core_095_not;
  wire popcount27_zzpw_core_096;
  wire popcount27_zzpw_core_098;
  wire popcount27_zzpw_core_099;
  wire popcount27_zzpw_core_100;
  wire popcount27_zzpw_core_101;
  wire popcount27_zzpw_core_104;
  wire popcount27_zzpw_core_106;
  wire popcount27_zzpw_core_107;
  wire popcount27_zzpw_core_108;
  wire popcount27_zzpw_core_109;
  wire popcount27_zzpw_core_110;
  wire popcount27_zzpw_core_114;
  wire popcount27_zzpw_core_116;
  wire popcount27_zzpw_core_117;
  wire popcount27_zzpw_core_119;
  wire popcount27_zzpw_core_120;
  wire popcount27_zzpw_core_122;
  wire popcount27_zzpw_core_123;
  wire popcount27_zzpw_core_124;
  wire popcount27_zzpw_core_126;
  wire popcount27_zzpw_core_127;
  wire popcount27_zzpw_core_128;
  wire popcount27_zzpw_core_129;
  wire popcount27_zzpw_core_130_not;
  wire popcount27_zzpw_core_131;
  wire popcount27_zzpw_core_134;
  wire popcount27_zzpw_core_135;
  wire popcount27_zzpw_core_140;
  wire popcount27_zzpw_core_141;
  wire popcount27_zzpw_core_144;
  wire popcount27_zzpw_core_146;
  wire popcount27_zzpw_core_147;
  wire popcount27_zzpw_core_148;
  wire popcount27_zzpw_core_149;
  wire popcount27_zzpw_core_151_not;
  wire popcount27_zzpw_core_152;
  wire popcount27_zzpw_core_154;
  wire popcount27_zzpw_core_156;
  wire popcount27_zzpw_core_157;
  wire popcount27_zzpw_core_158;
  wire popcount27_zzpw_core_159;
  wire popcount27_zzpw_core_160;
  wire popcount27_zzpw_core_161;
  wire popcount27_zzpw_core_162;
  wire popcount27_zzpw_core_165;
  wire popcount27_zzpw_core_166;
  wire popcount27_zzpw_core_167;
  wire popcount27_zzpw_core_169;
  wire popcount27_zzpw_core_173;
  wire popcount27_zzpw_core_174;
  wire popcount27_zzpw_core_176;
  wire popcount27_zzpw_core_177;
  wire popcount27_zzpw_core_178;
  wire popcount27_zzpw_core_180;
  wire popcount27_zzpw_core_181;
  wire popcount27_zzpw_core_182;
  wire popcount27_zzpw_core_183;
  wire popcount27_zzpw_core_184;
  wire popcount27_zzpw_core_185;
  wire popcount27_zzpw_core_187;
  wire popcount27_zzpw_core_190_not;
  wire popcount27_zzpw_core_191;
  wire popcount27_zzpw_core_192;
  wire popcount27_zzpw_core_193;
  wire popcount27_zzpw_core_194;
  wire popcount27_zzpw_core_195;

  assign popcount27_zzpw_core_029 = ~(input_a[17] | input_a[8]);
  assign popcount27_zzpw_core_030 = ~input_a[26];
  assign popcount27_zzpw_core_032 = input_a[21] | input_a[25];
  assign popcount27_zzpw_core_033 = ~(input_a[22] ^ input_a[6]);
  assign popcount27_zzpw_core_036 = ~(input_a[10] ^ input_a[23]);
  assign popcount27_zzpw_core_037 = input_a[6] ^ input_a[4];
  assign popcount27_zzpw_core_038 = input_a[8] & input_a[11];
  assign popcount27_zzpw_core_040 = ~(input_a[0] ^ input_a[16]);
  assign popcount27_zzpw_core_042 = ~input_a[4];
  assign popcount27_zzpw_core_043 = input_a[23] & input_a[4];
  assign popcount27_zzpw_core_044 = ~(input_a[20] & input_a[25]);
  assign popcount27_zzpw_core_046 = input_a[6] | input_a[1];
  assign popcount27_zzpw_core_049 = ~(input_a[18] | input_a[2]);
  assign popcount27_zzpw_core_050 = input_a[9] ^ input_a[18];
  assign popcount27_zzpw_core_051 = ~input_a[22];
  assign popcount27_zzpw_core_052 = ~(input_a[22] | input_a[18]);
  assign popcount27_zzpw_core_055 = input_a[18] & input_a[18];
  assign popcount27_zzpw_core_056 = input_a[19] | input_a[22];
  assign popcount27_zzpw_core_058 = input_a[20] | input_a[26];
  assign popcount27_zzpw_core_061 = ~(input_a[7] ^ input_a[3]);
  assign popcount27_zzpw_core_062 = ~input_a[18];
  assign popcount27_zzpw_core_064 = input_a[1] | input_a[4];
  assign popcount27_zzpw_core_066 = ~(input_a[7] ^ input_a[0]);
  assign popcount27_zzpw_core_067 = ~input_a[17];
  assign popcount27_zzpw_core_068 = ~(input_a[9] | input_a[24]);
  assign popcount27_zzpw_core_069 = input_a[13] ^ input_a[6];
  assign popcount27_zzpw_core_070 = ~(input_a[6] & input_a[6]);
  assign popcount27_zzpw_core_073 = ~(input_a[17] & input_a[5]);
  assign popcount27_zzpw_core_074 = ~(input_a[21] ^ input_a[4]);
  assign popcount27_zzpw_core_075 = input_a[20] ^ input_a[15];
  assign popcount27_zzpw_core_076 = ~(input_a[5] ^ input_a[16]);
  assign popcount27_zzpw_core_077 = ~(input_a[10] | input_a[3]);
  assign popcount27_zzpw_core_078 = ~(input_a[0] & input_a[11]);
  assign popcount27_zzpw_core_081 = ~(input_a[25] ^ input_a[17]);
  assign popcount27_zzpw_core_082 = ~(input_a[20] ^ input_a[26]);
  assign popcount27_zzpw_core_086 = input_a[25] & input_a[25];
  assign popcount27_zzpw_core_088 = input_a[17] & input_a[24];
  assign popcount27_zzpw_core_089_not = ~input_a[12];
  assign popcount27_zzpw_core_090 = ~(input_a[24] ^ input_a[5]);
  assign popcount27_zzpw_core_091 = ~(input_a[26] ^ input_a[6]);
  assign popcount27_zzpw_core_093 = ~(input_a[17] & input_a[23]);
  assign popcount27_zzpw_core_094 = input_a[25] ^ input_a[14];
  assign popcount27_zzpw_core_095_not = ~input_a[18];
  assign popcount27_zzpw_core_096 = input_a[16] & input_a[3];
  assign popcount27_zzpw_core_098 = input_a[1] ^ input_a[24];
  assign popcount27_zzpw_core_099 = ~input_a[13];
  assign popcount27_zzpw_core_100 = ~(input_a[1] & input_a[14]);
  assign popcount27_zzpw_core_101 = ~input_a[15];
  assign popcount27_zzpw_core_104 = ~input_a[15];
  assign popcount27_zzpw_core_106 = ~(input_a[3] ^ input_a[17]);
  assign popcount27_zzpw_core_107 = ~(input_a[3] ^ input_a[12]);
  assign popcount27_zzpw_core_108 = input_a[0] & input_a[17];
  assign popcount27_zzpw_core_109 = input_a[13] ^ input_a[18];
  assign popcount27_zzpw_core_110 = ~(input_a[8] | input_a[16]);
  assign popcount27_zzpw_core_114 = ~(input_a[13] ^ input_a[18]);
  assign popcount27_zzpw_core_116 = ~(input_a[14] & input_a[17]);
  assign popcount27_zzpw_core_117 = ~(input_a[21] & input_a[12]);
  assign popcount27_zzpw_core_119 = ~(input_a[23] & input_a[16]);
  assign popcount27_zzpw_core_120 = ~input_a[10];
  assign popcount27_zzpw_core_122 = ~(input_a[20] | input_a[22]);
  assign popcount27_zzpw_core_123 = ~(input_a[25] | input_a[5]);
  assign popcount27_zzpw_core_124 = ~(input_a[24] ^ input_a[10]);
  assign popcount27_zzpw_core_126 = ~(input_a[15] & input_a[11]);
  assign popcount27_zzpw_core_127 = ~(input_a[1] | input_a[6]);
  assign popcount27_zzpw_core_128 = ~input_a[2];
  assign popcount27_zzpw_core_129 = ~input_a[25];
  assign popcount27_zzpw_core_130_not = ~input_a[10];
  assign popcount27_zzpw_core_131 = input_a[10] & input_a[4];
  assign popcount27_zzpw_core_134 = ~(input_a[22] ^ input_a[7]);
  assign popcount27_zzpw_core_135 = ~(input_a[6] & input_a[2]);
  assign popcount27_zzpw_core_140 = ~(input_a[10] & input_a[25]);
  assign popcount27_zzpw_core_141 = input_a[23] | input_a[24];
  assign popcount27_zzpw_core_144 = input_a[0] & input_a[5];
  assign popcount27_zzpw_core_146 = ~input_a[13];
  assign popcount27_zzpw_core_147 = ~(input_a[24] | input_a[5]);
  assign popcount27_zzpw_core_148 = ~input_a[15];
  assign popcount27_zzpw_core_149 = input_a[8] | input_a[8];
  assign popcount27_zzpw_core_151_not = ~input_a[18];
  assign popcount27_zzpw_core_152 = input_a[2] & input_a[20];
  assign popcount27_zzpw_core_154 = ~(input_a[1] | input_a[2]);
  assign popcount27_zzpw_core_156 = input_a[3] | input_a[26];
  assign popcount27_zzpw_core_157 = input_a[23] & input_a[13];
  assign popcount27_zzpw_core_158 = input_a[15] ^ input_a[4];
  assign popcount27_zzpw_core_159 = ~(input_a[0] ^ input_a[2]);
  assign popcount27_zzpw_core_160 = input_a[21] ^ input_a[18];
  assign popcount27_zzpw_core_161 = input_a[23] | input_a[1];
  assign popcount27_zzpw_core_162 = input_a[22] & input_a[7];
  assign popcount27_zzpw_core_165 = input_a[16] | input_a[9];
  assign popcount27_zzpw_core_166 = ~(input_a[26] | input_a[4]);
  assign popcount27_zzpw_core_167 = input_a[5] ^ input_a[24];
  assign popcount27_zzpw_core_169 = ~(input_a[8] & input_a[24]);
  assign popcount27_zzpw_core_173 = input_a[12] ^ input_a[5];
  assign popcount27_zzpw_core_174 = ~(input_a[9] | input_a[17]);
  assign popcount27_zzpw_core_176 = ~input_a[24];
  assign popcount27_zzpw_core_177 = ~(input_a[1] ^ input_a[23]);
  assign popcount27_zzpw_core_178 = input_a[25] ^ input_a[6];
  assign popcount27_zzpw_core_180 = ~(input_a[0] ^ input_a[11]);
  assign popcount27_zzpw_core_181 = ~input_a[19];
  assign popcount27_zzpw_core_182 = ~input_a[25];
  assign popcount27_zzpw_core_183 = ~(input_a[25] & input_a[26]);
  assign popcount27_zzpw_core_184 = ~(input_a[5] | input_a[24]);
  assign popcount27_zzpw_core_185 = input_a[8] ^ input_a[23];
  assign popcount27_zzpw_core_187 = input_a[10] & input_a[22];
  assign popcount27_zzpw_core_190_not = ~input_a[22];
  assign popcount27_zzpw_core_191 = ~(input_a[10] | input_a[13]);
  assign popcount27_zzpw_core_192 = input_a[5] | input_a[8];
  assign popcount27_zzpw_core_193 = ~(input_a[11] | input_a[12]);
  assign popcount27_zzpw_core_194 = ~(input_a[8] | input_a[3]);
  assign popcount27_zzpw_core_195 = input_a[8] & input_a[16];

  assign popcount27_zzpw_out[0] = input_a[15];
  assign popcount27_zzpw_out[1] = 1'b1;
  assign popcount27_zzpw_out[2] = 1'b0;
  assign popcount27_zzpw_out[3] = 1'b1;
  assign popcount27_zzpw_out[4] = 1'b0;
endmodule