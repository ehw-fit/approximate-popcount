// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.99787
// WCE=20.0
// EP=0.843477%
// Printed PDK parameters:
//  Area=59274083.0
//  Delay=70444192.0
//  Power=3113900.0

module popcount40_jl9s(input [39:0] input_a, output [5:0] popcount40_jl9s_out);
  wire popcount40_jl9s_core_045;
  wire popcount40_jl9s_core_047;
  wire popcount40_jl9s_core_049_not;
  wire popcount40_jl9s_core_050;
  wire popcount40_jl9s_core_051;
  wire popcount40_jl9s_core_053;
  wire popcount40_jl9s_core_054;
  wire popcount40_jl9s_core_058;
  wire popcount40_jl9s_core_059;
  wire popcount40_jl9s_core_060;
  wire popcount40_jl9s_core_061;
  wire popcount40_jl9s_core_062;
  wire popcount40_jl9s_core_067;
  wire popcount40_jl9s_core_068;
  wire popcount40_jl9s_core_070;
  wire popcount40_jl9s_core_073_not;
  wire popcount40_jl9s_core_074;
  wire popcount40_jl9s_core_077;
  wire popcount40_jl9s_core_078;
  wire popcount40_jl9s_core_079;
  wire popcount40_jl9s_core_081;
  wire popcount40_jl9s_core_082;
  wire popcount40_jl9s_core_084;
  wire popcount40_jl9s_core_087;
  wire popcount40_jl9s_core_091;
  wire popcount40_jl9s_core_092;
  wire popcount40_jl9s_core_093;
  wire popcount40_jl9s_core_094;
  wire popcount40_jl9s_core_096;
  wire popcount40_jl9s_core_098;
  wire popcount40_jl9s_core_099_not;
  wire popcount40_jl9s_core_102;
  wire popcount40_jl9s_core_103;
  wire popcount40_jl9s_core_106;
  wire popcount40_jl9s_core_109_not;
  wire popcount40_jl9s_core_111;
  wire popcount40_jl9s_core_113;
  wire popcount40_jl9s_core_114;
  wire popcount40_jl9s_core_116;
  wire popcount40_jl9s_core_119;
  wire popcount40_jl9s_core_120;
  wire popcount40_jl9s_core_121;
  wire popcount40_jl9s_core_126;
  wire popcount40_jl9s_core_127;
  wire popcount40_jl9s_core_128;
  wire popcount40_jl9s_core_129;
  wire popcount40_jl9s_core_130;
  wire popcount40_jl9s_core_131;
  wire popcount40_jl9s_core_132;
  wire popcount40_jl9s_core_133;
  wire popcount40_jl9s_core_134;
  wire popcount40_jl9s_core_135;
  wire popcount40_jl9s_core_136;
  wire popcount40_jl9s_core_137;
  wire popcount40_jl9s_core_138;
  wire popcount40_jl9s_core_140;
  wire popcount40_jl9s_core_144;
  wire popcount40_jl9s_core_145;
  wire popcount40_jl9s_core_146_not;
  wire popcount40_jl9s_core_148;
  wire popcount40_jl9s_core_149;
  wire popcount40_jl9s_core_150;
  wire popcount40_jl9s_core_153;
  wire popcount40_jl9s_core_154;
  wire popcount40_jl9s_core_158;
  wire popcount40_jl9s_core_159;
  wire popcount40_jl9s_core_160;
  wire popcount40_jl9s_core_162;
  wire popcount40_jl9s_core_164;
  wire popcount40_jl9s_core_166;
  wire popcount40_jl9s_core_167;
  wire popcount40_jl9s_core_168;
  wire popcount40_jl9s_core_170;
  wire popcount40_jl9s_core_172;
  wire popcount40_jl9s_core_173;
  wire popcount40_jl9s_core_174;
  wire popcount40_jl9s_core_175;
  wire popcount40_jl9s_core_176;
  wire popcount40_jl9s_core_181;
  wire popcount40_jl9s_core_183;
  wire popcount40_jl9s_core_184;
  wire popcount40_jl9s_core_186;
  wire popcount40_jl9s_core_187_not;
  wire popcount40_jl9s_core_188;
  wire popcount40_jl9s_core_191;
  wire popcount40_jl9s_core_193;
  wire popcount40_jl9s_core_194;
  wire popcount40_jl9s_core_195;
  wire popcount40_jl9s_core_196;
  wire popcount40_jl9s_core_197;
  wire popcount40_jl9s_core_199;
  wire popcount40_jl9s_core_200;
  wire popcount40_jl9s_core_201;
  wire popcount40_jl9s_core_202;
  wire popcount40_jl9s_core_203;
  wire popcount40_jl9s_core_204;
  wire popcount40_jl9s_core_205;
  wire popcount40_jl9s_core_206;
  wire popcount40_jl9s_core_207;
  wire popcount40_jl9s_core_208;
  wire popcount40_jl9s_core_209;
  wire popcount40_jl9s_core_210;
  wire popcount40_jl9s_core_211;
  wire popcount40_jl9s_core_215;
  wire popcount40_jl9s_core_216;
  wire popcount40_jl9s_core_217;
  wire popcount40_jl9s_core_218;
  wire popcount40_jl9s_core_221;
  wire popcount40_jl9s_core_222_not;
  wire popcount40_jl9s_core_223;
  wire popcount40_jl9s_core_225;
  wire popcount40_jl9s_core_227;
  wire popcount40_jl9s_core_228;
  wire popcount40_jl9s_core_229;
  wire popcount40_jl9s_core_230;
  wire popcount40_jl9s_core_231;
  wire popcount40_jl9s_core_235;
  wire popcount40_jl9s_core_236;
  wire popcount40_jl9s_core_238;
  wire popcount40_jl9s_core_239;
  wire popcount40_jl9s_core_241;
  wire popcount40_jl9s_core_245;
  wire popcount40_jl9s_core_246;
  wire popcount40_jl9s_core_247;
  wire popcount40_jl9s_core_248;
  wire popcount40_jl9s_core_250;
  wire popcount40_jl9s_core_251;
  wire popcount40_jl9s_core_253;
  wire popcount40_jl9s_core_260;
  wire popcount40_jl9s_core_261;
  wire popcount40_jl9s_core_266;
  wire popcount40_jl9s_core_267;
  wire popcount40_jl9s_core_268;
  wire popcount40_jl9s_core_269;
  wire popcount40_jl9s_core_270;
  wire popcount40_jl9s_core_271;
  wire popcount40_jl9s_core_272;
  wire popcount40_jl9s_core_273;
  wire popcount40_jl9s_core_274;
  wire popcount40_jl9s_core_275;
  wire popcount40_jl9s_core_276;
  wire popcount40_jl9s_core_277;
  wire popcount40_jl9s_core_278;
  wire popcount40_jl9s_core_279;
  wire popcount40_jl9s_core_280;
  wire popcount40_jl9s_core_281;
  wire popcount40_jl9s_core_282;
  wire popcount40_jl9s_core_283;
  wire popcount40_jl9s_core_284;
  wire popcount40_jl9s_core_286;
  wire popcount40_jl9s_core_290;
  wire popcount40_jl9s_core_291;
  wire popcount40_jl9s_core_292;
  wire popcount40_jl9s_core_293;
  wire popcount40_jl9s_core_294;
  wire popcount40_jl9s_core_295;
  wire popcount40_jl9s_core_296;
  wire popcount40_jl9s_core_297;
  wire popcount40_jl9s_core_298;
  wire popcount40_jl9s_core_299;
  wire popcount40_jl9s_core_300;
  wire popcount40_jl9s_core_301;
  wire popcount40_jl9s_core_302;
  wire popcount40_jl9s_core_303;
  wire popcount40_jl9s_core_304;
  wire popcount40_jl9s_core_305;
  wire popcount40_jl9s_core_306;
  wire popcount40_jl9s_core_308;
  wire popcount40_jl9s_core_309;
  wire popcount40_jl9s_core_310;
  wire popcount40_jl9s_core_311;
  wire popcount40_jl9s_core_313;
  wire popcount40_jl9s_core_315;
  wire popcount40_jl9s_core_316;

  assign popcount40_jl9s_core_045 = input_a[2] | input_a[31];
  assign popcount40_jl9s_core_047 = input_a[38] ^ input_a[12];
  assign popcount40_jl9s_core_049_not = ~input_a[37];
  assign popcount40_jl9s_core_050 = ~(input_a[35] | input_a[28]);
  assign popcount40_jl9s_core_051 = input_a[30] & input_a[3];
  assign popcount40_jl9s_core_053 = ~(input_a[23] ^ input_a[16]);
  assign popcount40_jl9s_core_054 = ~input_a[17];
  assign popcount40_jl9s_core_058 = input_a[6] | input_a[39];
  assign popcount40_jl9s_core_059 = input_a[38] & input_a[15];
  assign popcount40_jl9s_core_060 = input_a[2] | input_a[6];
  assign popcount40_jl9s_core_061 = input_a[3] ^ input_a[6];
  assign popcount40_jl9s_core_062 = ~(input_a[4] | input_a[17]);
  assign popcount40_jl9s_core_067 = ~(input_a[22] ^ input_a[16]);
  assign popcount40_jl9s_core_068 = input_a[17] | input_a[22];
  assign popcount40_jl9s_core_070 = input_a[21] | input_a[10];
  assign popcount40_jl9s_core_073_not = ~input_a[14];
  assign popcount40_jl9s_core_074 = input_a[29] ^ input_a[25];
  assign popcount40_jl9s_core_077 = ~input_a[12];
  assign popcount40_jl9s_core_078 = input_a[23] ^ input_a[27];
  assign popcount40_jl9s_core_079 = input_a[38] & input_a[29];
  assign popcount40_jl9s_core_081 = ~input_a[13];
  assign popcount40_jl9s_core_082 = input_a[4] ^ input_a[21];
  assign popcount40_jl9s_core_084 = ~(input_a[20] | input_a[12]);
  assign popcount40_jl9s_core_087 = input_a[7] ^ input_a[15];
  assign popcount40_jl9s_core_091 = ~input_a[7];
  assign popcount40_jl9s_core_092 = ~(input_a[31] ^ input_a[7]);
  assign popcount40_jl9s_core_093 = input_a[23] ^ input_a[32];
  assign popcount40_jl9s_core_094 = input_a[10] & input_a[38];
  assign popcount40_jl9s_core_096 = input_a[26] | input_a[15];
  assign popcount40_jl9s_core_098 = input_a[18] & input_a[31];
  assign popcount40_jl9s_core_099_not = ~input_a[39];
  assign popcount40_jl9s_core_102 = ~(input_a[39] ^ input_a[26]);
  assign popcount40_jl9s_core_103 = ~popcount40_jl9s_core_094;
  assign popcount40_jl9s_core_106 = ~(input_a[3] ^ input_a[13]);
  assign popcount40_jl9s_core_109_not = ~input_a[24];
  assign popcount40_jl9s_core_111 = input_a[12] & input_a[22];
  assign popcount40_jl9s_core_113 = input_a[35] & input_a[19];
  assign popcount40_jl9s_core_114 = ~(input_a[36] & input_a[7]);
  assign popcount40_jl9s_core_116 = popcount40_jl9s_core_113 | input_a[13];
  assign popcount40_jl9s_core_119 = ~(input_a[5] & input_a[18]);
  assign popcount40_jl9s_core_120 = popcount40_jl9s_core_111 ^ popcount40_jl9s_core_116;
  assign popcount40_jl9s_core_121 = popcount40_jl9s_core_111 & popcount40_jl9s_core_116;
  assign popcount40_jl9s_core_126 = input_a[29] & input_a[28];
  assign popcount40_jl9s_core_127 = ~(input_a[10] ^ input_a[17]);
  assign popcount40_jl9s_core_128 = input_a[36] & input_a[29];
  assign popcount40_jl9s_core_129 = popcount40_jl9s_core_103 ^ popcount40_jl9s_core_120;
  assign popcount40_jl9s_core_130 = popcount40_jl9s_core_103 & popcount40_jl9s_core_120;
  assign popcount40_jl9s_core_131 = popcount40_jl9s_core_129 ^ popcount40_jl9s_core_128;
  assign popcount40_jl9s_core_132 = popcount40_jl9s_core_129 & popcount40_jl9s_core_128;
  assign popcount40_jl9s_core_133 = popcount40_jl9s_core_130 | popcount40_jl9s_core_132;
  assign popcount40_jl9s_core_134 = popcount40_jl9s_core_094 ^ popcount40_jl9s_core_121;
  assign popcount40_jl9s_core_135 = popcount40_jl9s_core_094 & popcount40_jl9s_core_121;
  assign popcount40_jl9s_core_136 = popcount40_jl9s_core_134 ^ popcount40_jl9s_core_133;
  assign popcount40_jl9s_core_137 = popcount40_jl9s_core_134 & popcount40_jl9s_core_133;
  assign popcount40_jl9s_core_138 = popcount40_jl9s_core_135 | popcount40_jl9s_core_137;
  assign popcount40_jl9s_core_140 = ~(input_a[30] & input_a[13]);
  assign popcount40_jl9s_core_144 = input_a[12] | input_a[1];
  assign popcount40_jl9s_core_145 = input_a[32] & input_a[39];
  assign popcount40_jl9s_core_146_not = ~popcount40_jl9s_core_131;
  assign popcount40_jl9s_core_148 = popcount40_jl9s_core_146_not ^ popcount40_jl9s_core_145;
  assign popcount40_jl9s_core_149 = popcount40_jl9s_core_146_not & popcount40_jl9s_core_145;
  assign popcount40_jl9s_core_150 = popcount40_jl9s_core_131 | popcount40_jl9s_core_149;
  assign popcount40_jl9s_core_153 = popcount40_jl9s_core_136 ^ popcount40_jl9s_core_150;
  assign popcount40_jl9s_core_154 = popcount40_jl9s_core_136 & popcount40_jl9s_core_150;
  assign popcount40_jl9s_core_158 = popcount40_jl9s_core_138 ^ popcount40_jl9s_core_154;
  assign popcount40_jl9s_core_159 = ~(input_a[37] ^ input_a[5]);
  assign popcount40_jl9s_core_160 = ~input_a[23];
  assign popcount40_jl9s_core_162 = input_a[30] & input_a[5];
  assign popcount40_jl9s_core_164 = ~(input_a[27] ^ input_a[3]);
  assign popcount40_jl9s_core_166 = input_a[27] | input_a[27];
  assign popcount40_jl9s_core_167 = input_a[20] & input_a[21];
  assign popcount40_jl9s_core_168 = ~(input_a[0] ^ input_a[32]);
  assign popcount40_jl9s_core_170 = ~(input_a[27] ^ input_a[8]);
  assign popcount40_jl9s_core_172 = ~(input_a[31] & input_a[37]);
  assign popcount40_jl9s_core_173 = input_a[31] & input_a[37];
  assign popcount40_jl9s_core_174 = input_a[26] ^ input_a[5];
  assign popcount40_jl9s_core_175 = ~(input_a[14] | input_a[19]);
  assign popcount40_jl9s_core_176 = popcount40_jl9s_core_167 ^ popcount40_jl9s_core_172;
  assign popcount40_jl9s_core_181 = popcount40_jl9s_core_173 | popcount40_jl9s_core_167;
  assign popcount40_jl9s_core_183 = ~(input_a[3] & input_a[3]);
  assign popcount40_jl9s_core_184 = input_a[25] & input_a[11];
  assign popcount40_jl9s_core_186 = input_a[28] & input_a[9];
  assign popcount40_jl9s_core_187_not = ~input_a[8];
  assign popcount40_jl9s_core_188 = input_a[4] ^ input_a[21];
  assign popcount40_jl9s_core_191 = ~(popcount40_jl9s_core_183 & popcount40_jl9s_core_187_not);
  assign popcount40_jl9s_core_193 = popcount40_jl9s_core_184 ^ input_a[18];
  assign popcount40_jl9s_core_194 = popcount40_jl9s_core_184 & input_a[18];
  assign popcount40_jl9s_core_195 = popcount40_jl9s_core_193 ^ popcount40_jl9s_core_183;
  assign popcount40_jl9s_core_196 = popcount40_jl9s_core_193 & popcount40_jl9s_core_183;
  assign popcount40_jl9s_core_197 = popcount40_jl9s_core_194 | popcount40_jl9s_core_196;
  assign popcount40_jl9s_core_199 = input_a[24] ^ input_a[33];
  assign popcount40_jl9s_core_200 = ~input_a[10];
  assign popcount40_jl9s_core_201 = input_a[14] & popcount40_jl9s_core_191;
  assign popcount40_jl9s_core_202 = popcount40_jl9s_core_176 ^ popcount40_jl9s_core_195;
  assign popcount40_jl9s_core_203 = popcount40_jl9s_core_176 & popcount40_jl9s_core_195;
  assign popcount40_jl9s_core_204 = popcount40_jl9s_core_202 ^ popcount40_jl9s_core_201;
  assign popcount40_jl9s_core_205 = popcount40_jl9s_core_202 & popcount40_jl9s_core_201;
  assign popcount40_jl9s_core_206 = popcount40_jl9s_core_203 | popcount40_jl9s_core_205;
  assign popcount40_jl9s_core_207 = popcount40_jl9s_core_181 ^ popcount40_jl9s_core_197;
  assign popcount40_jl9s_core_208 = popcount40_jl9s_core_181 & popcount40_jl9s_core_197;
  assign popcount40_jl9s_core_209 = popcount40_jl9s_core_207 ^ popcount40_jl9s_core_206;
  assign popcount40_jl9s_core_210 = popcount40_jl9s_core_207 & popcount40_jl9s_core_206;
  assign popcount40_jl9s_core_211 = popcount40_jl9s_core_208 | popcount40_jl9s_core_210;
  assign popcount40_jl9s_core_215 = ~input_a[29];
  assign popcount40_jl9s_core_216 = input_a[13] | input_a[21];
  assign popcount40_jl9s_core_217 = ~input_a[34];
  assign popcount40_jl9s_core_218 = input_a[30] & input_a[26];
  assign popcount40_jl9s_core_221 = input_a[10] | input_a[2];
  assign popcount40_jl9s_core_222_not = ~input_a[9];
  assign popcount40_jl9s_core_223 = input_a[5] | input_a[34];
  assign popcount40_jl9s_core_225 = ~(input_a[31] & input_a[22]);
  assign popcount40_jl9s_core_227 = popcount40_jl9s_core_218 ^ popcount40_jl9s_core_223;
  assign popcount40_jl9s_core_228 = popcount40_jl9s_core_218 & popcount40_jl9s_core_223;
  assign popcount40_jl9s_core_229 = popcount40_jl9s_core_227 ^ input_a[3];
  assign popcount40_jl9s_core_230 = popcount40_jl9s_core_227 & input_a[3];
  assign popcount40_jl9s_core_231 = popcount40_jl9s_core_228 | popcount40_jl9s_core_230;
  assign popcount40_jl9s_core_235 = input_a[28] & input_a[15];
  assign popcount40_jl9s_core_236 = input_a[30] | input_a[1];
  assign popcount40_jl9s_core_238 = ~(input_a[19] ^ input_a[15]);
  assign popcount40_jl9s_core_239 = ~(input_a[23] | input_a[10]);
  assign popcount40_jl9s_core_241 = ~(input_a[28] & input_a[27]);
  assign popcount40_jl9s_core_245 = ~(input_a[24] | input_a[12]);
  assign popcount40_jl9s_core_246 = input_a[27] & input_a[34];
  assign popcount40_jl9s_core_247 = ~(input_a[4] & input_a[34]);
  assign popcount40_jl9s_core_248 = input_a[22] ^ input_a[23];
  assign popcount40_jl9s_core_250 = input_a[20] ^ input_a[4];
  assign popcount40_jl9s_core_251 = ~(input_a[8] ^ input_a[5]);
  assign popcount40_jl9s_core_253 = ~popcount40_jl9s_core_229;
  assign popcount40_jl9s_core_260 = popcount40_jl9s_core_231 ^ popcount40_jl9s_core_229;
  assign popcount40_jl9s_core_261 = popcount40_jl9s_core_231 & popcount40_jl9s_core_229;
  assign popcount40_jl9s_core_266 = ~(input_a[33] ^ input_a[10]);
  assign popcount40_jl9s_core_267 = ~input_a[32];
  assign popcount40_jl9s_core_268 = input_a[32] | input_a[25];
  assign popcount40_jl9s_core_269 = input_a[1] & input_a[16];
  assign popcount40_jl9s_core_270 = popcount40_jl9s_core_204 ^ popcount40_jl9s_core_253;
  assign popcount40_jl9s_core_271 = popcount40_jl9s_core_204 & popcount40_jl9s_core_253;
  assign popcount40_jl9s_core_272 = popcount40_jl9s_core_270 ^ popcount40_jl9s_core_269;
  assign popcount40_jl9s_core_273 = popcount40_jl9s_core_270 & popcount40_jl9s_core_269;
  assign popcount40_jl9s_core_274 = popcount40_jl9s_core_271 | popcount40_jl9s_core_273;
  assign popcount40_jl9s_core_275 = popcount40_jl9s_core_209 ^ popcount40_jl9s_core_260;
  assign popcount40_jl9s_core_276 = popcount40_jl9s_core_209 & popcount40_jl9s_core_260;
  assign popcount40_jl9s_core_277 = popcount40_jl9s_core_275 ^ popcount40_jl9s_core_274;
  assign popcount40_jl9s_core_278 = popcount40_jl9s_core_275 & popcount40_jl9s_core_274;
  assign popcount40_jl9s_core_279 = popcount40_jl9s_core_276 | popcount40_jl9s_core_278;
  assign popcount40_jl9s_core_280 = popcount40_jl9s_core_211 ^ popcount40_jl9s_core_261;
  assign popcount40_jl9s_core_281 = popcount40_jl9s_core_211 & popcount40_jl9s_core_261;
  assign popcount40_jl9s_core_282 = popcount40_jl9s_core_280 ^ popcount40_jl9s_core_279;
  assign popcount40_jl9s_core_283 = popcount40_jl9s_core_280 & popcount40_jl9s_core_279;
  assign popcount40_jl9s_core_284 = popcount40_jl9s_core_281 | popcount40_jl9s_core_283;
  assign popcount40_jl9s_core_286 = input_a[8] ^ input_a[29];
  assign popcount40_jl9s_core_290 = input_a[13] | input_a[13];
  assign popcount40_jl9s_core_291 = input_a[0] & input_a[4];
  assign popcount40_jl9s_core_292 = popcount40_jl9s_core_148 ^ popcount40_jl9s_core_272;
  assign popcount40_jl9s_core_293 = popcount40_jl9s_core_148 & popcount40_jl9s_core_272;
  assign popcount40_jl9s_core_294 = popcount40_jl9s_core_292 ^ popcount40_jl9s_core_291;
  assign popcount40_jl9s_core_295 = popcount40_jl9s_core_292 & popcount40_jl9s_core_291;
  assign popcount40_jl9s_core_296 = popcount40_jl9s_core_293 | popcount40_jl9s_core_295;
  assign popcount40_jl9s_core_297 = popcount40_jl9s_core_153 ^ popcount40_jl9s_core_277;
  assign popcount40_jl9s_core_298 = popcount40_jl9s_core_153 & popcount40_jl9s_core_277;
  assign popcount40_jl9s_core_299 = popcount40_jl9s_core_297 ^ popcount40_jl9s_core_296;
  assign popcount40_jl9s_core_300 = popcount40_jl9s_core_297 & popcount40_jl9s_core_296;
  assign popcount40_jl9s_core_301 = popcount40_jl9s_core_298 | popcount40_jl9s_core_300;
  assign popcount40_jl9s_core_302 = popcount40_jl9s_core_158 ^ popcount40_jl9s_core_282;
  assign popcount40_jl9s_core_303 = popcount40_jl9s_core_158 & popcount40_jl9s_core_282;
  assign popcount40_jl9s_core_304 = popcount40_jl9s_core_302 ^ popcount40_jl9s_core_301;
  assign popcount40_jl9s_core_305 = popcount40_jl9s_core_302 & popcount40_jl9s_core_301;
  assign popcount40_jl9s_core_306 = popcount40_jl9s_core_303 | popcount40_jl9s_core_305;
  assign popcount40_jl9s_core_308 = ~(input_a[15] ^ input_a[26]);
  assign popcount40_jl9s_core_309 = popcount40_jl9s_core_284 | popcount40_jl9s_core_306;
  assign popcount40_jl9s_core_310 = input_a[1] & input_a[29];
  assign popcount40_jl9s_core_311 = ~(input_a[21] ^ input_a[38]);
  assign popcount40_jl9s_core_313 = input_a[10] & input_a[27];
  assign popcount40_jl9s_core_315 = ~input_a[13];
  assign popcount40_jl9s_core_316 = input_a[39] & input_a[16];

  assign popcount40_jl9s_out[0] = input_a[27];
  assign popcount40_jl9s_out[1] = popcount40_jl9s_core_294;
  assign popcount40_jl9s_out[2] = popcount40_jl9s_core_299;
  assign popcount40_jl9s_out[3] = popcount40_jl9s_core_304;
  assign popcount40_jl9s_out[4] = popcount40_jl9s_core_309;
  assign popcount40_jl9s_out[5] = 1'b0;
endmodule