// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.56944
// WCE=24.0
// EP=0.975355%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_zdtu(input [26:0] input_a, output [4:0] popcount27_zdtu_out);
  wire popcount27_zdtu_core_032;
  wire popcount27_zdtu_core_035;
  wire popcount27_zdtu_core_037;
  wire popcount27_zdtu_core_038;
  wire popcount27_zdtu_core_039;
  wire popcount27_zdtu_core_040;
  wire popcount27_zdtu_core_041;
  wire popcount27_zdtu_core_043;
  wire popcount27_zdtu_core_044;
  wire popcount27_zdtu_core_047;
  wire popcount27_zdtu_core_049;
  wire popcount27_zdtu_core_051;
  wire popcount27_zdtu_core_052;
  wire popcount27_zdtu_core_054;
  wire popcount27_zdtu_core_055_not;
  wire popcount27_zdtu_core_056;
  wire popcount27_zdtu_core_057;
  wire popcount27_zdtu_core_062;
  wire popcount27_zdtu_core_063;
  wire popcount27_zdtu_core_064;
  wire popcount27_zdtu_core_065;
  wire popcount27_zdtu_core_066;
  wire popcount27_zdtu_core_067;
  wire popcount27_zdtu_core_068;
  wire popcount27_zdtu_core_071;
  wire popcount27_zdtu_core_073;
  wire popcount27_zdtu_core_076;
  wire popcount27_zdtu_core_079;
  wire popcount27_zdtu_core_083;
  wire popcount27_zdtu_core_084;
  wire popcount27_zdtu_core_086;
  wire popcount27_zdtu_core_088_not;
  wire popcount27_zdtu_core_089;
  wire popcount27_zdtu_core_091;
  wire popcount27_zdtu_core_093;
  wire popcount27_zdtu_core_095_not;
  wire popcount27_zdtu_core_097;
  wire popcount27_zdtu_core_098;
  wire popcount27_zdtu_core_099;
  wire popcount27_zdtu_core_101;
  wire popcount27_zdtu_core_102;
  wire popcount27_zdtu_core_103;
  wire popcount27_zdtu_core_105;
  wire popcount27_zdtu_core_108;
  wire popcount27_zdtu_core_109;
  wire popcount27_zdtu_core_112;
  wire popcount27_zdtu_core_114;
  wire popcount27_zdtu_core_115;
  wire popcount27_zdtu_core_119;
  wire popcount27_zdtu_core_120;
  wire popcount27_zdtu_core_121_not;
  wire popcount27_zdtu_core_122;
  wire popcount27_zdtu_core_124;
  wire popcount27_zdtu_core_125;
  wire popcount27_zdtu_core_129;
  wire popcount27_zdtu_core_130;
  wire popcount27_zdtu_core_132;
  wire popcount27_zdtu_core_133;
  wire popcount27_zdtu_core_134;
  wire popcount27_zdtu_core_135;
  wire popcount27_zdtu_core_137;
  wire popcount27_zdtu_core_138;
  wire popcount27_zdtu_core_139;
  wire popcount27_zdtu_core_142;
  wire popcount27_zdtu_core_144;
  wire popcount27_zdtu_core_148;
  wire popcount27_zdtu_core_150;
  wire popcount27_zdtu_core_152;
  wire popcount27_zdtu_core_153;
  wire popcount27_zdtu_core_154;
  wire popcount27_zdtu_core_155;
  wire popcount27_zdtu_core_156;
  wire popcount27_zdtu_core_159;
  wire popcount27_zdtu_core_161;
  wire popcount27_zdtu_core_162_not;
  wire popcount27_zdtu_core_163;
  wire popcount27_zdtu_core_170;
  wire popcount27_zdtu_core_171;
  wire popcount27_zdtu_core_172;
  wire popcount27_zdtu_core_173;
  wire popcount27_zdtu_core_174;
  wire popcount27_zdtu_core_177;
  wire popcount27_zdtu_core_179_not;
  wire popcount27_zdtu_core_181;
  wire popcount27_zdtu_core_182;
  wire popcount27_zdtu_core_184;
  wire popcount27_zdtu_core_185;
  wire popcount27_zdtu_core_187;
  wire popcount27_zdtu_core_188;
  wire popcount27_zdtu_core_191;
  wire popcount27_zdtu_core_192;
  wire popcount27_zdtu_core_193;
  wire popcount27_zdtu_core_194;

  assign popcount27_zdtu_core_032 = ~(input_a[18] ^ input_a[16]);
  assign popcount27_zdtu_core_035 = ~(input_a[12] | input_a[12]);
  assign popcount27_zdtu_core_037 = input_a[11] ^ input_a[19];
  assign popcount27_zdtu_core_038 = input_a[6] | input_a[13];
  assign popcount27_zdtu_core_039 = ~(input_a[25] ^ input_a[10]);
  assign popcount27_zdtu_core_040 = ~(input_a[24] ^ input_a[24]);
  assign popcount27_zdtu_core_041 = ~input_a[11];
  assign popcount27_zdtu_core_043 = input_a[2] & input_a[16];
  assign popcount27_zdtu_core_044 = input_a[2] & input_a[16];
  assign popcount27_zdtu_core_047 = ~(input_a[20] | input_a[25]);
  assign popcount27_zdtu_core_049 = input_a[7] & input_a[9];
  assign popcount27_zdtu_core_051 = ~(input_a[0] ^ input_a[3]);
  assign popcount27_zdtu_core_052 = input_a[26] & input_a[16];
  assign popcount27_zdtu_core_054 = ~(input_a[0] & input_a[18]);
  assign popcount27_zdtu_core_055_not = ~input_a[4];
  assign popcount27_zdtu_core_056 = input_a[0] ^ input_a[18];
  assign popcount27_zdtu_core_057 = ~(input_a[11] | input_a[6]);
  assign popcount27_zdtu_core_062 = ~(input_a[24] & input_a[12]);
  assign popcount27_zdtu_core_063 = ~(input_a[9] & input_a[4]);
  assign popcount27_zdtu_core_064 = input_a[8] ^ input_a[4];
  assign popcount27_zdtu_core_065 = input_a[15] ^ input_a[4];
  assign popcount27_zdtu_core_066 = ~input_a[7];
  assign popcount27_zdtu_core_067 = input_a[14] | input_a[13];
  assign popcount27_zdtu_core_068 = input_a[5] | input_a[0];
  assign popcount27_zdtu_core_071 = ~(input_a[19] ^ input_a[17]);
  assign popcount27_zdtu_core_073 = ~(input_a[11] | input_a[5]);
  assign popcount27_zdtu_core_076 = ~(input_a[1] & input_a[7]);
  assign popcount27_zdtu_core_079 = ~input_a[14];
  assign popcount27_zdtu_core_083 = input_a[17] ^ input_a[7];
  assign popcount27_zdtu_core_084 = ~(input_a[12] & input_a[17]);
  assign popcount27_zdtu_core_086 = ~(input_a[26] | input_a[19]);
  assign popcount27_zdtu_core_088_not = ~input_a[15];
  assign popcount27_zdtu_core_089 = input_a[10] | input_a[2];
  assign popcount27_zdtu_core_091 = input_a[18] & input_a[21];
  assign popcount27_zdtu_core_093 = ~(input_a[12] ^ input_a[6]);
  assign popcount27_zdtu_core_095_not = ~input_a[0];
  assign popcount27_zdtu_core_097 = input_a[21] ^ input_a[6];
  assign popcount27_zdtu_core_098 = ~(input_a[21] & input_a[23]);
  assign popcount27_zdtu_core_099 = ~input_a[24];
  assign popcount27_zdtu_core_101 = input_a[15] & input_a[9];
  assign popcount27_zdtu_core_102 = ~(input_a[18] & input_a[17]);
  assign popcount27_zdtu_core_103 = input_a[14] ^ input_a[15];
  assign popcount27_zdtu_core_105 = ~(input_a[14] | input_a[12]);
  assign popcount27_zdtu_core_108 = ~(input_a[26] & input_a[4]);
  assign popcount27_zdtu_core_109 = ~(input_a[12] ^ input_a[15]);
  assign popcount27_zdtu_core_112 = input_a[7] & input_a[24];
  assign popcount27_zdtu_core_114 = input_a[5] ^ input_a[7];
  assign popcount27_zdtu_core_115 = input_a[20] | input_a[12];
  assign popcount27_zdtu_core_119 = input_a[16] & input_a[5];
  assign popcount27_zdtu_core_120 = ~input_a[3];
  assign popcount27_zdtu_core_121_not = ~input_a[21];
  assign popcount27_zdtu_core_122 = input_a[9] ^ input_a[5];
  assign popcount27_zdtu_core_124 = input_a[13] & input_a[26];
  assign popcount27_zdtu_core_125 = ~(input_a[1] & input_a[24]);
  assign popcount27_zdtu_core_129 = ~(input_a[24] ^ input_a[15]);
  assign popcount27_zdtu_core_130 = input_a[8] ^ input_a[23];
  assign popcount27_zdtu_core_132 = ~(input_a[9] | input_a[23]);
  assign popcount27_zdtu_core_133 = input_a[11] | input_a[8];
  assign popcount27_zdtu_core_134 = input_a[23] ^ input_a[19];
  assign popcount27_zdtu_core_135 = ~(input_a[2] ^ input_a[9]);
  assign popcount27_zdtu_core_137 = input_a[4] ^ input_a[12];
  assign popcount27_zdtu_core_138 = ~(input_a[21] | input_a[1]);
  assign popcount27_zdtu_core_139 = ~input_a[6];
  assign popcount27_zdtu_core_142 = ~(input_a[17] & input_a[11]);
  assign popcount27_zdtu_core_144 = ~(input_a[13] ^ input_a[21]);
  assign popcount27_zdtu_core_148 = ~(input_a[24] | input_a[15]);
  assign popcount27_zdtu_core_150 = ~(input_a[18] & input_a[22]);
  assign popcount27_zdtu_core_152 = ~(input_a[2] & input_a[24]);
  assign popcount27_zdtu_core_153 = ~input_a[3];
  assign popcount27_zdtu_core_154 = ~(input_a[2] | input_a[22]);
  assign popcount27_zdtu_core_155 = input_a[15] ^ input_a[15];
  assign popcount27_zdtu_core_156 = ~input_a[7];
  assign popcount27_zdtu_core_159 = ~(input_a[9] | input_a[3]);
  assign popcount27_zdtu_core_161 = ~(input_a[6] & input_a[0]);
  assign popcount27_zdtu_core_162_not = ~input_a[6];
  assign popcount27_zdtu_core_163 = ~input_a[0];
  assign popcount27_zdtu_core_170 = input_a[17] ^ input_a[2];
  assign popcount27_zdtu_core_171 = ~(input_a[9] & input_a[8]);
  assign popcount27_zdtu_core_172 = ~(input_a[6] ^ input_a[24]);
  assign popcount27_zdtu_core_173 = ~(input_a[4] & input_a[23]);
  assign popcount27_zdtu_core_174 = ~(input_a[6] & input_a[7]);
  assign popcount27_zdtu_core_177 = ~(input_a[20] | input_a[13]);
  assign popcount27_zdtu_core_179_not = ~input_a[9];
  assign popcount27_zdtu_core_181 = input_a[2] ^ input_a[24];
  assign popcount27_zdtu_core_182 = ~(input_a[1] | input_a[24]);
  assign popcount27_zdtu_core_184 = ~(input_a[24] ^ input_a[26]);
  assign popcount27_zdtu_core_185 = ~(input_a[20] ^ input_a[7]);
  assign popcount27_zdtu_core_187 = input_a[26] | input_a[25];
  assign popcount27_zdtu_core_188 = ~input_a[17];
  assign popcount27_zdtu_core_191 = input_a[0] ^ input_a[9];
  assign popcount27_zdtu_core_192 = ~(input_a[20] & input_a[15]);
  assign popcount27_zdtu_core_193 = input_a[24] & input_a[15];
  assign popcount27_zdtu_core_194 = ~(input_a[6] | input_a[22]);

  assign popcount27_zdtu_out[0] = input_a[21];
  assign popcount27_zdtu_out[1] = input_a[21];
  assign popcount27_zdtu_out[2] = 1'b0;
  assign popcount27_zdtu_out[3] = input_a[26];
  assign popcount27_zdtu_out[4] = input_a[24];
endmodule