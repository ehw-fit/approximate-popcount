// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.61776
// WCE=6.0
// EP=0.812671%
// Printed PDK parameters:
//  Area=46814884.0
//  Delay=70635768.0
//  Power=2511000.0

module popcount28_jzqm(input [27:0] input_a, output [4:0] popcount28_jzqm_out);
  wire popcount28_jzqm_core_030;
  wire popcount28_jzqm_core_031;
  wire popcount28_jzqm_core_032;
  wire popcount28_jzqm_core_033;
  wire popcount28_jzqm_core_034;
  wire popcount28_jzqm_core_036;
  wire popcount28_jzqm_core_037;
  wire popcount28_jzqm_core_038;
  wire popcount28_jzqm_core_039;
  wire popcount28_jzqm_core_041;
  wire popcount28_jzqm_core_042;
  wire popcount28_jzqm_core_043;
  wire popcount28_jzqm_core_044;
  wire popcount28_jzqm_core_045;
  wire popcount28_jzqm_core_047;
  wire popcount28_jzqm_core_048;
  wire popcount28_jzqm_core_049;
  wire popcount28_jzqm_core_050;
  wire popcount28_jzqm_core_056;
  wire popcount28_jzqm_core_058;
  wire popcount28_jzqm_core_059;
  wire popcount28_jzqm_core_060;
  wire popcount28_jzqm_core_062;
  wire popcount28_jzqm_core_063;
  wire popcount28_jzqm_core_066;
  wire popcount28_jzqm_core_067;
  wire popcount28_jzqm_core_068;
  wire popcount28_jzqm_core_070;
  wire popcount28_jzqm_core_071;
  wire popcount28_jzqm_core_073;
  wire popcount28_jzqm_core_074;
  wire popcount28_jzqm_core_075;
  wire popcount28_jzqm_core_077;
  wire popcount28_jzqm_core_082;
  wire popcount28_jzqm_core_083;
  wire popcount28_jzqm_core_084;
  wire popcount28_jzqm_core_085;
  wire popcount28_jzqm_core_086;
  wire popcount28_jzqm_core_088;
  wire popcount28_jzqm_core_089;
  wire popcount28_jzqm_core_090_not;
  wire popcount28_jzqm_core_093;
  wire popcount28_jzqm_core_097;
  wire popcount28_jzqm_core_098;
  wire popcount28_jzqm_core_101;
  wire popcount28_jzqm_core_104;
  wire popcount28_jzqm_core_105;
  wire popcount28_jzqm_core_106;
  wire popcount28_jzqm_core_107;
  wire popcount28_jzqm_core_108;
  wire popcount28_jzqm_core_109;
  wire popcount28_jzqm_core_111;
  wire popcount28_jzqm_core_112;
  wire popcount28_jzqm_core_113;
  wire popcount28_jzqm_core_114;
  wire popcount28_jzqm_core_115;
  wire popcount28_jzqm_core_116;
  wire popcount28_jzqm_core_117;
  wire popcount28_jzqm_core_118;
  wire popcount28_jzqm_core_119;
  wire popcount28_jzqm_core_120;
  wire popcount28_jzqm_core_122;
  wire popcount28_jzqm_core_123;
  wire popcount28_jzqm_core_124;
  wire popcount28_jzqm_core_125;
  wire popcount28_jzqm_core_126;
  wire popcount28_jzqm_core_127;
  wire popcount28_jzqm_core_128;
  wire popcount28_jzqm_core_131;
  wire popcount28_jzqm_core_132;
  wire popcount28_jzqm_core_134;
  wire popcount28_jzqm_core_135;
  wire popcount28_jzqm_core_136;
  wire popcount28_jzqm_core_137;
  wire popcount28_jzqm_core_138;
  wire popcount28_jzqm_core_141;
  wire popcount28_jzqm_core_143;
  wire popcount28_jzqm_core_148;
  wire popcount28_jzqm_core_150;
  wire popcount28_jzqm_core_151;
  wire popcount28_jzqm_core_152;
  wire popcount28_jzqm_core_155;
  wire popcount28_jzqm_core_156;
  wire popcount28_jzqm_core_160;
  wire popcount28_jzqm_core_161;
  wire popcount28_jzqm_core_163;
  wire popcount28_jzqm_core_164;
  wire popcount28_jzqm_core_165;
  wire popcount28_jzqm_core_166;
  wire popcount28_jzqm_core_167;
  wire popcount28_jzqm_core_168;
  wire popcount28_jzqm_core_169;
  wire popcount28_jzqm_core_170;
  wire popcount28_jzqm_core_172;
  wire popcount28_jzqm_core_173;
  wire popcount28_jzqm_core_174;
  wire popcount28_jzqm_core_176;
  wire popcount28_jzqm_core_177;
  wire popcount28_jzqm_core_178;
  wire popcount28_jzqm_core_179;
  wire popcount28_jzqm_core_180;
  wire popcount28_jzqm_core_181;
  wire popcount28_jzqm_core_182;
  wire popcount28_jzqm_core_183;
  wire popcount28_jzqm_core_184;
  wire popcount28_jzqm_core_185;
  wire popcount28_jzqm_core_186;
  wire popcount28_jzqm_core_187;
  wire popcount28_jzqm_core_188;
  wire popcount28_jzqm_core_189;
  wire popcount28_jzqm_core_190;
  wire popcount28_jzqm_core_191;
  wire popcount28_jzqm_core_192;
  wire popcount28_jzqm_core_193;
  wire popcount28_jzqm_core_194;
  wire popcount28_jzqm_core_195;
  wire popcount28_jzqm_core_196;
  wire popcount28_jzqm_core_198;
  wire popcount28_jzqm_core_199;
  wire popcount28_jzqm_core_200;

  assign popcount28_jzqm_core_030 = ~(input_a[4] & input_a[12]);
  assign popcount28_jzqm_core_031 = input_a[1] & input_a[12];
  assign popcount28_jzqm_core_032 = ~(input_a[13] ^ input_a[1]);
  assign popcount28_jzqm_core_033 = input_a[0] & input_a[6];
  assign popcount28_jzqm_core_034 = popcount28_jzqm_core_031 | popcount28_jzqm_core_033;
  assign popcount28_jzqm_core_036 = ~(input_a[18] ^ input_a[21]);
  assign popcount28_jzqm_core_037 = input_a[3] & input_a[4];
  assign popcount28_jzqm_core_038 = input_a[2] ^ input_a[3];
  assign popcount28_jzqm_core_039 = input_a[5] & input_a[11];
  assign popcount28_jzqm_core_041 = input_a[2] & input_a[7];
  assign popcount28_jzqm_core_042 = popcount28_jzqm_core_037 | popcount28_jzqm_core_039;
  assign popcount28_jzqm_core_043 = popcount28_jzqm_core_037 & popcount28_jzqm_core_039;
  assign popcount28_jzqm_core_044 = popcount28_jzqm_core_042 | popcount28_jzqm_core_041;
  assign popcount28_jzqm_core_045 = input_a[23] | input_a[9];
  assign popcount28_jzqm_core_047 = ~(input_a[24] ^ input_a[12]);
  assign popcount28_jzqm_core_048 = ~(input_a[10] ^ input_a[5]);
  assign popcount28_jzqm_core_049 = ~(input_a[12] & input_a[26]);
  assign popcount28_jzqm_core_050 = popcount28_jzqm_core_034 & popcount28_jzqm_core_044;
  assign popcount28_jzqm_core_056 = popcount28_jzqm_core_043 | popcount28_jzqm_core_050;
  assign popcount28_jzqm_core_058 = input_a[18] | input_a[21];
  assign popcount28_jzqm_core_059 = ~(input_a[15] ^ input_a[8]);
  assign popcount28_jzqm_core_060 = input_a[8] & input_a[9];
  assign popcount28_jzqm_core_062 = input_a[26] & input_a[24];
  assign popcount28_jzqm_core_063 = popcount28_jzqm_core_060 | popcount28_jzqm_core_062;
  assign popcount28_jzqm_core_066 = ~(input_a[13] & input_a[23]);
  assign popcount28_jzqm_core_067 = ~(input_a[10] | input_a[19]);
  assign popcount28_jzqm_core_068 = ~(input_a[3] & input_a[25]);
  assign popcount28_jzqm_core_070 = ~(input_a[20] ^ input_a[10]);
  assign popcount28_jzqm_core_071 = input_a[24] ^ input_a[13];
  assign popcount28_jzqm_core_073 = input_a[27] & input_a[22];
  assign popcount28_jzqm_core_074 = ~(input_a[1] & input_a[21]);
  assign popcount28_jzqm_core_075 = ~(input_a[13] & input_a[19]);
  assign popcount28_jzqm_core_077 = ~(input_a[7] ^ input_a[21]);
  assign popcount28_jzqm_core_082 = input_a[12] | input_a[11];
  assign popcount28_jzqm_core_083 = input_a[16] | input_a[21];
  assign popcount28_jzqm_core_084 = input_a[14] & input_a[18];
  assign popcount28_jzqm_core_085 = ~(input_a[23] ^ input_a[16]);
  assign popcount28_jzqm_core_086 = ~input_a[18];
  assign popcount28_jzqm_core_088 = ~(input_a[2] | input_a[14]);
  assign popcount28_jzqm_core_089 = ~(input_a[19] | input_a[27]);
  assign popcount28_jzqm_core_090_not = ~popcount28_jzqm_core_063;
  assign popcount28_jzqm_core_093 = ~popcount28_jzqm_core_090_not;
  assign popcount28_jzqm_core_097 = popcount28_jzqm_core_056 ^ popcount28_jzqm_core_093;
  assign popcount28_jzqm_core_098 = popcount28_jzqm_core_056 & popcount28_jzqm_core_093;
  assign popcount28_jzqm_core_101 = input_a[12] & input_a[19];
  assign popcount28_jzqm_core_104 = input_a[11] ^ input_a[20];
  assign popcount28_jzqm_core_105 = input_a[15] ^ input_a[16];
  assign popcount28_jzqm_core_106 = input_a[15] & input_a[16];
  assign popcount28_jzqm_core_107 = input_a[14] ^ popcount28_jzqm_core_105;
  assign popcount28_jzqm_core_108 = input_a[14] & popcount28_jzqm_core_105;
  assign popcount28_jzqm_core_109 = popcount28_jzqm_core_106 | popcount28_jzqm_core_108;
  assign popcount28_jzqm_core_111 = input_a[17] ^ input_a[18];
  assign popcount28_jzqm_core_112 = input_a[17] & input_a[18];
  assign popcount28_jzqm_core_113 = input_a[19] ^ input_a[20];
  assign popcount28_jzqm_core_114 = input_a[19] & input_a[20];
  assign popcount28_jzqm_core_115 = popcount28_jzqm_core_111 ^ popcount28_jzqm_core_113;
  assign popcount28_jzqm_core_116 = popcount28_jzqm_core_111 & popcount28_jzqm_core_113;
  assign popcount28_jzqm_core_117 = popcount28_jzqm_core_112 ^ popcount28_jzqm_core_114;
  assign popcount28_jzqm_core_118 = popcount28_jzqm_core_112 & popcount28_jzqm_core_114;
  assign popcount28_jzqm_core_119 = popcount28_jzqm_core_117 | popcount28_jzqm_core_116;
  assign popcount28_jzqm_core_120 = input_a[16] | input_a[21];
  assign popcount28_jzqm_core_122 = popcount28_jzqm_core_107 ^ popcount28_jzqm_core_115;
  assign popcount28_jzqm_core_123 = popcount28_jzqm_core_107 & popcount28_jzqm_core_115;
  assign popcount28_jzqm_core_124 = popcount28_jzqm_core_109 ^ popcount28_jzqm_core_119;
  assign popcount28_jzqm_core_125 = popcount28_jzqm_core_109 & popcount28_jzqm_core_119;
  assign popcount28_jzqm_core_126 = popcount28_jzqm_core_124 ^ popcount28_jzqm_core_123;
  assign popcount28_jzqm_core_127 = popcount28_jzqm_core_124 & popcount28_jzqm_core_123;
  assign popcount28_jzqm_core_128 = popcount28_jzqm_core_125 | popcount28_jzqm_core_127;
  assign popcount28_jzqm_core_131 = popcount28_jzqm_core_118 | popcount28_jzqm_core_128;
  assign popcount28_jzqm_core_132 = ~input_a[19];
  assign popcount28_jzqm_core_134 = input_a[22] ^ input_a[23];
  assign popcount28_jzqm_core_135 = input_a[22] & input_a[23];
  assign popcount28_jzqm_core_136 = input_a[21] ^ popcount28_jzqm_core_134;
  assign popcount28_jzqm_core_137 = input_a[21] & popcount28_jzqm_core_134;
  assign popcount28_jzqm_core_138 = popcount28_jzqm_core_135 | popcount28_jzqm_core_137;
  assign popcount28_jzqm_core_141 = ~(input_a[21] | input_a[15]);
  assign popcount28_jzqm_core_143 = input_a[25] & input_a[27];
  assign popcount28_jzqm_core_148 = ~(input_a[8] | input_a[10]);
  assign popcount28_jzqm_core_150 = ~input_a[22];
  assign popcount28_jzqm_core_151 = popcount28_jzqm_core_136 ^ input_a[10];
  assign popcount28_jzqm_core_152 = popcount28_jzqm_core_136 & input_a[10];
  assign popcount28_jzqm_core_155 = popcount28_jzqm_core_138 ^ popcount28_jzqm_core_152;
  assign popcount28_jzqm_core_156 = input_a[22] & popcount28_jzqm_core_152;
  assign popcount28_jzqm_core_160 = ~(input_a[21] & popcount28_jzqm_core_156);
  assign popcount28_jzqm_core_161 = input_a[23] & popcount28_jzqm_core_156;
  assign popcount28_jzqm_core_163 = popcount28_jzqm_core_122 ^ popcount28_jzqm_core_151;
  assign popcount28_jzqm_core_164 = popcount28_jzqm_core_122 & popcount28_jzqm_core_151;
  assign popcount28_jzqm_core_165 = popcount28_jzqm_core_126 ^ popcount28_jzqm_core_155;
  assign popcount28_jzqm_core_166 = popcount28_jzqm_core_126 & popcount28_jzqm_core_155;
  assign popcount28_jzqm_core_167 = popcount28_jzqm_core_165 ^ popcount28_jzqm_core_164;
  assign popcount28_jzqm_core_168 = popcount28_jzqm_core_165 & popcount28_jzqm_core_164;
  assign popcount28_jzqm_core_169 = popcount28_jzqm_core_166 | popcount28_jzqm_core_168;
  assign popcount28_jzqm_core_170 = popcount28_jzqm_core_131 ^ popcount28_jzqm_core_160;
  assign popcount28_jzqm_core_172 = popcount28_jzqm_core_170 ^ popcount28_jzqm_core_169;
  assign popcount28_jzqm_core_173 = popcount28_jzqm_core_170 & popcount28_jzqm_core_169;
  assign popcount28_jzqm_core_174 = popcount28_jzqm_core_131 | popcount28_jzqm_core_173;
  assign popcount28_jzqm_core_176 = input_a[25] | input_a[6];
  assign popcount28_jzqm_core_177 = popcount28_jzqm_core_161 | popcount28_jzqm_core_174;
  assign popcount28_jzqm_core_178 = input_a[2] & input_a[5];
  assign popcount28_jzqm_core_179 = ~(input_a[24] & input_a[5]);
  assign popcount28_jzqm_core_180 = input_a[13] ^ popcount28_jzqm_core_163;
  assign popcount28_jzqm_core_181 = input_a[13] & popcount28_jzqm_core_163;
  assign popcount28_jzqm_core_182 = popcount28_jzqm_core_090_not | popcount28_jzqm_core_167;
  assign popcount28_jzqm_core_183 = popcount28_jzqm_core_090_not & popcount28_jzqm_core_167;
  assign popcount28_jzqm_core_184 = ~(input_a[5] ^ input_a[11]);
  assign popcount28_jzqm_core_185 = popcount28_jzqm_core_182 & popcount28_jzqm_core_181;
  assign popcount28_jzqm_core_186 = popcount28_jzqm_core_183 | popcount28_jzqm_core_185;
  assign popcount28_jzqm_core_187 = popcount28_jzqm_core_097 ^ popcount28_jzqm_core_172;
  assign popcount28_jzqm_core_188 = popcount28_jzqm_core_097 & popcount28_jzqm_core_172;
  assign popcount28_jzqm_core_189 = popcount28_jzqm_core_187 ^ popcount28_jzqm_core_186;
  assign popcount28_jzqm_core_190 = popcount28_jzqm_core_187 & popcount28_jzqm_core_186;
  assign popcount28_jzqm_core_191 = popcount28_jzqm_core_188 | popcount28_jzqm_core_190;
  assign popcount28_jzqm_core_192 = popcount28_jzqm_core_098 ^ popcount28_jzqm_core_177;
  assign popcount28_jzqm_core_193 = popcount28_jzqm_core_098 & popcount28_jzqm_core_177;
  assign popcount28_jzqm_core_194 = popcount28_jzqm_core_192 ^ popcount28_jzqm_core_191;
  assign popcount28_jzqm_core_195 = popcount28_jzqm_core_192 & popcount28_jzqm_core_191;
  assign popcount28_jzqm_core_196 = popcount28_jzqm_core_193 | popcount28_jzqm_core_195;
  assign popcount28_jzqm_core_198 = input_a[18] & input_a[15];
  assign popcount28_jzqm_core_199 = ~(input_a[23] & input_a[7]);
  assign popcount28_jzqm_core_200 = ~(input_a[21] | input_a[7]);

  assign popcount28_jzqm_out[0] = popcount28_jzqm_core_180;
  assign popcount28_jzqm_out[1] = popcount28_jzqm_core_143;
  assign popcount28_jzqm_out[2] = popcount28_jzqm_core_189;
  assign popcount28_jzqm_out[3] = popcount28_jzqm_core_194;
  assign popcount28_jzqm_out[4] = popcount28_jzqm_core_196;
endmodule