// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.3151
// WCE=19.0
// EP=0.863499%
// Printed PDK parameters:
//  Area=108258289.0
//  Delay=96904376.0
//  Power=5299300.0

module popcount47_atj4(input [46:0] input_a, output [5:0] popcount47_atj4_out);
  wire popcount47_atj4_core_050;
  wire popcount47_atj4_core_051;
  wire popcount47_atj4_core_052;
  wire popcount47_atj4_core_053;
  wire popcount47_atj4_core_054;
  wire popcount47_atj4_core_056;
  wire popcount47_atj4_core_059;
  wire popcount47_atj4_core_061;
  wire popcount47_atj4_core_062;
  wire popcount47_atj4_core_063;
  wire popcount47_atj4_core_064;
  wire popcount47_atj4_core_065;
  wire popcount47_atj4_core_066;
  wire popcount47_atj4_core_067;
  wire popcount47_atj4_core_068;
  wire popcount47_atj4_core_069;
  wire popcount47_atj4_core_070;
  wire popcount47_atj4_core_071;
  wire popcount47_atj4_core_072;
  wire popcount47_atj4_core_073;
  wire popcount47_atj4_core_074;
  wire popcount47_atj4_core_075;
  wire popcount47_atj4_core_076;
  wire popcount47_atj4_core_079;
  wire popcount47_atj4_core_080;
  wire popcount47_atj4_core_081;
  wire popcount47_atj4_core_082;
  wire popcount47_atj4_core_083;
  wire popcount47_atj4_core_084;
  wire popcount47_atj4_core_086;
  wire popcount47_atj4_core_087;
  wire popcount47_atj4_core_092;
  wire popcount47_atj4_core_093;
  wire popcount47_atj4_core_097;
  wire popcount47_atj4_core_098;
  wire popcount47_atj4_core_099;
  wire popcount47_atj4_core_100;
  wire popcount47_atj4_core_101;
  wire popcount47_atj4_core_104;
  wire popcount47_atj4_core_105;
  wire popcount47_atj4_core_107;
  wire popcount47_atj4_core_108;
  wire popcount47_atj4_core_109;
  wire popcount47_atj4_core_110;
  wire popcount47_atj4_core_111;
  wire popcount47_atj4_core_112;
  wire popcount47_atj4_core_113;
  wire popcount47_atj4_core_114;
  wire popcount47_atj4_core_115;
  wire popcount47_atj4_core_116;
  wire popcount47_atj4_core_117;
  wire popcount47_atj4_core_118;
  wire popcount47_atj4_core_119;
  wire popcount47_atj4_core_120;
  wire popcount47_atj4_core_121;
  wire popcount47_atj4_core_122;
  wire popcount47_atj4_core_123;
  wire popcount47_atj4_core_124;
  wire popcount47_atj4_core_125;
  wire popcount47_atj4_core_127;
  wire popcount47_atj4_core_128;
  wire popcount47_atj4_core_131;
  wire popcount47_atj4_core_132;
  wire popcount47_atj4_core_133;
  wire popcount47_atj4_core_137;
  wire popcount47_atj4_core_140;
  wire popcount47_atj4_core_144;
  wire popcount47_atj4_core_146;
  wire popcount47_atj4_core_155;
  wire popcount47_atj4_core_156;
  wire popcount47_atj4_core_159;
  wire popcount47_atj4_core_160;
  wire popcount47_atj4_core_162;
  wire popcount47_atj4_core_163;
  wire popcount47_atj4_core_164;
  wire popcount47_atj4_core_165;
  wire popcount47_atj4_core_166;
  wire popcount47_atj4_core_172;
  wire popcount47_atj4_core_173;
  wire popcount47_atj4_core_174;
  wire popcount47_atj4_core_175;
  wire popcount47_atj4_core_176;
  wire popcount47_atj4_core_177;
  wire popcount47_atj4_core_178;
  wire popcount47_atj4_core_179;
  wire popcount47_atj4_core_180;
  wire popcount47_atj4_core_181;
  wire popcount47_atj4_core_182;
  wire popcount47_atj4_core_183;
  wire popcount47_atj4_core_184;
  wire popcount47_atj4_core_185;
  wire popcount47_atj4_core_186;
  wire popcount47_atj4_core_187;
  wire popcount47_atj4_core_188;
  wire popcount47_atj4_core_191;
  wire popcount47_atj4_core_195;
  wire popcount47_atj4_core_200;
  wire popcount47_atj4_core_201;
  wire popcount47_atj4_core_203;
  wire popcount47_atj4_core_205;
  wire popcount47_atj4_core_208_not;
  wire popcount47_atj4_core_214;
  wire popcount47_atj4_core_215;
  wire popcount47_atj4_core_218;
  wire popcount47_atj4_core_219;
  wire popcount47_atj4_core_220;
  wire popcount47_atj4_core_221;
  wire popcount47_atj4_core_222;
  wire popcount47_atj4_core_224;
  wire popcount47_atj4_core_225;
  wire popcount47_atj4_core_226;
  wire popcount47_atj4_core_228;
  wire popcount47_atj4_core_230;
  wire popcount47_atj4_core_231;
  wire popcount47_atj4_core_232;
  wire popcount47_atj4_core_233;
  wire popcount47_atj4_core_238;
  wire popcount47_atj4_core_242;
  wire popcount47_atj4_core_243;
  wire popcount47_atj4_core_244;
  wire popcount47_atj4_core_245;
  wire popcount47_atj4_core_246;
  wire popcount47_atj4_core_247;
  wire popcount47_atj4_core_248;
  wire popcount47_atj4_core_249;
  wire popcount47_atj4_core_250;
  wire popcount47_atj4_core_251;
  wire popcount47_atj4_core_252;
  wire popcount47_atj4_core_253;
  wire popcount47_atj4_core_256;
  wire popcount47_atj4_core_257;
  wire popcount47_atj4_core_259;
  wire popcount47_atj4_core_260;
  wire popcount47_atj4_core_261;
  wire popcount47_atj4_core_262;
  wire popcount47_atj4_core_263;
  wire popcount47_atj4_core_264;
  wire popcount47_atj4_core_266;
  wire popcount47_atj4_core_267;
  wire popcount47_atj4_core_271;
  wire popcount47_atj4_core_272;
  wire popcount47_atj4_core_273;
  wire popcount47_atj4_core_274;
  wire popcount47_atj4_core_275;
  wire popcount47_atj4_core_276;
  wire popcount47_atj4_core_277;
  wire popcount47_atj4_core_280;
  wire popcount47_atj4_core_281;
  wire popcount47_atj4_core_283;
  wire popcount47_atj4_core_284;
  wire popcount47_atj4_core_285;
  wire popcount47_atj4_core_286;
  wire popcount47_atj4_core_287;
  wire popcount47_atj4_core_290;
  wire popcount47_atj4_core_291;
  wire popcount47_atj4_core_292;
  wire popcount47_atj4_core_293;
  wire popcount47_atj4_core_294;
  wire popcount47_atj4_core_296;
  wire popcount47_atj4_core_297;
  wire popcount47_atj4_core_298;
  wire popcount47_atj4_core_299;
  wire popcount47_atj4_core_300;
  wire popcount47_atj4_core_301;
  wire popcount47_atj4_core_304;
  wire popcount47_atj4_core_309;
  wire popcount47_atj4_core_310;
  wire popcount47_atj4_core_311;
  wire popcount47_atj4_core_312;
  wire popcount47_atj4_core_313;
  wire popcount47_atj4_core_314;
  wire popcount47_atj4_core_315;
  wire popcount47_atj4_core_316;
  wire popcount47_atj4_core_317;
  wire popcount47_atj4_core_318;
  wire popcount47_atj4_core_321;
  wire popcount47_atj4_core_322;
  wire popcount47_atj4_core_323;
  wire popcount47_atj4_core_326;
  wire popcount47_atj4_core_327;
  wire popcount47_atj4_core_328;
  wire popcount47_atj4_core_329;
  wire popcount47_atj4_core_330;
  wire popcount47_atj4_core_331;
  wire popcount47_atj4_core_332;
  wire popcount47_atj4_core_333;
  wire popcount47_atj4_core_334;
  wire popcount47_atj4_core_335;
  wire popcount47_atj4_core_336;
  wire popcount47_atj4_core_337;
  wire popcount47_atj4_core_338;
  wire popcount47_atj4_core_339;
  wire popcount47_atj4_core_340;
  wire popcount47_atj4_core_343;
  wire popcount47_atj4_core_344;
  wire popcount47_atj4_core_347;
  wire popcount47_atj4_core_348;
  wire popcount47_atj4_core_349;
  wire popcount47_atj4_core_350;
  wire popcount47_atj4_core_351;
  wire popcount47_atj4_core_352;
  wire popcount47_atj4_core_353;
  wire popcount47_atj4_core_354;
  wire popcount47_atj4_core_355;
  wire popcount47_atj4_core_356;
  wire popcount47_atj4_core_357;
  wire popcount47_atj4_core_358;
  wire popcount47_atj4_core_359;
  wire popcount47_atj4_core_360;
  wire popcount47_atj4_core_361;
  wire popcount47_atj4_core_362;
  wire popcount47_atj4_core_363;
  wire popcount47_atj4_core_364;
  wire popcount47_atj4_core_365;
  wire popcount47_atj4_core_366;
  wire popcount47_atj4_core_367;
  wire popcount47_atj4_core_368;
  wire popcount47_atj4_core_369;
  wire popcount47_atj4_core_370;
  wire popcount47_atj4_core_371;
  wire popcount47_atj4_core_372;

  assign popcount47_atj4_core_050 = input_a[0] & input_a[1];
  assign popcount47_atj4_core_051 = input_a[3] ^ input_a[4];
  assign popcount47_atj4_core_052 = input_a[3] & input_a[4];
  assign popcount47_atj4_core_053 = input_a[39] ^ popcount47_atj4_core_051;
  assign popcount47_atj4_core_054 = input_a[11] & popcount47_atj4_core_051;
  assign popcount47_atj4_core_056 = popcount47_atj4_core_052 & popcount47_atj4_core_054;
  assign popcount47_atj4_core_059 = ~(popcount47_atj4_core_050 & input_a[42]);
  assign popcount47_atj4_core_061 = popcount47_atj4_core_059 ^ input_a[0];
  assign popcount47_atj4_core_062 = popcount47_atj4_core_059 & input_a[0];
  assign popcount47_atj4_core_063 = popcount47_atj4_core_050 | popcount47_atj4_core_062;
  assign popcount47_atj4_core_064 = popcount47_atj4_core_056 | popcount47_atj4_core_063;
  assign popcount47_atj4_core_065 = popcount47_atj4_core_056 & input_a[7];
  assign popcount47_atj4_core_066 = input_a[6] ^ input_a[7];
  assign popcount47_atj4_core_067 = input_a[6] & input_a[7];
  assign popcount47_atj4_core_068 = input_a[5] | popcount47_atj4_core_066;
  assign popcount47_atj4_core_069 = input_a[5] & popcount47_atj4_core_066;
  assign popcount47_atj4_core_070 = popcount47_atj4_core_067 ^ popcount47_atj4_core_069;
  assign popcount47_atj4_core_071 = popcount47_atj4_core_067 & popcount47_atj4_core_069;
  assign popcount47_atj4_core_072 = input_a[9] ^ input_a[10];
  assign popcount47_atj4_core_073 = input_a[9] & input_a[10];
  assign popcount47_atj4_core_074 = input_a[8] ^ popcount47_atj4_core_072;
  assign popcount47_atj4_core_075 = input_a[8] & popcount47_atj4_core_072;
  assign popcount47_atj4_core_076 = popcount47_atj4_core_073 ^ popcount47_atj4_core_075;
  assign popcount47_atj4_core_079 = input_a[40] & popcount47_atj4_core_074;
  assign popcount47_atj4_core_080 = popcount47_atj4_core_070 ^ popcount47_atj4_core_076;
  assign popcount47_atj4_core_081 = popcount47_atj4_core_070 & popcount47_atj4_core_076;
  assign popcount47_atj4_core_082 = popcount47_atj4_core_080 ^ popcount47_atj4_core_079;
  assign popcount47_atj4_core_083 = popcount47_atj4_core_080 & popcount47_atj4_core_079;
  assign popcount47_atj4_core_084 = popcount47_atj4_core_081 | popcount47_atj4_core_083;
  assign popcount47_atj4_core_086 = ~input_a[46];
  assign popcount47_atj4_core_087 = popcount47_atj4_core_071 ^ popcount47_atj4_core_084;
  assign popcount47_atj4_core_092 = popcount47_atj4_core_061 ^ popcount47_atj4_core_082;
  assign popcount47_atj4_core_093 = popcount47_atj4_core_061 & popcount47_atj4_core_082;
  assign popcount47_atj4_core_097 = input_a[0] ^ popcount47_atj4_core_087;
  assign popcount47_atj4_core_098 = popcount47_atj4_core_064 & popcount47_atj4_core_087;
  assign popcount47_atj4_core_099 = popcount47_atj4_core_097 ^ popcount47_atj4_core_093;
  assign popcount47_atj4_core_100 = popcount47_atj4_core_097 & popcount47_atj4_core_093;
  assign popcount47_atj4_core_101 = popcount47_atj4_core_098 | popcount47_atj4_core_100;
  assign popcount47_atj4_core_104 = popcount47_atj4_core_065 ^ popcount47_atj4_core_101;
  assign popcount47_atj4_core_105 = popcount47_atj4_core_065 & input_a[4];
  assign popcount47_atj4_core_107 = input_a[12] ^ input_a[13];
  assign popcount47_atj4_core_108 = input_a[12] & input_a[13];
  assign popcount47_atj4_core_109 = input_a[11] ^ popcount47_atj4_core_107;
  assign popcount47_atj4_core_110 = input_a[11] & popcount47_atj4_core_107;
  assign popcount47_atj4_core_111 = popcount47_atj4_core_108 ^ popcount47_atj4_core_110;
  assign popcount47_atj4_core_112 = popcount47_atj4_core_108 & popcount47_atj4_core_110;
  assign popcount47_atj4_core_113 = input_a[15] ^ input_a[16];
  assign popcount47_atj4_core_114 = input_a[15] & input_a[16];
  assign popcount47_atj4_core_115 = input_a[14] ^ popcount47_atj4_core_113;
  assign popcount47_atj4_core_116 = input_a[14] & popcount47_atj4_core_113;
  assign popcount47_atj4_core_117 = popcount47_atj4_core_114 ^ popcount47_atj4_core_116;
  assign popcount47_atj4_core_118 = popcount47_atj4_core_114 & input_a[33];
  assign popcount47_atj4_core_119 = popcount47_atj4_core_109 ^ popcount47_atj4_core_115;
  assign popcount47_atj4_core_120 = popcount47_atj4_core_109 & popcount47_atj4_core_115;
  assign popcount47_atj4_core_121 = popcount47_atj4_core_111 ^ popcount47_atj4_core_117;
  assign popcount47_atj4_core_122 = popcount47_atj4_core_111 & popcount47_atj4_core_117;
  assign popcount47_atj4_core_123 = popcount47_atj4_core_121 ^ popcount47_atj4_core_120;
  assign popcount47_atj4_core_124 = popcount47_atj4_core_121 & popcount47_atj4_core_120;
  assign popcount47_atj4_core_125 = popcount47_atj4_core_122 | popcount47_atj4_core_124;
  assign popcount47_atj4_core_127 = input_a[20] & popcount47_atj4_core_118;
  assign popcount47_atj4_core_128 = popcount47_atj4_core_112 | popcount47_atj4_core_125;
  assign popcount47_atj4_core_131 = ~(input_a[19] & input_a[19]);
  assign popcount47_atj4_core_132 = input_a[3] & input_a[20];
  assign popcount47_atj4_core_133 = ~(input_a[14] & input_a[27]);
  assign popcount47_atj4_core_137 = input_a[21] ^ input_a[22];
  assign popcount47_atj4_core_140 = input_a[44] & input_a[18];
  assign popcount47_atj4_core_144 = popcount47_atj4_core_133 & input_a[26];
  assign popcount47_atj4_core_146 = popcount47_atj4_core_132 & popcount47_atj4_core_140;
  assign popcount47_atj4_core_155 = input_a[31] ^ input_a[6];
  assign popcount47_atj4_core_156 = popcount47_atj4_core_119 & input_a[6];
  assign popcount47_atj4_core_159 = popcount47_atj4_core_123 ^ popcount47_atj4_core_156;
  assign popcount47_atj4_core_160 = popcount47_atj4_core_123 & popcount47_atj4_core_156;
  assign popcount47_atj4_core_162 = popcount47_atj4_core_128 ^ popcount47_atj4_core_146;
  assign popcount47_atj4_core_163 = popcount47_atj4_core_128 & popcount47_atj4_core_146;
  assign popcount47_atj4_core_164 = popcount47_atj4_core_162 ^ popcount47_atj4_core_160;
  assign popcount47_atj4_core_165 = popcount47_atj4_core_162 & popcount47_atj4_core_160;
  assign popcount47_atj4_core_166 = popcount47_atj4_core_163 | popcount47_atj4_core_165;
  assign popcount47_atj4_core_172 = input_a[27] ^ popcount47_atj4_core_155;
  assign popcount47_atj4_core_173 = input_a[17] & input_a[18];
  assign popcount47_atj4_core_174 = popcount47_atj4_core_092 ^ popcount47_atj4_core_159;
  assign popcount47_atj4_core_175 = popcount47_atj4_core_092 & popcount47_atj4_core_159;
  assign popcount47_atj4_core_176 = popcount47_atj4_core_174 ^ popcount47_atj4_core_173;
  assign popcount47_atj4_core_177 = popcount47_atj4_core_174 & popcount47_atj4_core_173;
  assign popcount47_atj4_core_178 = popcount47_atj4_core_175 | popcount47_atj4_core_177;
  assign popcount47_atj4_core_179 = popcount47_atj4_core_099 ^ popcount47_atj4_core_164;
  assign popcount47_atj4_core_180 = popcount47_atj4_core_099 & popcount47_atj4_core_164;
  assign popcount47_atj4_core_181 = popcount47_atj4_core_179 ^ popcount47_atj4_core_178;
  assign popcount47_atj4_core_182 = popcount47_atj4_core_179 & popcount47_atj4_core_178;
  assign popcount47_atj4_core_183 = popcount47_atj4_core_180 | popcount47_atj4_core_182;
  assign popcount47_atj4_core_184 = popcount47_atj4_core_104 ^ popcount47_atj4_core_166;
  assign popcount47_atj4_core_185 = popcount47_atj4_core_104 & popcount47_atj4_core_166;
  assign popcount47_atj4_core_186 = popcount47_atj4_core_184 ^ popcount47_atj4_core_183;
  assign popcount47_atj4_core_187 = popcount47_atj4_core_184 & popcount47_atj4_core_183;
  assign popcount47_atj4_core_188 = popcount47_atj4_core_185 | popcount47_atj4_core_187;
  assign popcount47_atj4_core_191 = popcount47_atj4_core_105 ^ popcount47_atj4_core_188;
  assign popcount47_atj4_core_195 = input_a[24] & input_a[25];
  assign popcount47_atj4_core_200 = ~(input_a[27] & input_a[28]);
  assign popcount47_atj4_core_201 = input_a[27] & input_a[28];
  assign popcount47_atj4_core_203 = input_a[26] & popcount47_atj4_core_200;
  assign popcount47_atj4_core_205 = popcount47_atj4_core_201 & popcount47_atj4_core_203;
  assign popcount47_atj4_core_208_not = ~popcount47_atj4_core_195;
  assign popcount47_atj4_core_214 = input_a[20] & popcount47_atj4_core_205;
  assign popcount47_atj4_core_215 = popcount47_atj4_core_205 ^ popcount47_atj4_core_195;
  assign popcount47_atj4_core_218 = input_a[30] ^ input_a[31];
  assign popcount47_atj4_core_219 = input_a[30] & input_a[31];
  assign popcount47_atj4_core_220 = input_a[29] ^ popcount47_atj4_core_218;
  assign popcount47_atj4_core_221 = input_a[29] & popcount47_atj4_core_218;
  assign popcount47_atj4_core_222 = popcount47_atj4_core_219 ^ popcount47_atj4_core_221;
  assign popcount47_atj4_core_224 = ~(input_a[2] & input_a[34]);
  assign popcount47_atj4_core_225 = ~(input_a[46] | input_a[34]);
  assign popcount47_atj4_core_226 = input_a[29] ^ input_a[34];
  assign popcount47_atj4_core_228 = input_a[21] ^ input_a[4];
  assign popcount47_atj4_core_230 = popcount47_atj4_core_220 & input_a[12];
  assign popcount47_atj4_core_231 = input_a[3] & popcount47_atj4_core_226;
  assign popcount47_atj4_core_232 = ~(popcount47_atj4_core_222 & popcount47_atj4_core_228);
  assign popcount47_atj4_core_233 = popcount47_atj4_core_222 & popcount47_atj4_core_228;
  assign popcount47_atj4_core_238 = input_a[35] & input_a[30];
  assign popcount47_atj4_core_242 = input_a[16] & input_a[42];
  assign popcount47_atj4_core_243 = input_a[23] & input_a[2];
  assign popcount47_atj4_core_244 = popcount47_atj4_core_208_not ^ popcount47_atj4_core_232;
  assign popcount47_atj4_core_245 = popcount47_atj4_core_208_not & popcount47_atj4_core_232;
  assign popcount47_atj4_core_246 = popcount47_atj4_core_244 ^ popcount47_atj4_core_243;
  assign popcount47_atj4_core_247 = input_a[43] & popcount47_atj4_core_243;
  assign popcount47_atj4_core_248 = popcount47_atj4_core_245 | popcount47_atj4_core_247;
  assign popcount47_atj4_core_249 = popcount47_atj4_core_215 ^ popcount47_atj4_core_233;
  assign popcount47_atj4_core_250 = popcount47_atj4_core_215 & popcount47_atj4_core_233;
  assign popcount47_atj4_core_251 = popcount47_atj4_core_249 ^ popcount47_atj4_core_248;
  assign popcount47_atj4_core_252 = popcount47_atj4_core_249 & popcount47_atj4_core_248;
  assign popcount47_atj4_core_253 = popcount47_atj4_core_250 | popcount47_atj4_core_252;
  assign popcount47_atj4_core_256 = popcount47_atj4_core_214 ^ popcount47_atj4_core_253;
  assign popcount47_atj4_core_257 = popcount47_atj4_core_214 & popcount47_atj4_core_253;
  assign popcount47_atj4_core_259 = input_a[36] ^ input_a[37];
  assign popcount47_atj4_core_260 = input_a[36] & input_a[37];
  assign popcount47_atj4_core_261 = input_a[35] ^ popcount47_atj4_core_259;
  assign popcount47_atj4_core_262 = input_a[35] & popcount47_atj4_core_259;
  assign popcount47_atj4_core_263 = popcount47_atj4_core_260 ^ popcount47_atj4_core_262;
  assign popcount47_atj4_core_264 = popcount47_atj4_core_260 & popcount47_atj4_core_262;
  assign popcount47_atj4_core_266 = input_a[39] & input_a[27];
  assign popcount47_atj4_core_267 = input_a[9] ^ input_a[4];
  assign popcount47_atj4_core_271 = popcount47_atj4_core_261 ^ popcount47_atj4_core_267;
  assign popcount47_atj4_core_272 = popcount47_atj4_core_261 & popcount47_atj4_core_267;
  assign popcount47_atj4_core_273 = popcount47_atj4_core_263 ^ popcount47_atj4_core_266;
  assign popcount47_atj4_core_274 = popcount47_atj4_core_263 & popcount47_atj4_core_266;
  assign popcount47_atj4_core_275 = popcount47_atj4_core_273 ^ popcount47_atj4_core_272;
  assign popcount47_atj4_core_276 = popcount47_atj4_core_273 & popcount47_atj4_core_272;
  assign popcount47_atj4_core_277 = popcount47_atj4_core_274 | popcount47_atj4_core_276;
  assign popcount47_atj4_core_280 = popcount47_atj4_core_264 ^ popcount47_atj4_core_277;
  assign popcount47_atj4_core_281 = popcount47_atj4_core_264 & popcount47_atj4_core_277;
  assign popcount47_atj4_core_283 = input_a[42] ^ input_a[43];
  assign popcount47_atj4_core_284 = input_a[26] & input_a[43];
  assign popcount47_atj4_core_285 = ~(input_a[24] & input_a[11]);
  assign popcount47_atj4_core_286 = input_a[28] & popcount47_atj4_core_283;
  assign popcount47_atj4_core_287 = popcount47_atj4_core_284 ^ popcount47_atj4_core_286;
  assign popcount47_atj4_core_290 = input_a[33] & input_a[46];
  assign popcount47_atj4_core_291 = input_a[44] ^ input_a[45];
  assign popcount47_atj4_core_292 = input_a[44] & input_a[45];
  assign popcount47_atj4_core_293 = popcount47_atj4_core_290 ^ popcount47_atj4_core_292;
  assign popcount47_atj4_core_294 = popcount47_atj4_core_290 & popcount47_atj4_core_292;
  assign popcount47_atj4_core_296 = input_a[4] & popcount47_atj4_core_291;
  assign popcount47_atj4_core_297 = popcount47_atj4_core_287 ^ popcount47_atj4_core_293;
  assign popcount47_atj4_core_298 = popcount47_atj4_core_287 & popcount47_atj4_core_293;
  assign popcount47_atj4_core_299 = popcount47_atj4_core_297 ^ popcount47_atj4_core_296;
  assign popcount47_atj4_core_300 = popcount47_atj4_core_297 & popcount47_atj4_core_296;
  assign popcount47_atj4_core_301 = popcount47_atj4_core_298 | popcount47_atj4_core_300;
  assign popcount47_atj4_core_304 = popcount47_atj4_core_294 ^ popcount47_atj4_core_301;
  assign popcount47_atj4_core_309 = popcount47_atj4_core_275 ^ popcount47_atj4_core_299;
  assign popcount47_atj4_core_310 = popcount47_atj4_core_275 & popcount47_atj4_core_299;
  assign popcount47_atj4_core_311 = popcount47_atj4_core_309 ^ popcount47_atj4_core_271;
  assign popcount47_atj4_core_312 = popcount47_atj4_core_309 & popcount47_atj4_core_271;
  assign popcount47_atj4_core_313 = popcount47_atj4_core_310 | popcount47_atj4_core_312;
  assign popcount47_atj4_core_314 = popcount47_atj4_core_280 ^ popcount47_atj4_core_304;
  assign popcount47_atj4_core_315 = popcount47_atj4_core_280 & popcount47_atj4_core_304;
  assign popcount47_atj4_core_316 = popcount47_atj4_core_314 ^ popcount47_atj4_core_313;
  assign popcount47_atj4_core_317 = popcount47_atj4_core_314 & popcount47_atj4_core_313;
  assign popcount47_atj4_core_318 = popcount47_atj4_core_315 | popcount47_atj4_core_317;
  assign popcount47_atj4_core_321 = popcount47_atj4_core_281 ^ popcount47_atj4_core_318;
  assign popcount47_atj4_core_322 = popcount47_atj4_core_281 & input_a[25];
  assign popcount47_atj4_core_323 = input_a[25] ^ input_a[9];
  assign popcount47_atj4_core_326 = popcount47_atj4_core_246 ^ popcount47_atj4_core_311;
  assign popcount47_atj4_core_327 = popcount47_atj4_core_246 & popcount47_atj4_core_311;
  assign popcount47_atj4_core_328 = popcount47_atj4_core_326 ^ input_a[34];
  assign popcount47_atj4_core_329 = popcount47_atj4_core_326 & input_a[34];
  assign popcount47_atj4_core_330 = popcount47_atj4_core_327 | popcount47_atj4_core_329;
  assign popcount47_atj4_core_331 = popcount47_atj4_core_251 ^ popcount47_atj4_core_316;
  assign popcount47_atj4_core_332 = popcount47_atj4_core_251 & popcount47_atj4_core_316;
  assign popcount47_atj4_core_333 = popcount47_atj4_core_331 ^ popcount47_atj4_core_330;
  assign popcount47_atj4_core_334 = popcount47_atj4_core_331 & popcount47_atj4_core_330;
  assign popcount47_atj4_core_335 = popcount47_atj4_core_332 | popcount47_atj4_core_334;
  assign popcount47_atj4_core_336 = popcount47_atj4_core_256 ^ popcount47_atj4_core_321;
  assign popcount47_atj4_core_337 = popcount47_atj4_core_256 & popcount47_atj4_core_321;
  assign popcount47_atj4_core_338 = popcount47_atj4_core_336 ^ popcount47_atj4_core_335;
  assign popcount47_atj4_core_339 = popcount47_atj4_core_336 & popcount47_atj4_core_335;
  assign popcount47_atj4_core_340 = popcount47_atj4_core_337 | popcount47_atj4_core_339;
  assign popcount47_atj4_core_343 = popcount47_atj4_core_257 | popcount47_atj4_core_340;
  assign popcount47_atj4_core_344 = input_a[33] & popcount47_atj4_core_340;
  assign popcount47_atj4_core_347 = ~(input_a[0] & input_a[34]);
  assign popcount47_atj4_core_348 = popcount47_atj4_core_176 ^ popcount47_atj4_core_328;
  assign popcount47_atj4_core_349 = popcount47_atj4_core_176 & popcount47_atj4_core_328;
  assign popcount47_atj4_core_350 = popcount47_atj4_core_348 ^ popcount47_atj4_core_347;
  assign popcount47_atj4_core_351 = popcount47_atj4_core_348 & popcount47_atj4_core_347;
  assign popcount47_atj4_core_352 = popcount47_atj4_core_349 | popcount47_atj4_core_351;
  assign popcount47_atj4_core_353 = popcount47_atj4_core_181 ^ popcount47_atj4_core_333;
  assign popcount47_atj4_core_354 = popcount47_atj4_core_181 & popcount47_atj4_core_333;
  assign popcount47_atj4_core_355 = popcount47_atj4_core_353 ^ popcount47_atj4_core_352;
  assign popcount47_atj4_core_356 = popcount47_atj4_core_353 & popcount47_atj4_core_352;
  assign popcount47_atj4_core_357 = popcount47_atj4_core_354 | popcount47_atj4_core_356;
  assign popcount47_atj4_core_358 = popcount47_atj4_core_186 ^ popcount47_atj4_core_338;
  assign popcount47_atj4_core_359 = popcount47_atj4_core_186 & popcount47_atj4_core_338;
  assign popcount47_atj4_core_360 = popcount47_atj4_core_358 ^ popcount47_atj4_core_357;
  assign popcount47_atj4_core_361 = popcount47_atj4_core_358 & popcount47_atj4_core_357;
  assign popcount47_atj4_core_362 = popcount47_atj4_core_359 | popcount47_atj4_core_361;
  assign popcount47_atj4_core_363 = popcount47_atj4_core_191 ^ popcount47_atj4_core_343;
  assign popcount47_atj4_core_364 = popcount47_atj4_core_191 & popcount47_atj4_core_343;
  assign popcount47_atj4_core_365 = popcount47_atj4_core_363 ^ popcount47_atj4_core_362;
  assign popcount47_atj4_core_366 = popcount47_atj4_core_363 & popcount47_atj4_core_362;
  assign popcount47_atj4_core_367 = popcount47_atj4_core_364 | popcount47_atj4_core_366;
  assign popcount47_atj4_core_368 = popcount47_atj4_core_105 & input_a[32];
  assign popcount47_atj4_core_369 = input_a[42] ^ input_a[32];
  assign popcount47_atj4_core_370 = popcount47_atj4_core_368 ^ popcount47_atj4_core_367;
  assign popcount47_atj4_core_371 = input_a[7] ^ input_a[18];
  assign popcount47_atj4_core_372 = ~(input_a[29] | input_a[1]);

  assign popcount47_atj4_out[0] = 1'b1;
  assign popcount47_atj4_out[1] = popcount47_atj4_core_350;
  assign popcount47_atj4_out[2] = popcount47_atj4_core_355;
  assign popcount47_atj4_out[3] = popcount47_atj4_core_360;
  assign popcount47_atj4_out[4] = popcount47_atj4_core_365;
  assign popcount47_atj4_out[5] = popcount47_atj4_core_370;
endmodule