// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.73629
// WCE=28.0
// EP=0.968996%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_62mx(input [27:0] input_a, output [4:0] popcount28_62mx_out);
  wire popcount28_62mx_core_030;
  wire popcount28_62mx_core_034;
  wire popcount28_62mx_core_035;
  wire popcount28_62mx_core_036;
  wire popcount28_62mx_core_038;
  wire popcount28_62mx_core_040;
  wire popcount28_62mx_core_041;
  wire popcount28_62mx_core_042;
  wire popcount28_62mx_core_043;
  wire popcount28_62mx_core_044_not;
  wire popcount28_62mx_core_048;
  wire popcount28_62mx_core_050;
  wire popcount28_62mx_core_053;
  wire popcount28_62mx_core_054;
  wire popcount28_62mx_core_055;
  wire popcount28_62mx_core_056;
  wire popcount28_62mx_core_058;
  wire popcount28_62mx_core_059;
  wire popcount28_62mx_core_060;
  wire popcount28_62mx_core_061;
  wire popcount28_62mx_core_062;
  wire popcount28_62mx_core_064;
  wire popcount28_62mx_core_065;
  wire popcount28_62mx_core_067;
  wire popcount28_62mx_core_068;
  wire popcount28_62mx_core_070;
  wire popcount28_62mx_core_073;
  wire popcount28_62mx_core_074;
  wire popcount28_62mx_core_076;
  wire popcount28_62mx_core_077;
  wire popcount28_62mx_core_078;
  wire popcount28_62mx_core_079;
  wire popcount28_62mx_core_080;
  wire popcount28_62mx_core_081;
  wire popcount28_62mx_core_083;
  wire popcount28_62mx_core_084;
  wire popcount28_62mx_core_085;
  wire popcount28_62mx_core_087;
  wire popcount28_62mx_core_088;
  wire popcount28_62mx_core_091;
  wire popcount28_62mx_core_093;
  wire popcount28_62mx_core_095;
  wire popcount28_62mx_core_096;
  wire popcount28_62mx_core_098;
  wire popcount28_62mx_core_101;
  wire popcount28_62mx_core_102;
  wire popcount28_62mx_core_103;
  wire popcount28_62mx_core_104;
  wire popcount28_62mx_core_106;
  wire popcount28_62mx_core_107;
  wire popcount28_62mx_core_112;
  wire popcount28_62mx_core_113;
  wire popcount28_62mx_core_114;
  wire popcount28_62mx_core_118;
  wire popcount28_62mx_core_119_not;
  wire popcount28_62mx_core_120;
  wire popcount28_62mx_core_124;
  wire popcount28_62mx_core_128;
  wire popcount28_62mx_core_129;
  wire popcount28_62mx_core_134;
  wire popcount28_62mx_core_136;
  wire popcount28_62mx_core_137;
  wire popcount28_62mx_core_138;
  wire popcount28_62mx_core_142;
  wire popcount28_62mx_core_143;
  wire popcount28_62mx_core_145;
  wire popcount28_62mx_core_146;
  wire popcount28_62mx_core_148;
  wire popcount28_62mx_core_150;
  wire popcount28_62mx_core_151;
  wire popcount28_62mx_core_152;
  wire popcount28_62mx_core_155;
  wire popcount28_62mx_core_158;
  wire popcount28_62mx_core_159;
  wire popcount28_62mx_core_160;
  wire popcount28_62mx_core_161;
  wire popcount28_62mx_core_163;
  wire popcount28_62mx_core_165;
  wire popcount28_62mx_core_166;
  wire popcount28_62mx_core_167;
  wire popcount28_62mx_core_170;
  wire popcount28_62mx_core_171;
  wire popcount28_62mx_core_173;
  wire popcount28_62mx_core_174;
  wire popcount28_62mx_core_176;
  wire popcount28_62mx_core_181;
  wire popcount28_62mx_core_182;
  wire popcount28_62mx_core_184;
  wire popcount28_62mx_core_185;
  wire popcount28_62mx_core_186;
  wire popcount28_62mx_core_188;
  wire popcount28_62mx_core_189;
  wire popcount28_62mx_core_190;
  wire popcount28_62mx_core_191;
  wire popcount28_62mx_core_192;
  wire popcount28_62mx_core_193;
  wire popcount28_62mx_core_195;
  wire popcount28_62mx_core_196;
  wire popcount28_62mx_core_197;
  wire popcount28_62mx_core_198;
  wire popcount28_62mx_core_199;
  wire popcount28_62mx_core_200;
  wire popcount28_62mx_core_201;

  assign popcount28_62mx_core_030 = ~(input_a[17] & input_a[11]);
  assign popcount28_62mx_core_034 = ~(input_a[27] | input_a[17]);
  assign popcount28_62mx_core_035 = input_a[13] & input_a[10];
  assign popcount28_62mx_core_036 = ~input_a[2];
  assign popcount28_62mx_core_038 = input_a[25] | input_a[8];
  assign popcount28_62mx_core_040 = input_a[9] | input_a[26];
  assign popcount28_62mx_core_041 = ~input_a[9];
  assign popcount28_62mx_core_042 = ~(input_a[2] | input_a[3]);
  assign popcount28_62mx_core_043 = ~(input_a[27] & input_a[8]);
  assign popcount28_62mx_core_044_not = ~input_a[21];
  assign popcount28_62mx_core_048 = ~input_a[20];
  assign popcount28_62mx_core_050 = input_a[22] & input_a[4];
  assign popcount28_62mx_core_053 = input_a[23] ^ input_a[27];
  assign popcount28_62mx_core_054 = input_a[27] & input_a[7];
  assign popcount28_62mx_core_055 = ~(input_a[0] ^ input_a[20]);
  assign popcount28_62mx_core_056 = ~(input_a[4] | input_a[22]);
  assign popcount28_62mx_core_058 = ~input_a[23];
  assign popcount28_62mx_core_059 = ~(input_a[10] ^ input_a[16]);
  assign popcount28_62mx_core_060 = ~(input_a[26] | input_a[19]);
  assign popcount28_62mx_core_061 = ~(input_a[27] & input_a[18]);
  assign popcount28_62mx_core_062 = input_a[2] | input_a[0];
  assign popcount28_62mx_core_064 = input_a[16] | input_a[0];
  assign popcount28_62mx_core_065 = ~(input_a[8] ^ input_a[2]);
  assign popcount28_62mx_core_067 = input_a[1] & input_a[11];
  assign popcount28_62mx_core_068 = input_a[11] & input_a[5];
  assign popcount28_62mx_core_070 = ~(input_a[10] & input_a[3]);
  assign popcount28_62mx_core_073 = ~(input_a[14] ^ input_a[12]);
  assign popcount28_62mx_core_074 = input_a[5] & input_a[25];
  assign popcount28_62mx_core_076 = ~input_a[17];
  assign popcount28_62mx_core_077 = ~(input_a[4] & input_a[4]);
  assign popcount28_62mx_core_078 = ~input_a[17];
  assign popcount28_62mx_core_079 = input_a[10] ^ input_a[1];
  assign popcount28_62mx_core_080 = input_a[6] ^ input_a[13];
  assign popcount28_62mx_core_081 = input_a[0] & input_a[22];
  assign popcount28_62mx_core_083 = ~input_a[2];
  assign popcount28_62mx_core_084 = ~(input_a[27] | input_a[21]);
  assign popcount28_62mx_core_085 = input_a[22] ^ input_a[8];
  assign popcount28_62mx_core_087 = input_a[24] ^ input_a[15];
  assign popcount28_62mx_core_088 = input_a[0] | input_a[21];
  assign popcount28_62mx_core_091 = input_a[3] & input_a[5];
  assign popcount28_62mx_core_093 = ~(input_a[20] | input_a[18]);
  assign popcount28_62mx_core_095 = ~(input_a[18] & input_a[20]);
  assign popcount28_62mx_core_096 = ~(input_a[17] | input_a[26]);
  assign popcount28_62mx_core_098 = input_a[27] | input_a[17];
  assign popcount28_62mx_core_101 = input_a[6] ^ input_a[17];
  assign popcount28_62mx_core_102 = input_a[0] | input_a[23];
  assign popcount28_62mx_core_103 = ~(input_a[18] & input_a[26]);
  assign popcount28_62mx_core_104 = input_a[10] ^ input_a[4];
  assign popcount28_62mx_core_106 = ~(input_a[18] & input_a[0]);
  assign popcount28_62mx_core_107 = input_a[16] | input_a[15];
  assign popcount28_62mx_core_112 = ~(input_a[16] & input_a[9]);
  assign popcount28_62mx_core_113 = ~(input_a[8] ^ input_a[12]);
  assign popcount28_62mx_core_114 = ~input_a[26];
  assign popcount28_62mx_core_118 = ~input_a[5];
  assign popcount28_62mx_core_119_not = ~input_a[22];
  assign popcount28_62mx_core_120 = ~(input_a[0] | input_a[8]);
  assign popcount28_62mx_core_124 = ~(input_a[9] | input_a[9]);
  assign popcount28_62mx_core_128 = ~input_a[14];
  assign popcount28_62mx_core_129 = input_a[21] | input_a[25];
  assign popcount28_62mx_core_134 = ~(input_a[6] | input_a[18]);
  assign popcount28_62mx_core_136 = input_a[15] ^ input_a[9];
  assign popcount28_62mx_core_137 = ~input_a[15];
  assign popcount28_62mx_core_138 = ~(input_a[26] ^ input_a[18]);
  assign popcount28_62mx_core_142 = ~(input_a[0] | input_a[15]);
  assign popcount28_62mx_core_143 = input_a[17] ^ input_a[14];
  assign popcount28_62mx_core_145 = ~(input_a[9] & input_a[9]);
  assign popcount28_62mx_core_146 = input_a[14] & input_a[19];
  assign popcount28_62mx_core_148 = input_a[15] | input_a[26];
  assign popcount28_62mx_core_150 = ~(input_a[17] & input_a[19]);
  assign popcount28_62mx_core_151 = ~(input_a[11] | input_a[25]);
  assign popcount28_62mx_core_152 = ~(input_a[1] & input_a[8]);
  assign popcount28_62mx_core_155 = ~(input_a[7] ^ input_a[3]);
  assign popcount28_62mx_core_158 = ~(input_a[24] | input_a[10]);
  assign popcount28_62mx_core_159 = ~(input_a[8] | input_a[24]);
  assign popcount28_62mx_core_160 = ~(input_a[27] ^ input_a[25]);
  assign popcount28_62mx_core_161 = input_a[10] & input_a[11];
  assign popcount28_62mx_core_163 = input_a[6] & input_a[15];
  assign popcount28_62mx_core_165 = ~input_a[0];
  assign popcount28_62mx_core_166 = ~(input_a[20] | input_a[6]);
  assign popcount28_62mx_core_167 = input_a[8] ^ input_a[13];
  assign popcount28_62mx_core_170 = input_a[26] & input_a[17];
  assign popcount28_62mx_core_171 = input_a[11] & input_a[19];
  assign popcount28_62mx_core_173 = ~(input_a[27] | input_a[15]);
  assign popcount28_62mx_core_174 = ~(input_a[18] | input_a[6]);
  assign popcount28_62mx_core_176 = input_a[20] ^ input_a[3];
  assign popcount28_62mx_core_181 = ~(input_a[25] | input_a[16]);
  assign popcount28_62mx_core_182 = ~(input_a[11] & input_a[10]);
  assign popcount28_62mx_core_184 = input_a[3] & input_a[14];
  assign popcount28_62mx_core_185 = ~(input_a[14] ^ input_a[24]);
  assign popcount28_62mx_core_186 = ~(input_a[2] & input_a[26]);
  assign popcount28_62mx_core_188 = ~(input_a[24] | input_a[1]);
  assign popcount28_62mx_core_189 = ~(input_a[9] & input_a[8]);
  assign popcount28_62mx_core_190 = ~(input_a[20] | input_a[21]);
  assign popcount28_62mx_core_191 = ~(input_a[17] | input_a[9]);
  assign popcount28_62mx_core_192 = input_a[8] & input_a[21];
  assign popcount28_62mx_core_193 = input_a[26] ^ input_a[5];
  assign popcount28_62mx_core_195 = input_a[10] & input_a[12];
  assign popcount28_62mx_core_196 = ~(input_a[17] ^ input_a[2]);
  assign popcount28_62mx_core_197 = ~input_a[7];
  assign popcount28_62mx_core_198 = ~input_a[8];
  assign popcount28_62mx_core_199 = ~(input_a[11] | input_a[16]);
  assign popcount28_62mx_core_200 = input_a[26] | input_a[17];
  assign popcount28_62mx_core_201 = input_a[17] | input_a[10];

  assign popcount28_62mx_out[0] = 1'b0;
  assign popcount28_62mx_out[1] = 1'b0;
  assign popcount28_62mx_out[2] = input_a[9];
  assign popcount28_62mx_out[3] = input_a[24];
  assign popcount28_62mx_out[4] = input_a[8];
endmodule