// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.78253
// WCE=18.0
// EP=0.890235%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_mod1(input [31:0] input_a, output [5:0] popcount32_mod1_out);
  wire popcount32_mod1_core_035;
  wire popcount32_mod1_core_037;
  wire popcount32_mod1_core_038;
  wire popcount32_mod1_core_039;
  wire popcount32_mod1_core_041;
  wire popcount32_mod1_core_042;
  wire popcount32_mod1_core_043;
  wire popcount32_mod1_core_044;
  wire popcount32_mod1_core_045;
  wire popcount32_mod1_core_046;
  wire popcount32_mod1_core_047;
  wire popcount32_mod1_core_048;
  wire popcount32_mod1_core_050;
  wire popcount32_mod1_core_051;
  wire popcount32_mod1_core_053;
  wire popcount32_mod1_core_054;
  wire popcount32_mod1_core_055;
  wire popcount32_mod1_core_057;
  wire popcount32_mod1_core_058;
  wire popcount32_mod1_core_059;
  wire popcount32_mod1_core_060;
  wire popcount32_mod1_core_061;
  wire popcount32_mod1_core_062;
  wire popcount32_mod1_core_063;
  wire popcount32_mod1_core_066;
  wire popcount32_mod1_core_067;
  wire popcount32_mod1_core_069;
  wire popcount32_mod1_core_071;
  wire popcount32_mod1_core_074;
  wire popcount32_mod1_core_075;
  wire popcount32_mod1_core_076;
  wire popcount32_mod1_core_078;
  wire popcount32_mod1_core_080;
  wire popcount32_mod1_core_081;
  wire popcount32_mod1_core_082;
  wire popcount32_mod1_core_085;
  wire popcount32_mod1_core_086;
  wire popcount32_mod1_core_090;
  wire popcount32_mod1_core_091;
  wire popcount32_mod1_core_099;
  wire popcount32_mod1_core_100;
  wire popcount32_mod1_core_102;
  wire popcount32_mod1_core_103;
  wire popcount32_mod1_core_105;
  wire popcount32_mod1_core_107;
  wire popcount32_mod1_core_108;
  wire popcount32_mod1_core_109;
  wire popcount32_mod1_core_110;
  wire popcount32_mod1_core_112;
  wire popcount32_mod1_core_114;
  wire popcount32_mod1_core_115;
  wire popcount32_mod1_core_116;
  wire popcount32_mod1_core_118;
  wire popcount32_mod1_core_121;
  wire popcount32_mod1_core_124;
  wire popcount32_mod1_core_125;
  wire popcount32_mod1_core_127;
  wire popcount32_mod1_core_128;
  wire popcount32_mod1_core_131;
  wire popcount32_mod1_core_135_not;
  wire popcount32_mod1_core_138;
  wire popcount32_mod1_core_139;
  wire popcount32_mod1_core_140;
  wire popcount32_mod1_core_141;
  wire popcount32_mod1_core_142;
  wire popcount32_mod1_core_146;
  wire popcount32_mod1_core_147;
  wire popcount32_mod1_core_149;
  wire popcount32_mod1_core_150;
  wire popcount32_mod1_core_152;
  wire popcount32_mod1_core_154;
  wire popcount32_mod1_core_157;
  wire popcount32_mod1_core_158;
  wire popcount32_mod1_core_159;
  wire popcount32_mod1_core_160;
  wire popcount32_mod1_core_161;
  wire popcount32_mod1_core_163;
  wire popcount32_mod1_core_164;
  wire popcount32_mod1_core_166;
  wire popcount32_mod1_core_167;
  wire popcount32_mod1_core_170;
  wire popcount32_mod1_core_171;
  wire popcount32_mod1_core_173;
  wire popcount32_mod1_core_174;
  wire popcount32_mod1_core_177;
  wire popcount32_mod1_core_178;
  wire popcount32_mod1_core_179;
  wire popcount32_mod1_core_180;
  wire popcount32_mod1_core_181;
  wire popcount32_mod1_core_183;
  wire popcount32_mod1_core_184;
  wire popcount32_mod1_core_186;
  wire popcount32_mod1_core_187;
  wire popcount32_mod1_core_189;
  wire popcount32_mod1_core_192;
  wire popcount32_mod1_core_193;
  wire popcount32_mod1_core_194;
  wire popcount32_mod1_core_195;
  wire popcount32_mod1_core_196;
  wire popcount32_mod1_core_197;
  wire popcount32_mod1_core_199;
  wire popcount32_mod1_core_201;
  wire popcount32_mod1_core_202;
  wire popcount32_mod1_core_203;
  wire popcount32_mod1_core_204;
  wire popcount32_mod1_core_206;
  wire popcount32_mod1_core_210;
  wire popcount32_mod1_core_211;
  wire popcount32_mod1_core_214;
  wire popcount32_mod1_core_215;
  wire popcount32_mod1_core_217;
  wire popcount32_mod1_core_218;
  wire popcount32_mod1_core_219;
  wire popcount32_mod1_core_222;

  assign popcount32_mod1_core_035 = ~(input_a[12] & input_a[9]);
  assign popcount32_mod1_core_037 = ~(input_a[10] ^ input_a[9]);
  assign popcount32_mod1_core_038 = input_a[30] ^ input_a[24];
  assign popcount32_mod1_core_039 = ~(input_a[15] & input_a[20]);
  assign popcount32_mod1_core_041 = ~(input_a[3] | input_a[23]);
  assign popcount32_mod1_core_042 = ~input_a[7];
  assign popcount32_mod1_core_043 = ~input_a[6];
  assign popcount32_mod1_core_044 = ~(input_a[15] ^ input_a[2]);
  assign popcount32_mod1_core_045 = input_a[31] | input_a[28];
  assign popcount32_mod1_core_046 = ~(input_a[10] ^ input_a[4]);
  assign popcount32_mod1_core_047 = ~(input_a[29] & input_a[21]);
  assign popcount32_mod1_core_048 = ~(input_a[4] ^ input_a[0]);
  assign popcount32_mod1_core_050 = ~input_a[5];
  assign popcount32_mod1_core_051 = input_a[19] ^ input_a[2];
  assign popcount32_mod1_core_053 = input_a[27] | input_a[19];
  assign popcount32_mod1_core_054 = input_a[26] ^ input_a[24];
  assign popcount32_mod1_core_055 = ~input_a[26];
  assign popcount32_mod1_core_057 = ~(input_a[31] ^ input_a[30]);
  assign popcount32_mod1_core_058 = ~(input_a[23] & input_a[14]);
  assign popcount32_mod1_core_059 = ~input_a[18];
  assign popcount32_mod1_core_060 = ~(input_a[5] | input_a[0]);
  assign popcount32_mod1_core_061 = ~(input_a[31] | input_a[17]);
  assign popcount32_mod1_core_062 = ~(input_a[0] | input_a[17]);
  assign popcount32_mod1_core_063 = ~(input_a[0] | input_a[10]);
  assign popcount32_mod1_core_066 = input_a[13] & input_a[1];
  assign popcount32_mod1_core_067 = input_a[22] ^ input_a[16];
  assign popcount32_mod1_core_069 = ~input_a[20];
  assign popcount32_mod1_core_071 = ~input_a[9];
  assign popcount32_mod1_core_074 = ~(input_a[8] ^ input_a[3]);
  assign popcount32_mod1_core_075 = input_a[14] | input_a[5];
  assign popcount32_mod1_core_076 = ~(input_a[28] | input_a[22]);
  assign popcount32_mod1_core_078 = input_a[6] | input_a[24];
  assign popcount32_mod1_core_080 = ~(input_a[12] ^ input_a[23]);
  assign popcount32_mod1_core_081 = input_a[11] ^ input_a[27];
  assign popcount32_mod1_core_082 = ~(input_a[5] & input_a[15]);
  assign popcount32_mod1_core_085 = ~(input_a[20] | input_a[10]);
  assign popcount32_mod1_core_086 = ~(input_a[6] | input_a[25]);
  assign popcount32_mod1_core_090 = ~(input_a[14] & input_a[8]);
  assign popcount32_mod1_core_091 = ~(input_a[6] & input_a[10]);
  assign popcount32_mod1_core_099 = ~input_a[26];
  assign popcount32_mod1_core_100 = ~input_a[27];
  assign popcount32_mod1_core_102 = ~(input_a[25] ^ input_a[25]);
  assign popcount32_mod1_core_103 = ~(input_a[5] ^ input_a[21]);
  assign popcount32_mod1_core_105 = ~(input_a[6] | input_a[28]);
  assign popcount32_mod1_core_107 = ~input_a[0];
  assign popcount32_mod1_core_108 = input_a[31] ^ input_a[7];
  assign popcount32_mod1_core_109 = input_a[9] | input_a[27];
  assign popcount32_mod1_core_110 = input_a[22] & input_a[4];
  assign popcount32_mod1_core_112 = ~(input_a[4] ^ input_a[31]);
  assign popcount32_mod1_core_114 = input_a[1] & input_a[9];
  assign popcount32_mod1_core_115 = ~input_a[0];
  assign popcount32_mod1_core_116 = input_a[19] & input_a[28];
  assign popcount32_mod1_core_118 = input_a[31] & input_a[29];
  assign popcount32_mod1_core_121 = ~(input_a[12] ^ input_a[18]);
  assign popcount32_mod1_core_124 = input_a[12] | input_a[19];
  assign popcount32_mod1_core_125 = input_a[5] | input_a[12];
  assign popcount32_mod1_core_127 = ~input_a[4];
  assign popcount32_mod1_core_128 = ~(input_a[13] ^ input_a[29]);
  assign popcount32_mod1_core_131 = ~(input_a[23] | input_a[5]);
  assign popcount32_mod1_core_135_not = ~input_a[23];
  assign popcount32_mod1_core_138 = input_a[6] | input_a[17];
  assign popcount32_mod1_core_139 = input_a[28] & input_a[26];
  assign popcount32_mod1_core_140 = ~(input_a[13] & input_a[14]);
  assign popcount32_mod1_core_141 = ~(input_a[14] | input_a[30]);
  assign popcount32_mod1_core_142 = input_a[5] ^ input_a[25];
  assign popcount32_mod1_core_146 = ~(input_a[24] | input_a[21]);
  assign popcount32_mod1_core_147 = ~input_a[29];
  assign popcount32_mod1_core_149 = input_a[13] | input_a[13];
  assign popcount32_mod1_core_150 = ~(input_a[8] ^ input_a[6]);
  assign popcount32_mod1_core_152 = ~(input_a[4] ^ input_a[20]);
  assign popcount32_mod1_core_154 = ~(input_a[18] & input_a[11]);
  assign popcount32_mod1_core_157 = input_a[27] | input_a[17];
  assign popcount32_mod1_core_158 = input_a[7] ^ input_a[6];
  assign popcount32_mod1_core_159 = ~input_a[7];
  assign popcount32_mod1_core_160 = ~(input_a[29] ^ input_a[15]);
  assign popcount32_mod1_core_161 = ~(input_a[5] & input_a[11]);
  assign popcount32_mod1_core_163 = ~(input_a[21] ^ input_a[19]);
  assign popcount32_mod1_core_164 = ~(input_a[11] | input_a[8]);
  assign popcount32_mod1_core_166 = ~input_a[19];
  assign popcount32_mod1_core_167 = input_a[4] & input_a[14];
  assign popcount32_mod1_core_170 = input_a[9] | input_a[8];
  assign popcount32_mod1_core_171 = input_a[17] ^ input_a[12];
  assign popcount32_mod1_core_173 = ~(input_a[0] & input_a[23]);
  assign popcount32_mod1_core_174 = ~(input_a[26] | input_a[7]);
  assign popcount32_mod1_core_177 = input_a[24] | input_a[9];
  assign popcount32_mod1_core_178 = ~(input_a[18] | input_a[8]);
  assign popcount32_mod1_core_179 = ~input_a[13];
  assign popcount32_mod1_core_180 = ~(input_a[1] | input_a[13]);
  assign popcount32_mod1_core_181 = input_a[16] | input_a[31];
  assign popcount32_mod1_core_183 = input_a[25] | input_a[11];
  assign popcount32_mod1_core_184 = input_a[10] | input_a[14];
  assign popcount32_mod1_core_186 = input_a[3] | input_a[11];
  assign popcount32_mod1_core_187 = ~(input_a[3] | input_a[5]);
  assign popcount32_mod1_core_189 = ~(input_a[11] ^ input_a[15]);
  assign popcount32_mod1_core_192 = input_a[13] | input_a[7];
  assign popcount32_mod1_core_193 = input_a[10] & input_a[20];
  assign popcount32_mod1_core_194 = input_a[21] ^ input_a[27];
  assign popcount32_mod1_core_195 = input_a[23] | input_a[13];
  assign popcount32_mod1_core_196 = input_a[18] | input_a[23];
  assign popcount32_mod1_core_197 = input_a[1] ^ input_a[9];
  assign popcount32_mod1_core_199 = ~(input_a[13] & input_a[14]);
  assign popcount32_mod1_core_201 = input_a[11] ^ input_a[12];
  assign popcount32_mod1_core_202 = ~(input_a[13] | input_a[0]);
  assign popcount32_mod1_core_203 = input_a[7] | input_a[16];
  assign popcount32_mod1_core_204 = ~(input_a[15] & input_a[10]);
  assign popcount32_mod1_core_206 = ~(input_a[20] ^ input_a[26]);
  assign popcount32_mod1_core_210 = input_a[11] | input_a[14];
  assign popcount32_mod1_core_211 = input_a[4] | input_a[14];
  assign popcount32_mod1_core_214 = ~input_a[9];
  assign popcount32_mod1_core_215 = ~input_a[25];
  assign popcount32_mod1_core_217 = input_a[31] & input_a[19];
  assign popcount32_mod1_core_218 = input_a[6] & input_a[13];
  assign popcount32_mod1_core_219 = input_a[9] & input_a[24];
  assign popcount32_mod1_core_222 = ~(input_a[20] ^ input_a[31]);

  assign popcount32_mod1_out[0] = 1'b1;
  assign popcount32_mod1_out[1] = input_a[10];
  assign popcount32_mod1_out[2] = 1'b1;
  assign popcount32_mod1_out[3] = 1'b1;
  assign popcount32_mod1_out[4] = 1'b0;
  assign popcount32_mod1_out[5] = 1'b0;
endmodule