// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.12993
// WCE=23.0
// EP=0.901238%
// Printed PDK parameters:
//  Area=3015890.0
//  Delay=9540127.0
//  Power=161710.0

module popcount45_dtro(input [44:0] input_a, output [5:0] popcount45_dtro_out);
  wire popcount45_dtro_core_047_not;
  wire popcount45_dtro_core_048;
  wire popcount45_dtro_core_049;
  wire popcount45_dtro_core_050_not;
  wire popcount45_dtro_core_051;
  wire popcount45_dtro_core_053;
  wire popcount45_dtro_core_056;
  wire popcount45_dtro_core_058;
  wire popcount45_dtro_core_060;
  wire popcount45_dtro_core_061;
  wire popcount45_dtro_core_062;
  wire popcount45_dtro_core_065;
  wire popcount45_dtro_core_066;
  wire popcount45_dtro_core_067;
  wire popcount45_dtro_core_068;
  wire popcount45_dtro_core_069;
  wire popcount45_dtro_core_070;
  wire popcount45_dtro_core_071;
  wire popcount45_dtro_core_073;
  wire popcount45_dtro_core_074;
  wire popcount45_dtro_core_075;
  wire popcount45_dtro_core_078;
  wire popcount45_dtro_core_079;
  wire popcount45_dtro_core_082;
  wire popcount45_dtro_core_083;
  wire popcount45_dtro_core_084;
  wire popcount45_dtro_core_085;
  wire popcount45_dtro_core_086;
  wire popcount45_dtro_core_087;
  wire popcount45_dtro_core_088;
  wire popcount45_dtro_core_089;
  wire popcount45_dtro_core_091;
  wire popcount45_dtro_core_092;
  wire popcount45_dtro_core_095;
  wire popcount45_dtro_core_097;
  wire popcount45_dtro_core_099;
  wire popcount45_dtro_core_100;
  wire popcount45_dtro_core_101;
  wire popcount45_dtro_core_103;
  wire popcount45_dtro_core_104;
  wire popcount45_dtro_core_106_not;
  wire popcount45_dtro_core_107_not;
  wire popcount45_dtro_core_110;
  wire popcount45_dtro_core_113;
  wire popcount45_dtro_core_114;
  wire popcount45_dtro_core_117;
  wire popcount45_dtro_core_118;
  wire popcount45_dtro_core_119;
  wire popcount45_dtro_core_121;
  wire popcount45_dtro_core_122;
  wire popcount45_dtro_core_123;
  wire popcount45_dtro_core_124;
  wire popcount45_dtro_core_125;
  wire popcount45_dtro_core_126;
  wire popcount45_dtro_core_127;
  wire popcount45_dtro_core_129;
  wire popcount45_dtro_core_130;
  wire popcount45_dtro_core_131;
  wire popcount45_dtro_core_132;
  wire popcount45_dtro_core_133;
  wire popcount45_dtro_core_137;
  wire popcount45_dtro_core_138;
  wire popcount45_dtro_core_139;
  wire popcount45_dtro_core_140;
  wire popcount45_dtro_core_141;
  wire popcount45_dtro_core_143;
  wire popcount45_dtro_core_145;
  wire popcount45_dtro_core_146;
  wire popcount45_dtro_core_147;
  wire popcount45_dtro_core_148;
  wire popcount45_dtro_core_149;
  wire popcount45_dtro_core_150;
  wire popcount45_dtro_core_151;
  wire popcount45_dtro_core_152;
  wire popcount45_dtro_core_153;
  wire popcount45_dtro_core_155;
  wire popcount45_dtro_core_156;
  wire popcount45_dtro_core_157;
  wire popcount45_dtro_core_159;
  wire popcount45_dtro_core_160;
  wire popcount45_dtro_core_162;
  wire popcount45_dtro_core_164;
  wire popcount45_dtro_core_166;
  wire popcount45_dtro_core_167;
  wire popcount45_dtro_core_169;
  wire popcount45_dtro_core_170;
  wire popcount45_dtro_core_171;
  wire popcount45_dtro_core_173;
  wire popcount45_dtro_core_175;
  wire popcount45_dtro_core_176;
  wire popcount45_dtro_core_178;
  wire popcount45_dtro_core_179;
  wire popcount45_dtro_core_180;
  wire popcount45_dtro_core_182;
  wire popcount45_dtro_core_185;
  wire popcount45_dtro_core_186;
  wire popcount45_dtro_core_187;
  wire popcount45_dtro_core_188;
  wire popcount45_dtro_core_189;
  wire popcount45_dtro_core_192;
  wire popcount45_dtro_core_193;
  wire popcount45_dtro_core_196;
  wire popcount45_dtro_core_197;
  wire popcount45_dtro_core_198;
  wire popcount45_dtro_core_203;
  wire popcount45_dtro_core_204;
  wire popcount45_dtro_core_205;
  wire popcount45_dtro_core_206;
  wire popcount45_dtro_core_208;
  wire popcount45_dtro_core_209;
  wire popcount45_dtro_core_210;
  wire popcount45_dtro_core_211;
  wire popcount45_dtro_core_212;
  wire popcount45_dtro_core_213;
  wire popcount45_dtro_core_214;
  wire popcount45_dtro_core_215;
  wire popcount45_dtro_core_216;
  wire popcount45_dtro_core_219;
  wire popcount45_dtro_core_220;
  wire popcount45_dtro_core_221;
  wire popcount45_dtro_core_222;
  wire popcount45_dtro_core_223;
  wire popcount45_dtro_core_224;
  wire popcount45_dtro_core_225;
  wire popcount45_dtro_core_226;
  wire popcount45_dtro_core_227;
  wire popcount45_dtro_core_228;
  wire popcount45_dtro_core_231;
  wire popcount45_dtro_core_232;
  wire popcount45_dtro_core_235;
  wire popcount45_dtro_core_236;
  wire popcount45_dtro_core_237;
  wire popcount45_dtro_core_238;
  wire popcount45_dtro_core_239;
  wire popcount45_dtro_core_240;
  wire popcount45_dtro_core_241;
  wire popcount45_dtro_core_242;
  wire popcount45_dtro_core_244;
  wire popcount45_dtro_core_247;
  wire popcount45_dtro_core_248;
  wire popcount45_dtro_core_250;
  wire popcount45_dtro_core_251;
  wire popcount45_dtro_core_254;
  wire popcount45_dtro_core_255;
  wire popcount45_dtro_core_256;
  wire popcount45_dtro_core_257;
  wire popcount45_dtro_core_258;
  wire popcount45_dtro_core_259;
  wire popcount45_dtro_core_260;
  wire popcount45_dtro_core_261;
  wire popcount45_dtro_core_262;
  wire popcount45_dtro_core_263;
  wire popcount45_dtro_core_264;
  wire popcount45_dtro_core_266;
  wire popcount45_dtro_core_267;
  wire popcount45_dtro_core_268;
  wire popcount45_dtro_core_269;
  wire popcount45_dtro_core_270;
  wire popcount45_dtro_core_272;
  wire popcount45_dtro_core_274;
  wire popcount45_dtro_core_275;
  wire popcount45_dtro_core_277;
  wire popcount45_dtro_core_278;
  wire popcount45_dtro_core_279;
  wire popcount45_dtro_core_280;
  wire popcount45_dtro_core_282;
  wire popcount45_dtro_core_283;
  wire popcount45_dtro_core_284;
  wire popcount45_dtro_core_287;
  wire popcount45_dtro_core_289;
  wire popcount45_dtro_core_290;
  wire popcount45_dtro_core_291;
  wire popcount45_dtro_core_292;
  wire popcount45_dtro_core_294;
  wire popcount45_dtro_core_295_not;
  wire popcount45_dtro_core_296;
  wire popcount45_dtro_core_297;
  wire popcount45_dtro_core_298;
  wire popcount45_dtro_core_301;
  wire popcount45_dtro_core_303;
  wire popcount45_dtro_core_305;
  wire popcount45_dtro_core_306;
  wire popcount45_dtro_core_307;
  wire popcount45_dtro_core_308;
  wire popcount45_dtro_core_310;
  wire popcount45_dtro_core_312;
  wire popcount45_dtro_core_314;
  wire popcount45_dtro_core_316;
  wire popcount45_dtro_core_317;
  wire popcount45_dtro_core_318;
  wire popcount45_dtro_core_321;
  wire popcount45_dtro_core_322;
  wire popcount45_dtro_core_326;
  wire popcount45_dtro_core_327;
  wire popcount45_dtro_core_329;
  wire popcount45_dtro_core_331;
  wire popcount45_dtro_core_333;
  wire popcount45_dtro_core_334;
  wire popcount45_dtro_core_336;
  wire popcount45_dtro_core_337_not;
  wire popcount45_dtro_core_340;
  wire popcount45_dtro_core_342_not;
  wire popcount45_dtro_core_343;
  wire popcount45_dtro_core_344;
  wire popcount45_dtro_core_345;
  wire popcount45_dtro_core_346;
  wire popcount45_dtro_core_347;
  wire popcount45_dtro_core_348;
  wire popcount45_dtro_core_349;
  wire popcount45_dtro_core_350;
  wire popcount45_dtro_core_352;
  wire popcount45_dtro_core_353;
  wire popcount45_dtro_core_354;
  wire popcount45_dtro_core_355;

  assign popcount45_dtro_core_047_not = ~input_a[12];
  assign popcount45_dtro_core_048 = input_a[34] | input_a[40];
  assign popcount45_dtro_core_049 = ~input_a[16];
  assign popcount45_dtro_core_050_not = ~input_a[6];
  assign popcount45_dtro_core_051 = input_a[30] & input_a[3];
  assign popcount45_dtro_core_053 = ~(input_a[34] | input_a[34]);
  assign popcount45_dtro_core_056 = ~(input_a[41] | input_a[18]);
  assign popcount45_dtro_core_058 = input_a[15] & input_a[31];
  assign popcount45_dtro_core_060 = ~(input_a[40] & input_a[11]);
  assign popcount45_dtro_core_061 = ~(input_a[5] ^ input_a[3]);
  assign popcount45_dtro_core_062 = input_a[36] | input_a[29];
  assign popcount45_dtro_core_065 = ~(input_a[33] | input_a[41]);
  assign popcount45_dtro_core_066 = input_a[25] ^ input_a[29];
  assign popcount45_dtro_core_067 = ~(input_a[23] | input_a[23]);
  assign popcount45_dtro_core_068 = ~(input_a[25] ^ input_a[42]);
  assign popcount45_dtro_core_069 = ~input_a[44];
  assign popcount45_dtro_core_070 = input_a[35] ^ input_a[32];
  assign popcount45_dtro_core_071 = ~(input_a[17] | input_a[35]);
  assign popcount45_dtro_core_073 = ~(input_a[44] & input_a[18]);
  assign popcount45_dtro_core_074 = input_a[42] | input_a[22];
  assign popcount45_dtro_core_075 = input_a[32] | input_a[21];
  assign popcount45_dtro_core_078 = input_a[13] & input_a[21];
  assign popcount45_dtro_core_079 = input_a[37] & input_a[34];
  assign popcount45_dtro_core_082 = input_a[37] ^ input_a[20];
  assign popcount45_dtro_core_083 = ~(input_a[27] & input_a[37]);
  assign popcount45_dtro_core_084 = ~input_a[33];
  assign popcount45_dtro_core_085 = ~(input_a[3] & input_a[1]);
  assign popcount45_dtro_core_086 = ~(input_a[8] & input_a[35]);
  assign popcount45_dtro_core_087 = input_a[20] | input_a[20];
  assign popcount45_dtro_core_088 = input_a[10] & input_a[33];
  assign popcount45_dtro_core_089 = ~(input_a[36] & input_a[30]);
  assign popcount45_dtro_core_091 = ~(input_a[31] | input_a[28]);
  assign popcount45_dtro_core_092 = input_a[13] | input_a[15];
  assign popcount45_dtro_core_095 = ~(input_a[20] & input_a[17]);
  assign popcount45_dtro_core_097 = input_a[9] ^ input_a[38];
  assign popcount45_dtro_core_099 = ~input_a[6];
  assign popcount45_dtro_core_100 = input_a[18] ^ input_a[19];
  assign popcount45_dtro_core_101 = ~(input_a[33] & input_a[20]);
  assign popcount45_dtro_core_103 = input_a[24] ^ input_a[2];
  assign popcount45_dtro_core_104 = ~(input_a[14] & input_a[13]);
  assign popcount45_dtro_core_106_not = ~input_a[25];
  assign popcount45_dtro_core_107_not = ~input_a[32];
  assign popcount45_dtro_core_110 = input_a[25] & input_a[29];
  assign popcount45_dtro_core_113 = input_a[35] | input_a[15];
  assign popcount45_dtro_core_114 = input_a[12] & input_a[18];
  assign popcount45_dtro_core_117 = ~(input_a[12] | input_a[25]);
  assign popcount45_dtro_core_118 = input_a[12] ^ input_a[34];
  assign popcount45_dtro_core_119 = ~(input_a[2] & input_a[7]);
  assign popcount45_dtro_core_121 = ~input_a[23];
  assign popcount45_dtro_core_122 = ~input_a[12];
  assign popcount45_dtro_core_123 = ~(input_a[35] & input_a[15]);
  assign popcount45_dtro_core_124 = ~(input_a[14] & input_a[15]);
  assign popcount45_dtro_core_125 = input_a[41] | input_a[1];
  assign popcount45_dtro_core_126 = ~(input_a[35] | input_a[31]);
  assign popcount45_dtro_core_127 = input_a[3] & input_a[44];
  assign popcount45_dtro_core_129 = ~(input_a[17] ^ input_a[22]);
  assign popcount45_dtro_core_130 = input_a[10] | input_a[34];
  assign popcount45_dtro_core_131 = ~(input_a[22] & input_a[21]);
  assign popcount45_dtro_core_132 = ~(input_a[35] | input_a[10]);
  assign popcount45_dtro_core_133 = ~(input_a[42] & input_a[38]);
  assign popcount45_dtro_core_137 = ~(input_a[38] | input_a[29]);
  assign popcount45_dtro_core_138 = ~(input_a[37] ^ input_a[43]);
  assign popcount45_dtro_core_139 = ~(input_a[27] & input_a[13]);
  assign popcount45_dtro_core_140 = input_a[12] ^ input_a[30];
  assign popcount45_dtro_core_141 = ~(input_a[8] & input_a[17]);
  assign popcount45_dtro_core_143 = input_a[32] | input_a[34];
  assign popcount45_dtro_core_145 = ~(input_a[31] ^ input_a[33]);
  assign popcount45_dtro_core_146 = input_a[13] ^ input_a[4];
  assign popcount45_dtro_core_147 = input_a[4] | input_a[21];
  assign popcount45_dtro_core_148 = input_a[29] | input_a[1];
  assign popcount45_dtro_core_149 = ~input_a[9];
  assign popcount45_dtro_core_150 = ~input_a[43];
  assign popcount45_dtro_core_151 = ~(input_a[36] | input_a[19]);
  assign popcount45_dtro_core_152 = input_a[7] & input_a[30];
  assign popcount45_dtro_core_153 = ~(input_a[19] | input_a[42]);
  assign popcount45_dtro_core_155 = input_a[39] & input_a[3];
  assign popcount45_dtro_core_156 = input_a[25] | input_a[34];
  assign popcount45_dtro_core_157 = input_a[28] & input_a[28];
  assign popcount45_dtro_core_159 = ~(input_a[22] | input_a[37]);
  assign popcount45_dtro_core_160 = ~input_a[41];
  assign popcount45_dtro_core_162 = ~input_a[33];
  assign popcount45_dtro_core_164 = ~(input_a[28] ^ input_a[27]);
  assign popcount45_dtro_core_166 = input_a[20] | input_a[24];
  assign popcount45_dtro_core_167 = ~input_a[28];
  assign popcount45_dtro_core_169 = input_a[32] | input_a[6];
  assign popcount45_dtro_core_170 = input_a[12] | input_a[14];
  assign popcount45_dtro_core_171 = input_a[35] ^ input_a[44];
  assign popcount45_dtro_core_173 = input_a[43] | input_a[30];
  assign popcount45_dtro_core_175 = input_a[12] ^ input_a[16];
  assign popcount45_dtro_core_176 = ~(input_a[17] ^ input_a[13]);
  assign popcount45_dtro_core_178 = ~(input_a[7] & input_a[0]);
  assign popcount45_dtro_core_179 = ~(input_a[39] | input_a[37]);
  assign popcount45_dtro_core_180 = input_a[1] | input_a[11];
  assign popcount45_dtro_core_182 = ~(input_a[36] & input_a[0]);
  assign popcount45_dtro_core_185 = input_a[22] & input_a[35];
  assign popcount45_dtro_core_186 = input_a[3] | input_a[17];
  assign popcount45_dtro_core_187 = ~(input_a[11] | input_a[44]);
  assign popcount45_dtro_core_188 = ~(input_a[12] | input_a[9]);
  assign popcount45_dtro_core_189 = ~input_a[41];
  assign popcount45_dtro_core_192 = ~(input_a[2] ^ input_a[17]);
  assign popcount45_dtro_core_193 = ~(input_a[20] | input_a[2]);
  assign popcount45_dtro_core_196 = ~(input_a[39] ^ input_a[2]);
  assign popcount45_dtro_core_197 = ~(input_a[9] & input_a[1]);
  assign popcount45_dtro_core_198 = ~(input_a[10] ^ input_a[8]);
  assign popcount45_dtro_core_203 = input_a[14] | input_a[25];
  assign popcount45_dtro_core_204 = ~(input_a[1] | input_a[41]);
  assign popcount45_dtro_core_205 = input_a[1] & input_a[37];
  assign popcount45_dtro_core_206 = input_a[38] ^ input_a[28];
  assign popcount45_dtro_core_208 = ~input_a[16];
  assign popcount45_dtro_core_209 = ~(input_a[32] | input_a[18]);
  assign popcount45_dtro_core_210 = ~(input_a[24] ^ input_a[39]);
  assign popcount45_dtro_core_211 = ~input_a[27];
  assign popcount45_dtro_core_212 = ~input_a[5];
  assign popcount45_dtro_core_213 = ~(input_a[33] & input_a[0]);
  assign popcount45_dtro_core_214 = ~input_a[14];
  assign popcount45_dtro_core_215 = ~(input_a[30] | input_a[18]);
  assign popcount45_dtro_core_216 = input_a[26] ^ input_a[31];
  assign popcount45_dtro_core_219 = ~input_a[25];
  assign popcount45_dtro_core_220 = ~(input_a[39] | input_a[18]);
  assign popcount45_dtro_core_221 = ~(input_a[0] & input_a[14]);
  assign popcount45_dtro_core_222 = ~input_a[32];
  assign popcount45_dtro_core_223 = ~(input_a[39] & input_a[16]);
  assign popcount45_dtro_core_224 = ~(input_a[5] | input_a[10]);
  assign popcount45_dtro_core_225 = input_a[12] ^ input_a[10];
  assign popcount45_dtro_core_226 = ~(input_a[39] | input_a[4]);
  assign popcount45_dtro_core_227 = ~(input_a[7] ^ input_a[31]);
  assign popcount45_dtro_core_228 = ~(input_a[44] | input_a[23]);
  assign popcount45_dtro_core_231 = input_a[26] & input_a[13];
  assign popcount45_dtro_core_232 = input_a[40] | input_a[3];
  assign popcount45_dtro_core_235 = ~(input_a[5] & popcount45_dtro_core_232);
  assign popcount45_dtro_core_236 = input_a[36] ^ input_a[4];
  assign popcount45_dtro_core_237 = input_a[3] | input_a[40];
  assign popcount45_dtro_core_238 = ~input_a[23];
  assign popcount45_dtro_core_239 = input_a[34] ^ input_a[27];
  assign popcount45_dtro_core_240 = input_a[32] | popcount45_dtro_core_237;
  assign popcount45_dtro_core_241 = ~(input_a[30] | input_a[38]);
  assign popcount45_dtro_core_242 = input_a[37] & input_a[6];
  assign popcount45_dtro_core_244 = ~(input_a[6] ^ input_a[14]);
  assign popcount45_dtro_core_247 = ~(input_a[38] ^ input_a[24]);
  assign popcount45_dtro_core_248 = input_a[41] | input_a[6];
  assign popcount45_dtro_core_250 = input_a[5] & input_a[6];
  assign popcount45_dtro_core_251 = ~(input_a[8] ^ input_a[28]);
  assign popcount45_dtro_core_254 = input_a[14] | input_a[27];
  assign popcount45_dtro_core_255 = ~(input_a[10] | input_a[38]);
  assign popcount45_dtro_core_256 = ~(input_a[30] & input_a[25]);
  assign popcount45_dtro_core_257 = ~(input_a[5] | input_a[20]);
  assign popcount45_dtro_core_258 = input_a[1] | input_a[41];
  assign popcount45_dtro_core_259 = input_a[1] & input_a[16];
  assign popcount45_dtro_core_260 = ~input_a[25];
  assign popcount45_dtro_core_261 = ~(input_a[43] ^ input_a[35]);
  assign popcount45_dtro_core_262 = input_a[12] | input_a[0];
  assign popcount45_dtro_core_263 = ~(input_a[41] ^ input_a[4]);
  assign popcount45_dtro_core_264 = input_a[16] ^ input_a[2];
  assign popcount45_dtro_core_266 = ~input_a[21];
  assign popcount45_dtro_core_267 = input_a[1] ^ input_a[29];
  assign popcount45_dtro_core_268 = input_a[4] | input_a[42];
  assign popcount45_dtro_core_269 = ~input_a[33];
  assign popcount45_dtro_core_270 = input_a[28] ^ input_a[33];
  assign popcount45_dtro_core_272 = ~(input_a[41] | input_a[26]);
  assign popcount45_dtro_core_274 = ~(input_a[32] ^ input_a[31]);
  assign popcount45_dtro_core_275 = ~(input_a[32] | input_a[7]);
  assign popcount45_dtro_core_277 = ~(input_a[5] ^ input_a[9]);
  assign popcount45_dtro_core_278 = input_a[25] ^ input_a[12];
  assign popcount45_dtro_core_279 = ~(input_a[34] | input_a[25]);
  assign popcount45_dtro_core_280 = input_a[29] & input_a[15];
  assign popcount45_dtro_core_282 = ~(input_a[35] | input_a[31]);
  assign popcount45_dtro_core_283 = ~(input_a[10] | input_a[32]);
  assign popcount45_dtro_core_284 = input_a[42] & input_a[14];
  assign popcount45_dtro_core_287 = input_a[32] | input_a[32];
  assign popcount45_dtro_core_289 = input_a[30] & input_a[25];
  assign popcount45_dtro_core_290 = ~(input_a[28] | input_a[36]);
  assign popcount45_dtro_core_291 = ~(input_a[22] & input_a[24]);
  assign popcount45_dtro_core_292 = ~input_a[7];
  assign popcount45_dtro_core_294 = input_a[42] | input_a[4];
  assign popcount45_dtro_core_295_not = ~input_a[36];
  assign popcount45_dtro_core_296 = ~(input_a[44] & input_a[1]);
  assign popcount45_dtro_core_297 = ~input_a[5];
  assign popcount45_dtro_core_298 = ~(input_a[7] ^ input_a[21]);
  assign popcount45_dtro_core_301 = ~(input_a[18] | input_a[24]);
  assign popcount45_dtro_core_303 = ~(input_a[28] & input_a[16]);
  assign popcount45_dtro_core_305 = input_a[14] & input_a[8];
  assign popcount45_dtro_core_306 = input_a[41] & input_a[5];
  assign popcount45_dtro_core_307 = ~(input_a[34] | input_a[15]);
  assign popcount45_dtro_core_308 = input_a[30] & input_a[4];
  assign popcount45_dtro_core_310 = ~input_a[26];
  assign popcount45_dtro_core_312 = input_a[0] | input_a[35];
  assign popcount45_dtro_core_314 = input_a[5] | input_a[27];
  assign popcount45_dtro_core_316 = input_a[19] & input_a[41];
  assign popcount45_dtro_core_317 = popcount45_dtro_core_235 ^ input_a[32];
  assign popcount45_dtro_core_318 = ~(input_a[4] | input_a[33]);
  assign popcount45_dtro_core_321 = ~(input_a[40] | input_a[14]);
  assign popcount45_dtro_core_322 = popcount45_dtro_core_240 | popcount45_dtro_core_316;
  assign popcount45_dtro_core_326 = ~input_a[29];
  assign popcount45_dtro_core_327 = input_a[14] ^ input_a[44];
  assign popcount45_dtro_core_329 = ~input_a[41];
  assign popcount45_dtro_core_331 = input_a[36] | input_a[27];
  assign popcount45_dtro_core_333 = input_a[40] ^ input_a[41];
  assign popcount45_dtro_core_334 = input_a[1] | input_a[16];
  assign popcount45_dtro_core_336 = ~(input_a[42] & input_a[18]);
  assign popcount45_dtro_core_337_not = ~popcount45_dtro_core_317;
  assign popcount45_dtro_core_340 = ~(input_a[37] | input_a[2]);
  assign popcount45_dtro_core_342_not = ~popcount45_dtro_core_322;
  assign popcount45_dtro_core_343 = ~(input_a[19] & input_a[20]);
  assign popcount45_dtro_core_344 = popcount45_dtro_core_342_not ^ popcount45_dtro_core_317;
  assign popcount45_dtro_core_345 = input_a[34] | input_a[8];
  assign popcount45_dtro_core_346 = input_a[11] | input_a[8];
  assign popcount45_dtro_core_347 = input_a[23] & input_a[24];
  assign popcount45_dtro_core_348 = ~(input_a[42] ^ input_a[44]);
  assign popcount45_dtro_core_349 = ~(input_a[21] & input_a[40]);
  assign popcount45_dtro_core_350 = ~input_a[40];
  assign popcount45_dtro_core_352 = input_a[27] | input_a[5];
  assign popcount45_dtro_core_353 = ~(input_a[27] | input_a[7]);
  assign popcount45_dtro_core_354 = input_a[25] | input_a[27];
  assign popcount45_dtro_core_355 = input_a[36] | input_a[8];

  assign popcount45_dtro_out[0] = input_a[1];
  assign popcount45_dtro_out[1] = input_a[5];
  assign popcount45_dtro_out[2] = popcount45_dtro_core_337_not;
  assign popcount45_dtro_out[3] = popcount45_dtro_core_344;
  assign popcount45_dtro_out[4] = 1'b1;
  assign popcount45_dtro_out[5] = 1'b0;
endmodule