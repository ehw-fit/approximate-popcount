// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.70669
// WCE=8.0
// EP=0.820683%
// Printed PDK parameters:
//  Area=64907251.0
//  Delay=96404064.0
//  Power=3264900.0

module popcount38_5cwm(input [37:0] input_a, output [5:0] popcount38_5cwm_out);
  wire popcount38_5cwm_core_040;
  wire popcount38_5cwm_core_041;
  wire popcount38_5cwm_core_042;
  wire popcount38_5cwm_core_043;
  wire popcount38_5cwm_core_044;
  wire popcount38_5cwm_core_045;
  wire popcount38_5cwm_core_046;
  wire popcount38_5cwm_core_047;
  wire popcount38_5cwm_core_048;
  wire popcount38_5cwm_core_051;
  wire popcount38_5cwm_core_052;
  wire popcount38_5cwm_core_053;
  wire popcount38_5cwm_core_054;
  wire popcount38_5cwm_core_055;
  wire popcount38_5cwm_core_060;
  wire popcount38_5cwm_core_061;
  wire popcount38_5cwm_core_063;
  wire popcount38_5cwm_core_064;
  wire popcount38_5cwm_core_066;
  wire popcount38_5cwm_core_067;
  wire popcount38_5cwm_core_068;
  wire popcount38_5cwm_core_069;
  wire popcount38_5cwm_core_070;
  wire popcount38_5cwm_core_071;
  wire popcount38_5cwm_core_073;
  wire popcount38_5cwm_core_076;
  wire popcount38_5cwm_core_077;
  wire popcount38_5cwm_core_078;
  wire popcount38_5cwm_core_079;
  wire popcount38_5cwm_core_083;
  wire popcount38_5cwm_core_085;
  wire popcount38_5cwm_core_089;
  wire popcount38_5cwm_core_090;
  wire popcount38_5cwm_core_092;
  wire popcount38_5cwm_core_095;
  wire popcount38_5cwm_core_098;
  wire popcount38_5cwm_core_099;
  wire popcount38_5cwm_core_100;
  wire popcount38_5cwm_core_101;
  wire popcount38_5cwm_core_102;
  wire popcount38_5cwm_core_104;
  wire popcount38_5cwm_core_105;
  wire popcount38_5cwm_core_107;
  wire popcount38_5cwm_core_108;
  wire popcount38_5cwm_core_109;
  wire popcount38_5cwm_core_110;
  wire popcount38_5cwm_core_111;
  wire popcount38_5cwm_core_112;
  wire popcount38_5cwm_core_113;
  wire popcount38_5cwm_core_115;
  wire popcount38_5cwm_core_116;
  wire popcount38_5cwm_core_117;
  wire popcount38_5cwm_core_119;
  wire popcount38_5cwm_core_124;
  wire popcount38_5cwm_core_125;
  wire popcount38_5cwm_core_128;
  wire popcount38_5cwm_core_129;
  wire popcount38_5cwm_core_131;
  wire popcount38_5cwm_core_132;
  wire popcount38_5cwm_core_133;
  wire popcount38_5cwm_core_136;
  wire popcount38_5cwm_core_138;
  wire popcount38_5cwm_core_139;
  wire popcount38_5cwm_core_140;
  wire popcount38_5cwm_core_142;
  wire popcount38_5cwm_core_144;
  wire popcount38_5cwm_core_146_not;
  wire popcount38_5cwm_core_149;
  wire popcount38_5cwm_core_150;
  wire popcount38_5cwm_core_151;
  wire popcount38_5cwm_core_153;
  wire popcount38_5cwm_core_154;
  wire popcount38_5cwm_core_155;
  wire popcount38_5cwm_core_156;
  wire popcount38_5cwm_core_157;
  wire popcount38_5cwm_core_158;
  wire popcount38_5cwm_core_159;
  wire popcount38_5cwm_core_161;
  wire popcount38_5cwm_core_162;
  wire popcount38_5cwm_core_163;
  wire popcount38_5cwm_core_164;
  wire popcount38_5cwm_core_166;
  wire popcount38_5cwm_core_167;
  wire popcount38_5cwm_core_169;
  wire popcount38_5cwm_core_170;
  wire popcount38_5cwm_core_171;
  wire popcount38_5cwm_core_176;
  wire popcount38_5cwm_core_177;
  wire popcount38_5cwm_core_179_not;
  wire popcount38_5cwm_core_184;
  wire popcount38_5cwm_core_185;
  wire popcount38_5cwm_core_186;
  wire popcount38_5cwm_core_188;
  wire popcount38_5cwm_core_190;
  wire popcount38_5cwm_core_191;
  wire popcount38_5cwm_core_192;
  wire popcount38_5cwm_core_193;
  wire popcount38_5cwm_core_196;
  wire popcount38_5cwm_core_197;
  wire popcount38_5cwm_core_198;
  wire popcount38_5cwm_core_199;
  wire popcount38_5cwm_core_200;
  wire popcount38_5cwm_core_201;
  wire popcount38_5cwm_core_202;
  wire popcount38_5cwm_core_203;
  wire popcount38_5cwm_core_205;
  wire popcount38_5cwm_core_206;
  wire popcount38_5cwm_core_207;
  wire popcount38_5cwm_core_208;
  wire popcount38_5cwm_core_209;
  wire popcount38_5cwm_core_210;
  wire popcount38_5cwm_core_211;
  wire popcount38_5cwm_core_213;
  wire popcount38_5cwm_core_214;
  wire popcount38_5cwm_core_215;
  wire popcount38_5cwm_core_217;
  wire popcount38_5cwm_core_218;
  wire popcount38_5cwm_core_219;
  wire popcount38_5cwm_core_220;
  wire popcount38_5cwm_core_222;
  wire popcount38_5cwm_core_224;
  wire popcount38_5cwm_core_225;
  wire popcount38_5cwm_core_226;
  wire popcount38_5cwm_core_227;
  wire popcount38_5cwm_core_228;
  wire popcount38_5cwm_core_231;
  wire popcount38_5cwm_core_232;
  wire popcount38_5cwm_core_233;
  wire popcount38_5cwm_core_234;
  wire popcount38_5cwm_core_235;
  wire popcount38_5cwm_core_236;
  wire popcount38_5cwm_core_237;
  wire popcount38_5cwm_core_238;
  wire popcount38_5cwm_core_239;
  wire popcount38_5cwm_core_240;
  wire popcount38_5cwm_core_241;
  wire popcount38_5cwm_core_242;
  wire popcount38_5cwm_core_244;
  wire popcount38_5cwm_core_246;
  wire popcount38_5cwm_core_248_not;
  wire popcount38_5cwm_core_250;
  wire popcount38_5cwm_core_251;
  wire popcount38_5cwm_core_252;
  wire popcount38_5cwm_core_253;
  wire popcount38_5cwm_core_254;
  wire popcount38_5cwm_core_255;
  wire popcount38_5cwm_core_256;
  wire popcount38_5cwm_core_257;
  wire popcount38_5cwm_core_258;
  wire popcount38_5cwm_core_259;
  wire popcount38_5cwm_core_260;
  wire popcount38_5cwm_core_261;
  wire popcount38_5cwm_core_262;
  wire popcount38_5cwm_core_263;
  wire popcount38_5cwm_core_264;
  wire popcount38_5cwm_core_266;
  wire popcount38_5cwm_core_268;
  wire popcount38_5cwm_core_269;
  wire popcount38_5cwm_core_270;
  wire popcount38_5cwm_core_271;
  wire popcount38_5cwm_core_272;
  wire popcount38_5cwm_core_273;
  wire popcount38_5cwm_core_274;
  wire popcount38_5cwm_core_275;
  wire popcount38_5cwm_core_276;
  wire popcount38_5cwm_core_277;
  wire popcount38_5cwm_core_278;
  wire popcount38_5cwm_core_279;
  wire popcount38_5cwm_core_280;
  wire popcount38_5cwm_core_281;
  wire popcount38_5cwm_core_282;
  wire popcount38_5cwm_core_283;
  wire popcount38_5cwm_core_284;
  wire popcount38_5cwm_core_285;
  wire popcount38_5cwm_core_286;
  wire popcount38_5cwm_core_288;
  wire popcount38_5cwm_core_289;
  wire popcount38_5cwm_core_290;
  wire popcount38_5cwm_core_291;
  wire popcount38_5cwm_core_292;
  wire popcount38_5cwm_core_294;
  wire popcount38_5cwm_core_295;
  wire popcount38_5cwm_core_296;

  assign popcount38_5cwm_core_040 = input_a[26] | input_a[3];
  assign popcount38_5cwm_core_041 = input_a[7] & input_a[27];
  assign popcount38_5cwm_core_042 = input_a[2] ^ input_a[3];
  assign popcount38_5cwm_core_043 = input_a[2] & input_a[3];
  assign popcount38_5cwm_core_044 = input_a[13] ^ input_a[21];
  assign popcount38_5cwm_core_045 = input_a[11] & popcount38_5cwm_core_042;
  assign popcount38_5cwm_core_046 = popcount38_5cwm_core_041 ^ popcount38_5cwm_core_043;
  assign popcount38_5cwm_core_047 = popcount38_5cwm_core_041 & popcount38_5cwm_core_043;
  assign popcount38_5cwm_core_048 = popcount38_5cwm_core_046 | popcount38_5cwm_core_045;
  assign popcount38_5cwm_core_051 = ~(input_a[4] | input_a[15]);
  assign popcount38_5cwm_core_052 = input_a[29] | input_a[28];
  assign popcount38_5cwm_core_053 = ~input_a[19];
  assign popcount38_5cwm_core_054 = ~(input_a[13] & input_a[27]);
  assign popcount38_5cwm_core_055 = ~input_a[17];
  assign popcount38_5cwm_core_060 = input_a[13] | input_a[29];
  assign popcount38_5cwm_core_061 = ~input_a[15];
  assign popcount38_5cwm_core_063 = input_a[24] | input_a[5];
  assign popcount38_5cwm_core_064 = ~(input_a[19] ^ input_a[10]);
  assign popcount38_5cwm_core_066 = ~(input_a[26] & input_a[25]);
  assign popcount38_5cwm_core_067 = input_a[0] | input_a[28];
  assign popcount38_5cwm_core_068 = input_a[28] | input_a[5];
  assign popcount38_5cwm_core_069 = input_a[12] | input_a[8];
  assign popcount38_5cwm_core_070 = popcount38_5cwm_core_048 ^ popcount38_5cwm_core_063;
  assign popcount38_5cwm_core_071 = popcount38_5cwm_core_048 & popcount38_5cwm_core_063;
  assign popcount38_5cwm_core_073 = ~input_a[20];
  assign popcount38_5cwm_core_076 = ~(input_a[7] & input_a[16]);
  assign popcount38_5cwm_core_077 = popcount38_5cwm_core_047 | popcount38_5cwm_core_071;
  assign popcount38_5cwm_core_078 = ~input_a[6];
  assign popcount38_5cwm_core_079 = input_a[29] ^ input_a[4];
  assign popcount38_5cwm_core_083 = input_a[6] & input_a[10];
  assign popcount38_5cwm_core_085 = input_a[9] & input_a[8];
  assign popcount38_5cwm_core_089 = input_a[28] & input_a[35];
  assign popcount38_5cwm_core_090 = ~(input_a[18] ^ input_a[7]);
  assign popcount38_5cwm_core_092 = popcount38_5cwm_core_083 | popcount38_5cwm_core_085;
  assign popcount38_5cwm_core_095 = input_a[8] & input_a[27];
  assign popcount38_5cwm_core_098 = ~(input_a[2] | input_a[36]);
  assign popcount38_5cwm_core_099 = input_a[9] & input_a[14];
  assign popcount38_5cwm_core_100 = input_a[14] & input_a[15];
  assign popcount38_5cwm_core_101 = ~(input_a[31] ^ input_a[3]);
  assign popcount38_5cwm_core_102 = input_a[17] & input_a[12];
  assign popcount38_5cwm_core_104 = input_a[16] & input_a[22];
  assign popcount38_5cwm_core_105 = popcount38_5cwm_core_102 | popcount38_5cwm_core_104;
  assign popcount38_5cwm_core_107 = input_a[36] | input_a[1];
  assign popcount38_5cwm_core_108 = input_a[13] & input_a[25];
  assign popcount38_5cwm_core_109 = popcount38_5cwm_core_100 | popcount38_5cwm_core_105;
  assign popcount38_5cwm_core_110 = popcount38_5cwm_core_100 & popcount38_5cwm_core_105;
  assign popcount38_5cwm_core_111 = popcount38_5cwm_core_109 | popcount38_5cwm_core_108;
  assign popcount38_5cwm_core_112 = popcount38_5cwm_core_109 & popcount38_5cwm_core_108;
  assign popcount38_5cwm_core_113 = popcount38_5cwm_core_110 | popcount38_5cwm_core_112;
  assign popcount38_5cwm_core_115 = ~(input_a[31] | input_a[15]);
  assign popcount38_5cwm_core_116 = input_a[3] ^ input_a[1];
  assign popcount38_5cwm_core_117 = ~input_a[12];
  assign popcount38_5cwm_core_119 = popcount38_5cwm_core_092 & popcount38_5cwm_core_111;
  assign popcount38_5cwm_core_124 = ~(input_a[3] & input_a[34]);
  assign popcount38_5cwm_core_125 = popcount38_5cwm_core_113 | popcount38_5cwm_core_119;
  assign popcount38_5cwm_core_128 = ~(input_a[10] & input_a[4]);
  assign popcount38_5cwm_core_129 = ~(input_a[35] | input_a[32]);
  assign popcount38_5cwm_core_131 = ~(input_a[27] ^ input_a[16]);
  assign popcount38_5cwm_core_132 = input_a[0] ^ input_a[37];
  assign popcount38_5cwm_core_133 = input_a[5] & input_a[33];
  assign popcount38_5cwm_core_136 = input_a[14] & input_a[34];
  assign popcount38_5cwm_core_138 = ~(input_a[15] | input_a[36]);
  assign popcount38_5cwm_core_139 = ~(input_a[9] | input_a[3]);
  assign popcount38_5cwm_core_140 = popcount38_5cwm_core_077 ^ popcount38_5cwm_core_125;
  assign popcount38_5cwm_core_142 = ~popcount38_5cwm_core_140;
  assign popcount38_5cwm_core_144 = popcount38_5cwm_core_077 | popcount38_5cwm_core_140;
  assign popcount38_5cwm_core_146_not = ~input_a[26];
  assign popcount38_5cwm_core_149 = input_a[10] & input_a[30];
  assign popcount38_5cwm_core_150 = ~input_a[18];
  assign popcount38_5cwm_core_151 = ~(input_a[12] & input_a[31]);
  assign popcount38_5cwm_core_153 = input_a[11] ^ input_a[1];
  assign popcount38_5cwm_core_154 = input_a[33] | input_a[18];
  assign popcount38_5cwm_core_155 = input_a[19] ^ input_a[20];
  assign popcount38_5cwm_core_156 = input_a[19] & input_a[20];
  assign popcount38_5cwm_core_157 = input_a[7] | input_a[22];
  assign popcount38_5cwm_core_158 = ~input_a[26];
  assign popcount38_5cwm_core_159 = ~(input_a[29] & input_a[6]);
  assign popcount38_5cwm_core_161 = input_a[20] ^ input_a[21];
  assign popcount38_5cwm_core_162 = popcount38_5cwm_core_156 & input_a[21];
  assign popcount38_5cwm_core_163 = popcount38_5cwm_core_161 | popcount38_5cwm_core_155;
  assign popcount38_5cwm_core_164 = input_a[18] | input_a[15];
  assign popcount38_5cwm_core_166 = ~(input_a[15] | input_a[5]);
  assign popcount38_5cwm_core_167 = input_a[18] & input_a[35];
  assign popcount38_5cwm_core_169 = input_a[26] & input_a[23];
  assign popcount38_5cwm_core_170 = ~(input_a[37] | input_a[21]);
  assign popcount38_5cwm_core_171 = ~input_a[12];
  assign popcount38_5cwm_core_176 = popcount38_5cwm_core_167 ^ popcount38_5cwm_core_169;
  assign popcount38_5cwm_core_177 = popcount38_5cwm_core_167 & popcount38_5cwm_core_169;
  assign popcount38_5cwm_core_179_not = ~input_a[0];
  assign popcount38_5cwm_core_184 = ~input_a[1];
  assign popcount38_5cwm_core_185 = popcount38_5cwm_core_163 ^ popcount38_5cwm_core_176;
  assign popcount38_5cwm_core_186 = popcount38_5cwm_core_163 & popcount38_5cwm_core_176;
  assign popcount38_5cwm_core_188 = input_a[2] & input_a[24];
  assign popcount38_5cwm_core_190 = popcount38_5cwm_core_162 ^ popcount38_5cwm_core_177;
  assign popcount38_5cwm_core_191 = popcount38_5cwm_core_162 & popcount38_5cwm_core_177;
  assign popcount38_5cwm_core_192 = popcount38_5cwm_core_190 | popcount38_5cwm_core_186;
  assign popcount38_5cwm_core_193 = ~(input_a[16] & input_a[28]);
  assign popcount38_5cwm_core_196 = ~(input_a[37] & input_a[6]);
  assign popcount38_5cwm_core_197 = input_a[28] ^ input_a[29];
  assign popcount38_5cwm_core_198 = input_a[28] & input_a[29];
  assign popcount38_5cwm_core_199 = input_a[31] ^ input_a[32];
  assign popcount38_5cwm_core_200 = input_a[31] & input_a[32];
  assign popcount38_5cwm_core_201 = input_a[30] ^ popcount38_5cwm_core_199;
  assign popcount38_5cwm_core_202 = input_a[30] & popcount38_5cwm_core_199;
  assign popcount38_5cwm_core_203 = popcount38_5cwm_core_200 | popcount38_5cwm_core_202;
  assign popcount38_5cwm_core_205 = popcount38_5cwm_core_197 ^ popcount38_5cwm_core_201;
  assign popcount38_5cwm_core_206 = popcount38_5cwm_core_197 & popcount38_5cwm_core_201;
  assign popcount38_5cwm_core_207 = popcount38_5cwm_core_198 ^ popcount38_5cwm_core_203;
  assign popcount38_5cwm_core_208 = popcount38_5cwm_core_198 & popcount38_5cwm_core_203;
  assign popcount38_5cwm_core_209 = popcount38_5cwm_core_207 ^ popcount38_5cwm_core_206;
  assign popcount38_5cwm_core_210 = popcount38_5cwm_core_207 & popcount38_5cwm_core_206;
  assign popcount38_5cwm_core_211 = popcount38_5cwm_core_208 | popcount38_5cwm_core_210;
  assign popcount38_5cwm_core_213 = input_a[13] | input_a[22];
  assign popcount38_5cwm_core_214 = input_a[33] ^ input_a[34];
  assign popcount38_5cwm_core_215 = input_a[33] & input_a[34];
  assign popcount38_5cwm_core_217 = input_a[36] & input_a[37];
  assign popcount38_5cwm_core_218 = ~(input_a[22] & input_a[24]);
  assign popcount38_5cwm_core_219 = input_a[1] & input_a[0];
  assign popcount38_5cwm_core_220 = popcount38_5cwm_core_217 | popcount38_5cwm_core_219;
  assign popcount38_5cwm_core_222 = ~popcount38_5cwm_core_214;
  assign popcount38_5cwm_core_224 = popcount38_5cwm_core_215 ^ popcount38_5cwm_core_220;
  assign popcount38_5cwm_core_225 = input_a[34] & popcount38_5cwm_core_220;
  assign popcount38_5cwm_core_226 = popcount38_5cwm_core_224 ^ popcount38_5cwm_core_214;
  assign popcount38_5cwm_core_227 = popcount38_5cwm_core_224 & popcount38_5cwm_core_214;
  assign popcount38_5cwm_core_228 = popcount38_5cwm_core_225 | popcount38_5cwm_core_227;
  assign popcount38_5cwm_core_231 = popcount38_5cwm_core_205 ^ popcount38_5cwm_core_222;
  assign popcount38_5cwm_core_232 = popcount38_5cwm_core_205 & popcount38_5cwm_core_222;
  assign popcount38_5cwm_core_233 = popcount38_5cwm_core_209 ^ popcount38_5cwm_core_226;
  assign popcount38_5cwm_core_234 = popcount38_5cwm_core_209 & popcount38_5cwm_core_226;
  assign popcount38_5cwm_core_235 = popcount38_5cwm_core_233 ^ popcount38_5cwm_core_232;
  assign popcount38_5cwm_core_236 = popcount38_5cwm_core_233 & popcount38_5cwm_core_232;
  assign popcount38_5cwm_core_237 = popcount38_5cwm_core_234 | popcount38_5cwm_core_236;
  assign popcount38_5cwm_core_238 = popcount38_5cwm_core_211 ^ popcount38_5cwm_core_228;
  assign popcount38_5cwm_core_239 = popcount38_5cwm_core_211 & popcount38_5cwm_core_228;
  assign popcount38_5cwm_core_240 = popcount38_5cwm_core_238 ^ popcount38_5cwm_core_237;
  assign popcount38_5cwm_core_241 = popcount38_5cwm_core_238 & popcount38_5cwm_core_237;
  assign popcount38_5cwm_core_242 = popcount38_5cwm_core_239 | popcount38_5cwm_core_241;
  assign popcount38_5cwm_core_244 = input_a[29] ^ input_a[2];
  assign popcount38_5cwm_core_246 = ~(input_a[3] ^ input_a[36]);
  assign popcount38_5cwm_core_248_not = ~popcount38_5cwm_core_231;
  assign popcount38_5cwm_core_250 = popcount38_5cwm_core_185 ^ popcount38_5cwm_core_235;
  assign popcount38_5cwm_core_251 = popcount38_5cwm_core_185 & popcount38_5cwm_core_235;
  assign popcount38_5cwm_core_252 = popcount38_5cwm_core_250 ^ popcount38_5cwm_core_231;
  assign popcount38_5cwm_core_253 = popcount38_5cwm_core_250 & popcount38_5cwm_core_231;
  assign popcount38_5cwm_core_254 = popcount38_5cwm_core_251 | popcount38_5cwm_core_253;
  assign popcount38_5cwm_core_255 = popcount38_5cwm_core_192 ^ popcount38_5cwm_core_240;
  assign popcount38_5cwm_core_256 = popcount38_5cwm_core_192 & popcount38_5cwm_core_240;
  assign popcount38_5cwm_core_257 = popcount38_5cwm_core_255 ^ popcount38_5cwm_core_254;
  assign popcount38_5cwm_core_258 = popcount38_5cwm_core_255 & popcount38_5cwm_core_254;
  assign popcount38_5cwm_core_259 = popcount38_5cwm_core_256 | popcount38_5cwm_core_258;
  assign popcount38_5cwm_core_260 = popcount38_5cwm_core_191 ^ popcount38_5cwm_core_242;
  assign popcount38_5cwm_core_261 = popcount38_5cwm_core_191 & popcount38_5cwm_core_242;
  assign popcount38_5cwm_core_262 = popcount38_5cwm_core_260 ^ popcount38_5cwm_core_259;
  assign popcount38_5cwm_core_263 = popcount38_5cwm_core_260 & popcount38_5cwm_core_259;
  assign popcount38_5cwm_core_264 = popcount38_5cwm_core_261 | popcount38_5cwm_core_263;
  assign popcount38_5cwm_core_266 = ~input_a[37];
  assign popcount38_5cwm_core_268 = ~(input_a[7] ^ input_a[32]);
  assign popcount38_5cwm_core_269 = input_a[28] | input_a[2];
  assign popcount38_5cwm_core_270 = input_a[4] ^ popcount38_5cwm_core_248_not;
  assign popcount38_5cwm_core_271 = input_a[4] & popcount38_5cwm_core_248_not;
  assign popcount38_5cwm_core_272 = popcount38_5cwm_core_070 ^ popcount38_5cwm_core_252;
  assign popcount38_5cwm_core_273 = popcount38_5cwm_core_070 & popcount38_5cwm_core_252;
  assign popcount38_5cwm_core_274 = popcount38_5cwm_core_272 ^ popcount38_5cwm_core_271;
  assign popcount38_5cwm_core_275 = popcount38_5cwm_core_272 & popcount38_5cwm_core_271;
  assign popcount38_5cwm_core_276 = popcount38_5cwm_core_273 | popcount38_5cwm_core_275;
  assign popcount38_5cwm_core_277 = popcount38_5cwm_core_142 ^ popcount38_5cwm_core_257;
  assign popcount38_5cwm_core_278 = popcount38_5cwm_core_142 & popcount38_5cwm_core_257;
  assign popcount38_5cwm_core_279 = popcount38_5cwm_core_277 ^ popcount38_5cwm_core_276;
  assign popcount38_5cwm_core_280 = popcount38_5cwm_core_277 & popcount38_5cwm_core_276;
  assign popcount38_5cwm_core_281 = popcount38_5cwm_core_278 | popcount38_5cwm_core_280;
  assign popcount38_5cwm_core_282 = popcount38_5cwm_core_144 ^ popcount38_5cwm_core_262;
  assign popcount38_5cwm_core_283 = popcount38_5cwm_core_144 & popcount38_5cwm_core_262;
  assign popcount38_5cwm_core_284 = popcount38_5cwm_core_282 ^ popcount38_5cwm_core_281;
  assign popcount38_5cwm_core_285 = popcount38_5cwm_core_282 & popcount38_5cwm_core_281;
  assign popcount38_5cwm_core_286 = popcount38_5cwm_core_283 | popcount38_5cwm_core_285;
  assign popcount38_5cwm_core_288 = ~input_a[0];
  assign popcount38_5cwm_core_289 = popcount38_5cwm_core_264 ^ popcount38_5cwm_core_286;
  assign popcount38_5cwm_core_290 = popcount38_5cwm_core_264 & popcount38_5cwm_core_286;
  assign popcount38_5cwm_core_291 = ~(input_a[28] & input_a[30]);
  assign popcount38_5cwm_core_292 = input_a[0] & input_a[23];
  assign popcount38_5cwm_core_294 = ~(input_a[13] ^ input_a[1]);
  assign popcount38_5cwm_core_295 = ~(input_a[19] | input_a[11]);
  assign popcount38_5cwm_core_296 = input_a[24] & input_a[36];

  assign popcount38_5cwm_out[0] = popcount38_5cwm_core_270;
  assign popcount38_5cwm_out[1] = popcount38_5cwm_core_274;
  assign popcount38_5cwm_out[2] = popcount38_5cwm_core_279;
  assign popcount38_5cwm_out[3] = popcount38_5cwm_core_284;
  assign popcount38_5cwm_out[4] = popcount38_5cwm_core_289;
  assign popcount38_5cwm_out[5] = popcount38_5cwm_core_290;
endmodule