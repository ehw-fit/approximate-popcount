// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.94951
// WCE=20.0
// EP=0.836311%
// Printed PDK parameters:
//  Area=60000140.0
//  Delay=74411048.0
//  Power=3378300.0

module popcount39_wtue(input [38:0] input_a, output [5:0] popcount39_wtue_out);
  wire popcount39_wtue_core_041;
  wire popcount39_wtue_core_042;
  wire popcount39_wtue_core_043;
  wire popcount39_wtue_core_044;
  wire popcount39_wtue_core_045;
  wire popcount39_wtue_core_046;
  wire popcount39_wtue_core_049;
  wire popcount39_wtue_core_050;
  wire popcount39_wtue_core_053;
  wire popcount39_wtue_core_055;
  wire popcount39_wtue_core_056;
  wire popcount39_wtue_core_059;
  wire popcount39_wtue_core_060;
  wire popcount39_wtue_core_062;
  wire popcount39_wtue_core_064;
  wire popcount39_wtue_core_067;
  wire popcount39_wtue_core_069;
  wire popcount39_wtue_core_071;
  wire popcount39_wtue_core_072;
  wire popcount39_wtue_core_073;
  wire popcount39_wtue_core_075;
  wire popcount39_wtue_core_078;
  wire popcount39_wtue_core_079;
  wire popcount39_wtue_core_083;
  wire popcount39_wtue_core_084;
  wire popcount39_wtue_core_085;
  wire popcount39_wtue_core_086;
  wire popcount39_wtue_core_089;
  wire popcount39_wtue_core_090;
  wire popcount39_wtue_core_091;
  wire popcount39_wtue_core_092;
  wire popcount39_wtue_core_093;
  wire popcount39_wtue_core_096;
  wire popcount39_wtue_core_098;
  wire popcount39_wtue_core_100;
  wire popcount39_wtue_core_101;
  wire popcount39_wtue_core_102;
  wire popcount39_wtue_core_103;
  wire popcount39_wtue_core_104;
  wire popcount39_wtue_core_106;
  wire popcount39_wtue_core_107;
  wire popcount39_wtue_core_108;
  wire popcount39_wtue_core_109;
  wire popcount39_wtue_core_110;
  wire popcount39_wtue_core_111;
  wire popcount39_wtue_core_113;
  wire popcount39_wtue_core_115;
  wire popcount39_wtue_core_117;
  wire popcount39_wtue_core_118;
  wire popcount39_wtue_core_119;
  wire popcount39_wtue_core_120;
  wire popcount39_wtue_core_121;
  wire popcount39_wtue_core_122;
  wire popcount39_wtue_core_123;
  wire popcount39_wtue_core_124;
  wire popcount39_wtue_core_125;
  wire popcount39_wtue_core_126;
  wire popcount39_wtue_core_127;
  wire popcount39_wtue_core_128;
  wire popcount39_wtue_core_132;
  wire popcount39_wtue_core_133;
  wire popcount39_wtue_core_134;
  wire popcount39_wtue_core_135;
  wire popcount39_wtue_core_136;
  wire popcount39_wtue_core_137;
  wire popcount39_wtue_core_139;
  wire popcount39_wtue_core_141;
  wire popcount39_wtue_core_142;
  wire popcount39_wtue_core_143;
  wire popcount39_wtue_core_144;
  wire popcount39_wtue_core_145;
  wire popcount39_wtue_core_146;
  wire popcount39_wtue_core_148;
  wire popcount39_wtue_core_154;
  wire popcount39_wtue_core_156;
  wire popcount39_wtue_core_157;
  wire popcount39_wtue_core_158;
  wire popcount39_wtue_core_159;
  wire popcount39_wtue_core_160;
  wire popcount39_wtue_core_161;
  wire popcount39_wtue_core_162;
  wire popcount39_wtue_core_164;
  wire popcount39_wtue_core_165;
  wire popcount39_wtue_core_166;
  wire popcount39_wtue_core_167;
  wire popcount39_wtue_core_168;
  wire popcount39_wtue_core_169;
  wire popcount39_wtue_core_170;
  wire popcount39_wtue_core_173;
  wire popcount39_wtue_core_175;
  wire popcount39_wtue_core_176;
  wire popcount39_wtue_core_177;
  wire popcount39_wtue_core_178;
  wire popcount39_wtue_core_179;
  wire popcount39_wtue_core_180;
  wire popcount39_wtue_core_181;
  wire popcount39_wtue_core_182;
  wire popcount39_wtue_core_184;
  wire popcount39_wtue_core_185;
  wire popcount39_wtue_core_191;
  wire popcount39_wtue_core_192;
  wire popcount39_wtue_core_194;
  wire popcount39_wtue_core_195;
  wire popcount39_wtue_core_196;
  wire popcount39_wtue_core_199;
  wire popcount39_wtue_core_203;
  wire popcount39_wtue_core_205;
  wire popcount39_wtue_core_206;
  wire popcount39_wtue_core_207;
  wire popcount39_wtue_core_208;
  wire popcount39_wtue_core_211;
  wire popcount39_wtue_core_213;
  wire popcount39_wtue_core_214;
  wire popcount39_wtue_core_215;
  wire popcount39_wtue_core_216;
  wire popcount39_wtue_core_221;
  wire popcount39_wtue_core_225;
  wire popcount39_wtue_core_226;
  wire popcount39_wtue_core_227;
  wire popcount39_wtue_core_228;
  wire popcount39_wtue_core_229;
  wire popcount39_wtue_core_230;
  wire popcount39_wtue_core_232;
  wire popcount39_wtue_core_233;
  wire popcount39_wtue_core_234;
  wire popcount39_wtue_core_235;
  wire popcount39_wtue_core_236;
  wire popcount39_wtue_core_237;
  wire popcount39_wtue_core_238;
  wire popcount39_wtue_core_240;
  wire popcount39_wtue_core_241;
  wire popcount39_wtue_core_242;
  wire popcount39_wtue_core_243_not;
  wire popcount39_wtue_core_245;
  wire popcount39_wtue_core_246;
  wire popcount39_wtue_core_247;
  wire popcount39_wtue_core_250;
  wire popcount39_wtue_core_258;
  wire popcount39_wtue_core_259;
  wire popcount39_wtue_core_260;
  wire popcount39_wtue_core_261;
  wire popcount39_wtue_core_265;
  wire popcount39_wtue_core_266;
  wire popcount39_wtue_core_267;
  wire popcount39_wtue_core_268;
  wire popcount39_wtue_core_269;
  wire popcount39_wtue_core_270;
  wire popcount39_wtue_core_271;
  wire popcount39_wtue_core_272;
  wire popcount39_wtue_core_273;
  wire popcount39_wtue_core_275;
  wire popcount39_wtue_core_277;
  wire popcount39_wtue_core_278;
  wire popcount39_wtue_core_279;
  wire popcount39_wtue_core_281;
  wire popcount39_wtue_core_282;
  wire popcount39_wtue_core_283;
  wire popcount39_wtue_core_285;
  wire popcount39_wtue_core_287;
  wire popcount39_wtue_core_288;
  wire popcount39_wtue_core_289;
  wire popcount39_wtue_core_290;
  wire popcount39_wtue_core_291;
  wire popcount39_wtue_core_292;
  wire popcount39_wtue_core_293;
  wire popcount39_wtue_core_294;
  wire popcount39_wtue_core_295;
  wire popcount39_wtue_core_296;
  wire popcount39_wtue_core_298;
  wire popcount39_wtue_core_299;
  wire popcount39_wtue_core_302;
  wire popcount39_wtue_core_304;
  wire popcount39_wtue_core_305;

  assign popcount39_wtue_core_041 = input_a[27] | input_a[9];
  assign popcount39_wtue_core_042 = input_a[32] ^ input_a[28];
  assign popcount39_wtue_core_043 = ~(input_a[4] & input_a[3]);
  assign popcount39_wtue_core_044 = ~input_a[5];
  assign popcount39_wtue_core_045 = ~(input_a[35] & input_a[34]);
  assign popcount39_wtue_core_046 = input_a[12] & input_a[1];
  assign popcount39_wtue_core_049 = input_a[8] ^ popcount39_wtue_core_046;
  assign popcount39_wtue_core_050 = input_a[8] & popcount39_wtue_core_046;
  assign popcount39_wtue_core_053 = input_a[19] ^ input_a[29];
  assign popcount39_wtue_core_055 = input_a[34] & input_a[35];
  assign popcount39_wtue_core_056 = ~(input_a[2] | input_a[35]);
  assign popcount39_wtue_core_059 = ~(input_a[0] ^ input_a[6]);
  assign popcount39_wtue_core_060 = input_a[19] | input_a[35];
  assign popcount39_wtue_core_062 = input_a[23] | input_a[13];
  assign popcount39_wtue_core_064 = input_a[31] | input_a[29];
  assign popcount39_wtue_core_067 = ~(input_a[15] ^ input_a[18]);
  assign popcount39_wtue_core_069 = ~input_a[36];
  assign popcount39_wtue_core_071 = ~(popcount39_wtue_core_049 & popcount39_wtue_core_064);
  assign popcount39_wtue_core_072 = popcount39_wtue_core_049 & popcount39_wtue_core_064;
  assign popcount39_wtue_core_073 = popcount39_wtue_core_071 ^ input_a[16];
  assign popcount39_wtue_core_075 = popcount39_wtue_core_072 | input_a[16];
  assign popcount39_wtue_core_078 = popcount39_wtue_core_050 ^ popcount39_wtue_core_075;
  assign popcount39_wtue_core_079 = popcount39_wtue_core_050 & input_a[16];
  assign popcount39_wtue_core_083 = input_a[24] ^ input_a[5];
  assign popcount39_wtue_core_084 = input_a[36] & input_a[18];
  assign popcount39_wtue_core_085 = ~(input_a[10] & input_a[27]);
  assign popcount39_wtue_core_086 = input_a[3] | input_a[6];
  assign popcount39_wtue_core_089 = ~(input_a[28] & input_a[11]);
  assign popcount39_wtue_core_090 = input_a[28] & input_a[11];
  assign popcount39_wtue_core_091 = ~(input_a[17] & input_a[27]);
  assign popcount39_wtue_core_092 = ~(input_a[5] & input_a[5]);
  assign popcount39_wtue_core_093 = popcount39_wtue_core_084 ^ popcount39_wtue_core_089;
  assign popcount39_wtue_core_096 = ~(input_a[0] & input_a[33]);
  assign popcount39_wtue_core_098 = popcount39_wtue_core_090 | popcount39_wtue_core_084;
  assign popcount39_wtue_core_100 = ~(input_a[7] & input_a[16]);
  assign popcount39_wtue_core_101 = input_a[37] & input_a[7];
  assign popcount39_wtue_core_102 = input_a[32] ^ input_a[12];
  assign popcount39_wtue_core_103 = input_a[3] & input_a[9];
  assign popcount39_wtue_core_104 = ~input_a[20];
  assign popcount39_wtue_core_106 = popcount39_wtue_core_103 ^ input_a[6];
  assign popcount39_wtue_core_107 = popcount39_wtue_core_103 & input_a[6];
  assign popcount39_wtue_core_108 = input_a[28] | input_a[3];
  assign popcount39_wtue_core_109 = ~(input_a[18] ^ input_a[8]);
  assign popcount39_wtue_core_110 = popcount39_wtue_core_101 ^ popcount39_wtue_core_106;
  assign popcount39_wtue_core_111 = popcount39_wtue_core_101 & popcount39_wtue_core_106;
  assign popcount39_wtue_core_113 = ~(input_a[9] & input_a[4]);
  assign popcount39_wtue_core_115 = popcount39_wtue_core_107 | popcount39_wtue_core_111;
  assign popcount39_wtue_core_117 = input_a[33] | input_a[17];
  assign popcount39_wtue_core_118 = input_a[26] & input_a[27];
  assign popcount39_wtue_core_119 = popcount39_wtue_core_093 ^ popcount39_wtue_core_110;
  assign popcount39_wtue_core_120 = popcount39_wtue_core_093 & popcount39_wtue_core_110;
  assign popcount39_wtue_core_121 = popcount39_wtue_core_119 ^ popcount39_wtue_core_118;
  assign popcount39_wtue_core_122 = popcount39_wtue_core_119 & popcount39_wtue_core_118;
  assign popcount39_wtue_core_123 = popcount39_wtue_core_120 | popcount39_wtue_core_122;
  assign popcount39_wtue_core_124 = popcount39_wtue_core_098 ^ popcount39_wtue_core_115;
  assign popcount39_wtue_core_125 = popcount39_wtue_core_098 & popcount39_wtue_core_115;
  assign popcount39_wtue_core_126 = popcount39_wtue_core_124 ^ popcount39_wtue_core_123;
  assign popcount39_wtue_core_127 = popcount39_wtue_core_124 & popcount39_wtue_core_123;
  assign popcount39_wtue_core_128 = popcount39_wtue_core_125 | popcount39_wtue_core_127;
  assign popcount39_wtue_core_132 = ~input_a[29];
  assign popcount39_wtue_core_133 = input_a[27] | input_a[19];
  assign popcount39_wtue_core_134 = ~(input_a[20] & input_a[26]);
  assign popcount39_wtue_core_135 = input_a[31] ^ input_a[5];
  assign popcount39_wtue_core_136 = popcount39_wtue_core_073 ^ popcount39_wtue_core_121;
  assign popcount39_wtue_core_137 = popcount39_wtue_core_073 & popcount39_wtue_core_121;
  assign popcount39_wtue_core_139 = ~(input_a[26] ^ input_a[13]);
  assign popcount39_wtue_core_141 = popcount39_wtue_core_078 ^ popcount39_wtue_core_126;
  assign popcount39_wtue_core_142 = popcount39_wtue_core_078 & popcount39_wtue_core_126;
  assign popcount39_wtue_core_143 = popcount39_wtue_core_141 ^ popcount39_wtue_core_137;
  assign popcount39_wtue_core_144 = popcount39_wtue_core_141 & popcount39_wtue_core_137;
  assign popcount39_wtue_core_145 = popcount39_wtue_core_142 | popcount39_wtue_core_144;
  assign popcount39_wtue_core_146 = popcount39_wtue_core_079 | popcount39_wtue_core_128;
  assign popcount39_wtue_core_148 = popcount39_wtue_core_146 ^ popcount39_wtue_core_145;
  assign popcount39_wtue_core_154 = ~(input_a[30] | input_a[25]);
  assign popcount39_wtue_core_156 = input_a[19] ^ input_a[20];
  assign popcount39_wtue_core_157 = input_a[19] & input_a[20];
  assign popcount39_wtue_core_158 = ~(input_a[22] & input_a[23]);
  assign popcount39_wtue_core_159 = input_a[22] & input_a[23];
  assign popcount39_wtue_core_160 = input_a[21] ^ popcount39_wtue_core_158;
  assign popcount39_wtue_core_161 = ~(input_a[32] & input_a[29]);
  assign popcount39_wtue_core_162 = popcount39_wtue_core_159 | input_a[21];
  assign popcount39_wtue_core_164 = ~(input_a[33] & input_a[26]);
  assign popcount39_wtue_core_165 = popcount39_wtue_core_156 & popcount39_wtue_core_160;
  assign popcount39_wtue_core_166 = popcount39_wtue_core_157 ^ popcount39_wtue_core_162;
  assign popcount39_wtue_core_167 = popcount39_wtue_core_157 & popcount39_wtue_core_162;
  assign popcount39_wtue_core_168 = popcount39_wtue_core_166 ^ popcount39_wtue_core_165;
  assign popcount39_wtue_core_169 = input_a[21] & popcount39_wtue_core_165;
  assign popcount39_wtue_core_170 = popcount39_wtue_core_167 | popcount39_wtue_core_169;
  assign popcount39_wtue_core_173 = ~(input_a[35] & input_a[30]);
  assign popcount39_wtue_core_175 = input_a[36] & input_a[20];
  assign popcount39_wtue_core_176 = ~(input_a[16] & input_a[21]);
  assign popcount39_wtue_core_177 = input_a[34] ^ input_a[35];
  assign popcount39_wtue_core_178 = ~input_a[37];
  assign popcount39_wtue_core_179 = input_a[18] | input_a[14];
  assign popcount39_wtue_core_180 = input_a[19] | input_a[21];
  assign popcount39_wtue_core_181 = input_a[27] | input_a[21];
  assign popcount39_wtue_core_182 = ~(input_a[23] | input_a[30]);
  assign popcount39_wtue_core_184 = input_a[17] ^ input_a[12];
  assign popcount39_wtue_core_185 = input_a[8] ^ input_a[31];
  assign popcount39_wtue_core_191 = input_a[13] & input_a[4];
  assign popcount39_wtue_core_192 = ~popcount39_wtue_core_168;
  assign popcount39_wtue_core_194 = popcount39_wtue_core_192 ^ popcount39_wtue_core_191;
  assign popcount39_wtue_core_195 = input_a[4] & popcount39_wtue_core_191;
  assign popcount39_wtue_core_196 = popcount39_wtue_core_168 | popcount39_wtue_core_195;
  assign popcount39_wtue_core_199 = popcount39_wtue_core_170 ^ popcount39_wtue_core_196;
  assign popcount39_wtue_core_203 = input_a[26] ^ input_a[38];
  assign popcount39_wtue_core_205 = ~input_a[1];
  assign popcount39_wtue_core_206 = ~(input_a[31] ^ input_a[32]);
  assign popcount39_wtue_core_207 = input_a[3] ^ input_a[13];
  assign popcount39_wtue_core_208 = input_a[19] ^ input_a[2];
  assign popcount39_wtue_core_211 = ~(input_a[37] ^ input_a[31]);
  assign popcount39_wtue_core_213 = input_a[25] & input_a[29];
  assign popcount39_wtue_core_214 = input_a[20] | input_a[22];
  assign popcount39_wtue_core_215 = ~(input_a[28] | input_a[0]);
  assign popcount39_wtue_core_216 = input_a[7] ^ input_a[26];
  assign popcount39_wtue_core_221 = input_a[34] ^ input_a[33];
  assign popcount39_wtue_core_225 = input_a[32] & input_a[14];
  assign popcount39_wtue_core_226 = input_a[23] | input_a[22];
  assign popcount39_wtue_core_227 = input_a[10] & input_a[34];
  assign popcount39_wtue_core_228 = input_a[24] ^ input_a[2];
  assign popcount39_wtue_core_229 = input_a[30] & popcount39_wtue_core_226;
  assign popcount39_wtue_core_230 = popcount39_wtue_core_227 | popcount39_wtue_core_229;
  assign popcount39_wtue_core_232 = input_a[9] & input_a[19];
  assign popcount39_wtue_core_233 = input_a[2] & input_a[0];
  assign popcount39_wtue_core_234 = popcount39_wtue_core_225 ^ popcount39_wtue_core_230;
  assign popcount39_wtue_core_235 = popcount39_wtue_core_225 & popcount39_wtue_core_230;
  assign popcount39_wtue_core_236 = popcount39_wtue_core_234 ^ popcount39_wtue_core_233;
  assign popcount39_wtue_core_237 = popcount39_wtue_core_234 & popcount39_wtue_core_233;
  assign popcount39_wtue_core_238 = popcount39_wtue_core_235 | popcount39_wtue_core_237;
  assign popcount39_wtue_core_240 = ~(input_a[33] | input_a[5]);
  assign popcount39_wtue_core_241 = input_a[17] & input_a[5];
  assign popcount39_wtue_core_242 = input_a[25] & input_a[33];
  assign popcount39_wtue_core_243_not = ~popcount39_wtue_core_236;
  assign popcount39_wtue_core_245 = popcount39_wtue_core_243_not ^ popcount39_wtue_core_242;
  assign popcount39_wtue_core_246 = input_a[25] & input_a[33];
  assign popcount39_wtue_core_247 = popcount39_wtue_core_236 | popcount39_wtue_core_246;
  assign popcount39_wtue_core_250 = popcount39_wtue_core_238 ^ popcount39_wtue_core_247;
  assign popcount39_wtue_core_258 = ~(input_a[36] & input_a[12]);
  assign popcount39_wtue_core_259 = ~(input_a[36] | input_a[7]);
  assign popcount39_wtue_core_260 = popcount39_wtue_core_194 ^ popcount39_wtue_core_245;
  assign popcount39_wtue_core_261 = popcount39_wtue_core_194 & popcount39_wtue_core_245;
  assign popcount39_wtue_core_265 = ~(popcount39_wtue_core_199 & popcount39_wtue_core_250);
  assign popcount39_wtue_core_266 = popcount39_wtue_core_199 & popcount39_wtue_core_250;
  assign popcount39_wtue_core_267 = popcount39_wtue_core_265 ^ popcount39_wtue_core_261;
  assign popcount39_wtue_core_268 = popcount39_wtue_core_265 & popcount39_wtue_core_261;
  assign popcount39_wtue_core_269 = popcount39_wtue_core_266 | popcount39_wtue_core_268;
  assign popcount39_wtue_core_270 = popcount39_wtue_core_170 | popcount39_wtue_core_238;
  assign popcount39_wtue_core_271 = ~input_a[14];
  assign popcount39_wtue_core_272 = popcount39_wtue_core_270 | popcount39_wtue_core_269;
  assign popcount39_wtue_core_273 = ~input_a[7];
  assign popcount39_wtue_core_275 = input_a[18] | input_a[17];
  assign popcount39_wtue_core_277 = ~(input_a[12] | input_a[20]);
  assign popcount39_wtue_core_278 = input_a[7] | input_a[8];
  assign popcount39_wtue_core_279 = input_a[12] & input_a[2];
  assign popcount39_wtue_core_281 = input_a[1] ^ input_a[35];
  assign popcount39_wtue_core_282 = popcount39_wtue_core_136 ^ popcount39_wtue_core_260;
  assign popcount39_wtue_core_283 = popcount39_wtue_core_136 & popcount39_wtue_core_260;
  assign popcount39_wtue_core_285 = ~input_a[8];
  assign popcount39_wtue_core_287 = popcount39_wtue_core_143 ^ popcount39_wtue_core_267;
  assign popcount39_wtue_core_288 = popcount39_wtue_core_143 & popcount39_wtue_core_267;
  assign popcount39_wtue_core_289 = popcount39_wtue_core_287 ^ popcount39_wtue_core_283;
  assign popcount39_wtue_core_290 = popcount39_wtue_core_287 & popcount39_wtue_core_283;
  assign popcount39_wtue_core_291 = popcount39_wtue_core_288 | popcount39_wtue_core_290;
  assign popcount39_wtue_core_292 = popcount39_wtue_core_148 ^ popcount39_wtue_core_272;
  assign popcount39_wtue_core_293 = popcount39_wtue_core_148 & popcount39_wtue_core_272;
  assign popcount39_wtue_core_294 = popcount39_wtue_core_292 ^ popcount39_wtue_core_291;
  assign popcount39_wtue_core_295 = popcount39_wtue_core_292 & popcount39_wtue_core_291;
  assign popcount39_wtue_core_296 = popcount39_wtue_core_293 | popcount39_wtue_core_295;
  assign popcount39_wtue_core_298 = input_a[20] | input_a[11];
  assign popcount39_wtue_core_299 = popcount39_wtue_core_146 | popcount39_wtue_core_296;
  assign popcount39_wtue_core_302 = input_a[13] & input_a[11];
  assign popcount39_wtue_core_304 = input_a[11] ^ input_a[11];
  assign popcount39_wtue_core_305 = input_a[17] | input_a[25];

  assign popcount39_wtue_out[0] = input_a[5];
  assign popcount39_wtue_out[1] = popcount39_wtue_core_282;
  assign popcount39_wtue_out[2] = popcount39_wtue_core_289;
  assign popcount39_wtue_out[3] = popcount39_wtue_core_294;
  assign popcount39_wtue_out[4] = popcount39_wtue_core_299;
  assign popcount39_wtue_out[5] = 1'b0;
endmodule