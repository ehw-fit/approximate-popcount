// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.09224
// WCE=14.0
// EP=0.850554%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_gp0i(input [27:0] input_a, output [4:0] popcount28_gp0i_out);
  wire popcount28_gp0i_core_030;
  wire popcount28_gp0i_core_031;
  wire popcount28_gp0i_core_032;
  wire popcount28_gp0i_core_033;
  wire popcount28_gp0i_core_034;
  wire popcount28_gp0i_core_035;
  wire popcount28_gp0i_core_037;
  wire popcount28_gp0i_core_038;
  wire popcount28_gp0i_core_039;
  wire popcount28_gp0i_core_041;
  wire popcount28_gp0i_core_042;
  wire popcount28_gp0i_core_044;
  wire popcount28_gp0i_core_045;
  wire popcount28_gp0i_core_046;
  wire popcount28_gp0i_core_049;
  wire popcount28_gp0i_core_050;
  wire popcount28_gp0i_core_053;
  wire popcount28_gp0i_core_058;
  wire popcount28_gp0i_core_059;
  wire popcount28_gp0i_core_060;
  wire popcount28_gp0i_core_061;
  wire popcount28_gp0i_core_062;
  wire popcount28_gp0i_core_064;
  wire popcount28_gp0i_core_065;
  wire popcount28_gp0i_core_066;
  wire popcount28_gp0i_core_069;
  wire popcount28_gp0i_core_071;
  wire popcount28_gp0i_core_072;
  wire popcount28_gp0i_core_073;
  wire popcount28_gp0i_core_075;
  wire popcount28_gp0i_core_078;
  wire popcount28_gp0i_core_079;
  wire popcount28_gp0i_core_080;
  wire popcount28_gp0i_core_081;
  wire popcount28_gp0i_core_083;
  wire popcount28_gp0i_core_084;
  wire popcount28_gp0i_core_085;
  wire popcount28_gp0i_core_086;
  wire popcount28_gp0i_core_090;
  wire popcount28_gp0i_core_092;
  wire popcount28_gp0i_core_096;
  wire popcount28_gp0i_core_097;
  wire popcount28_gp0i_core_098;
  wire popcount28_gp0i_core_099;
  wire popcount28_gp0i_core_100;
  wire popcount28_gp0i_core_101;
  wire popcount28_gp0i_core_103;
  wire popcount28_gp0i_core_104;
  wire popcount28_gp0i_core_105;
  wire popcount28_gp0i_core_106_not;
  wire popcount28_gp0i_core_107;
  wire popcount28_gp0i_core_108;
  wire popcount28_gp0i_core_109;
  wire popcount28_gp0i_core_111;
  wire popcount28_gp0i_core_112;
  wire popcount28_gp0i_core_114;
  wire popcount28_gp0i_core_115;
  wire popcount28_gp0i_core_116;
  wire popcount28_gp0i_core_117_not;
  wire popcount28_gp0i_core_118;
  wire popcount28_gp0i_core_119;
  wire popcount28_gp0i_core_120;
  wire popcount28_gp0i_core_121;
  wire popcount28_gp0i_core_122;
  wire popcount28_gp0i_core_124;
  wire popcount28_gp0i_core_125;
  wire popcount28_gp0i_core_126;
  wire popcount28_gp0i_core_127;
  wire popcount28_gp0i_core_128;
  wire popcount28_gp0i_core_130;
  wire popcount28_gp0i_core_131;
  wire popcount28_gp0i_core_132;
  wire popcount28_gp0i_core_135;
  wire popcount28_gp0i_core_136;
  wire popcount28_gp0i_core_137;
  wire popcount28_gp0i_core_140;
  wire popcount28_gp0i_core_144;
  wire popcount28_gp0i_core_145;
  wire popcount28_gp0i_core_147;
  wire popcount28_gp0i_core_151;
  wire popcount28_gp0i_core_153;
  wire popcount28_gp0i_core_154;
  wire popcount28_gp0i_core_155;
  wire popcount28_gp0i_core_156;
  wire popcount28_gp0i_core_157;
  wire popcount28_gp0i_core_158;
  wire popcount28_gp0i_core_159;
  wire popcount28_gp0i_core_161;
  wire popcount28_gp0i_core_162;
  wire popcount28_gp0i_core_165;
  wire popcount28_gp0i_core_166;
  wire popcount28_gp0i_core_167;
  wire popcount28_gp0i_core_169;
  wire popcount28_gp0i_core_170_not;
  wire popcount28_gp0i_core_171;
  wire popcount28_gp0i_core_172;
  wire popcount28_gp0i_core_173;
  wire popcount28_gp0i_core_175_not;
  wire popcount28_gp0i_core_176;
  wire popcount28_gp0i_core_179;
  wire popcount28_gp0i_core_181;
  wire popcount28_gp0i_core_182;
  wire popcount28_gp0i_core_183;
  wire popcount28_gp0i_core_184;
  wire popcount28_gp0i_core_185;
  wire popcount28_gp0i_core_186;
  wire popcount28_gp0i_core_187;
  wire popcount28_gp0i_core_190;
  wire popcount28_gp0i_core_191;
  wire popcount28_gp0i_core_192_not;
  wire popcount28_gp0i_core_193;
  wire popcount28_gp0i_core_194;
  wire popcount28_gp0i_core_196;
  wire popcount28_gp0i_core_197;
  wire popcount28_gp0i_core_199;
  wire popcount28_gp0i_core_200;
  wire popcount28_gp0i_core_201;

  assign popcount28_gp0i_core_030 = input_a[9] & input_a[0];
  assign popcount28_gp0i_core_031 = ~(input_a[5] & input_a[5]);
  assign popcount28_gp0i_core_032 = ~(input_a[0] ^ input_a[24]);
  assign popcount28_gp0i_core_033 = input_a[10] & input_a[0];
  assign popcount28_gp0i_core_034 = input_a[11] | input_a[17];
  assign popcount28_gp0i_core_035 = ~input_a[12];
  assign popcount28_gp0i_core_037 = input_a[0] & input_a[12];
  assign popcount28_gp0i_core_038 = ~(input_a[3] | input_a[16]);
  assign popcount28_gp0i_core_039 = ~(input_a[19] ^ input_a[1]);
  assign popcount28_gp0i_core_041 = ~(input_a[0] & input_a[6]);
  assign popcount28_gp0i_core_042 = ~input_a[11];
  assign popcount28_gp0i_core_044 = input_a[15] & input_a[17];
  assign popcount28_gp0i_core_045 = ~(input_a[1] ^ input_a[23]);
  assign popcount28_gp0i_core_046 = input_a[12] & input_a[2];
  assign popcount28_gp0i_core_049 = ~input_a[19];
  assign popcount28_gp0i_core_050 = ~(input_a[16] ^ input_a[26]);
  assign popcount28_gp0i_core_053 = input_a[2] | input_a[20];
  assign popcount28_gp0i_core_058 = ~(input_a[15] | input_a[13]);
  assign popcount28_gp0i_core_059 = input_a[5] ^ input_a[10];
  assign popcount28_gp0i_core_060 = ~(input_a[16] | input_a[24]);
  assign popcount28_gp0i_core_061 = ~(input_a[20] & input_a[8]);
  assign popcount28_gp0i_core_062 = input_a[27] | input_a[14];
  assign popcount28_gp0i_core_064 = ~(input_a[27] ^ input_a[17]);
  assign popcount28_gp0i_core_065 = ~(input_a[20] ^ input_a[3]);
  assign popcount28_gp0i_core_066 = input_a[10] ^ input_a[3];
  assign popcount28_gp0i_core_069 = input_a[8] | input_a[10];
  assign popcount28_gp0i_core_071 = input_a[22] | input_a[12];
  assign popcount28_gp0i_core_072 = ~(input_a[21] ^ input_a[2]);
  assign popcount28_gp0i_core_073 = ~(input_a[16] | input_a[20]);
  assign popcount28_gp0i_core_075 = input_a[18] ^ input_a[4];
  assign popcount28_gp0i_core_078 = ~(input_a[1] ^ input_a[5]);
  assign popcount28_gp0i_core_079 = input_a[5] & input_a[15];
  assign popcount28_gp0i_core_080 = ~(input_a[18] ^ input_a[0]);
  assign popcount28_gp0i_core_081 = ~(input_a[26] & input_a[17]);
  assign popcount28_gp0i_core_083 = input_a[23] | input_a[26];
  assign popcount28_gp0i_core_084 = input_a[15] & input_a[8];
  assign popcount28_gp0i_core_085 = ~input_a[4];
  assign popcount28_gp0i_core_086 = input_a[21] ^ input_a[25];
  assign popcount28_gp0i_core_090 = input_a[0] | input_a[5];
  assign popcount28_gp0i_core_092 = input_a[8] | input_a[21];
  assign popcount28_gp0i_core_096 = input_a[7] & input_a[11];
  assign popcount28_gp0i_core_097 = input_a[0] & input_a[2];
  assign popcount28_gp0i_core_098 = input_a[17] & input_a[23];
  assign popcount28_gp0i_core_099 = ~(input_a[11] | input_a[13]);
  assign popcount28_gp0i_core_100 = ~(input_a[3] | input_a[26]);
  assign popcount28_gp0i_core_101 = input_a[14] ^ input_a[20];
  assign popcount28_gp0i_core_103 = ~(input_a[6] & input_a[6]);
  assign popcount28_gp0i_core_104 = input_a[21] ^ input_a[0];
  assign popcount28_gp0i_core_105 = input_a[7] & input_a[19];
  assign popcount28_gp0i_core_106_not = ~input_a[18];
  assign popcount28_gp0i_core_107 = input_a[15] & input_a[4];
  assign popcount28_gp0i_core_108 = ~(input_a[7] | input_a[16]);
  assign popcount28_gp0i_core_109 = input_a[13] & input_a[13];
  assign popcount28_gp0i_core_111 = input_a[21] ^ input_a[14];
  assign popcount28_gp0i_core_112 = ~(input_a[22] & input_a[23]);
  assign popcount28_gp0i_core_114 = ~input_a[26];
  assign popcount28_gp0i_core_115 = ~(input_a[7] | input_a[16]);
  assign popcount28_gp0i_core_116 = ~(input_a[4] ^ input_a[3]);
  assign popcount28_gp0i_core_117_not = ~input_a[27];
  assign popcount28_gp0i_core_118 = ~(input_a[10] & input_a[16]);
  assign popcount28_gp0i_core_119 = input_a[14] | input_a[3];
  assign popcount28_gp0i_core_120 = ~(input_a[8] & input_a[15]);
  assign popcount28_gp0i_core_121 = ~(input_a[1] ^ input_a[6]);
  assign popcount28_gp0i_core_122 = ~(input_a[24] & input_a[14]);
  assign popcount28_gp0i_core_124 = ~(input_a[1] | input_a[4]);
  assign popcount28_gp0i_core_125 = ~(input_a[14] ^ input_a[5]);
  assign popcount28_gp0i_core_126 = ~(input_a[0] ^ input_a[14]);
  assign popcount28_gp0i_core_127 = input_a[8] ^ input_a[15];
  assign popcount28_gp0i_core_128 = ~(input_a[4] | input_a[13]);
  assign popcount28_gp0i_core_130 = input_a[6] ^ input_a[5];
  assign popcount28_gp0i_core_131 = input_a[10] & input_a[7];
  assign popcount28_gp0i_core_132 = input_a[11] & input_a[27];
  assign popcount28_gp0i_core_135 = input_a[7] & input_a[1];
  assign popcount28_gp0i_core_136 = input_a[10] | input_a[8];
  assign popcount28_gp0i_core_137 = input_a[7] & input_a[26];
  assign popcount28_gp0i_core_140 = input_a[7] ^ input_a[18];
  assign popcount28_gp0i_core_144 = ~(input_a[2] | input_a[0]);
  assign popcount28_gp0i_core_145 = ~input_a[13];
  assign popcount28_gp0i_core_147 = input_a[24] & input_a[7];
  assign popcount28_gp0i_core_151 = ~(input_a[15] | input_a[8]);
  assign popcount28_gp0i_core_153 = ~(input_a[10] ^ input_a[27]);
  assign popcount28_gp0i_core_154 = input_a[24] & input_a[6];
  assign popcount28_gp0i_core_155 = ~(input_a[13] | input_a[18]);
  assign popcount28_gp0i_core_156 = ~(input_a[25] | input_a[2]);
  assign popcount28_gp0i_core_157 = input_a[20] | input_a[21];
  assign popcount28_gp0i_core_158 = ~(input_a[16] | input_a[25]);
  assign popcount28_gp0i_core_159 = ~input_a[7];
  assign popcount28_gp0i_core_161 = input_a[2] | input_a[3];
  assign popcount28_gp0i_core_162 = ~(input_a[17] ^ input_a[1]);
  assign popcount28_gp0i_core_165 = ~(input_a[20] ^ input_a[2]);
  assign popcount28_gp0i_core_166 = input_a[12] & input_a[10];
  assign popcount28_gp0i_core_167 = ~(input_a[11] & input_a[1]);
  assign popcount28_gp0i_core_169 = input_a[24] & input_a[4];
  assign popcount28_gp0i_core_170_not = ~input_a[19];
  assign popcount28_gp0i_core_171 = ~(input_a[6] & input_a[3]);
  assign popcount28_gp0i_core_172 = ~(input_a[14] | input_a[16]);
  assign popcount28_gp0i_core_173 = ~(input_a[10] & input_a[9]);
  assign popcount28_gp0i_core_175_not = ~input_a[15];
  assign popcount28_gp0i_core_176 = ~input_a[17];
  assign popcount28_gp0i_core_179 = ~(input_a[3] ^ input_a[0]);
  assign popcount28_gp0i_core_181 = ~(input_a[12] & input_a[0]);
  assign popcount28_gp0i_core_182 = input_a[13] ^ input_a[0];
  assign popcount28_gp0i_core_183 = ~(input_a[15] | input_a[11]);
  assign popcount28_gp0i_core_184 = input_a[5] & input_a[18];
  assign popcount28_gp0i_core_185 = ~(input_a[21] & input_a[27]);
  assign popcount28_gp0i_core_186 = ~input_a[13];
  assign popcount28_gp0i_core_187 = input_a[8] & input_a[6];
  assign popcount28_gp0i_core_190 = input_a[24] & input_a[14];
  assign popcount28_gp0i_core_191 = input_a[19] | input_a[5];
  assign popcount28_gp0i_core_192_not = ~input_a[22];
  assign popcount28_gp0i_core_193 = input_a[9] | input_a[26];
  assign popcount28_gp0i_core_194 = input_a[5] | input_a[12];
  assign popcount28_gp0i_core_196 = input_a[13] & input_a[25];
  assign popcount28_gp0i_core_197 = input_a[17] & input_a[8];
  assign popcount28_gp0i_core_199 = ~(input_a[24] | input_a[16]);
  assign popcount28_gp0i_core_200 = ~input_a[13];
  assign popcount28_gp0i_core_201 = ~input_a[4];

  assign popcount28_gp0i_out[0] = input_a[26];
  assign popcount28_gp0i_out[1] = 1'b1;
  assign popcount28_gp0i_out[2] = 1'b1;
  assign popcount28_gp0i_out[3] = 1'b1;
  assign popcount28_gp0i_out[4] = 1'b0;
endmodule