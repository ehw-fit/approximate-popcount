// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5001
// WCE=37.0
// EP=0.999861%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_y9gs(input [31:0] input_a, output [5:0] popcount32_y9gs_out);
  wire popcount32_y9gs_core_034;
  wire popcount32_y9gs_core_035;
  wire popcount32_y9gs_core_037;
  wire popcount32_y9gs_core_038;
  wire popcount32_y9gs_core_039;
  wire popcount32_y9gs_core_040;
  wire popcount32_y9gs_core_043;
  wire popcount32_y9gs_core_045_not;
  wire popcount32_y9gs_core_046_not;
  wire popcount32_y9gs_core_048;
  wire popcount32_y9gs_core_050;
  wire popcount32_y9gs_core_051;
  wire popcount32_y9gs_core_052;
  wire popcount32_y9gs_core_053;
  wire popcount32_y9gs_core_054;
  wire popcount32_y9gs_core_055;
  wire popcount32_y9gs_core_056;
  wire popcount32_y9gs_core_057;
  wire popcount32_y9gs_core_060;
  wire popcount32_y9gs_core_063;
  wire popcount32_y9gs_core_065;
  wire popcount32_y9gs_core_066;
  wire popcount32_y9gs_core_067;
  wire popcount32_y9gs_core_069;
  wire popcount32_y9gs_core_070;
  wire popcount32_y9gs_core_071;
  wire popcount32_y9gs_core_072;
  wire popcount32_y9gs_core_076;
  wire popcount32_y9gs_core_077;
  wire popcount32_y9gs_core_078;
  wire popcount32_y9gs_core_079;
  wire popcount32_y9gs_core_080;
  wire popcount32_y9gs_core_083;
  wire popcount32_y9gs_core_085;
  wire popcount32_y9gs_core_086;
  wire popcount32_y9gs_core_087;
  wire popcount32_y9gs_core_090;
  wire popcount32_y9gs_core_091;
  wire popcount32_y9gs_core_092;
  wire popcount32_y9gs_core_093;
  wire popcount32_y9gs_core_095;
  wire popcount32_y9gs_core_097;
  wire popcount32_y9gs_core_098;
  wire popcount32_y9gs_core_099;
  wire popcount32_y9gs_core_100;
  wire popcount32_y9gs_core_101;
  wire popcount32_y9gs_core_103;
  wire popcount32_y9gs_core_106;
  wire popcount32_y9gs_core_107_not;
  wire popcount32_y9gs_core_108;
  wire popcount32_y9gs_core_109;
  wire popcount32_y9gs_core_110;
  wire popcount32_y9gs_core_111;
  wire popcount32_y9gs_core_112;
  wire popcount32_y9gs_core_114;
  wire popcount32_y9gs_core_115;
  wire popcount32_y9gs_core_116;
  wire popcount32_y9gs_core_118;
  wire popcount32_y9gs_core_120;
  wire popcount32_y9gs_core_121;
  wire popcount32_y9gs_core_122;
  wire popcount32_y9gs_core_124;
  wire popcount32_y9gs_core_127;
  wire popcount32_y9gs_core_129;
  wire popcount32_y9gs_core_131;
  wire popcount32_y9gs_core_134;
  wire popcount32_y9gs_core_135;
  wire popcount32_y9gs_core_138;
  wire popcount32_y9gs_core_139;
  wire popcount32_y9gs_core_140;
  wire popcount32_y9gs_core_141;
  wire popcount32_y9gs_core_142;
  wire popcount32_y9gs_core_143;
  wire popcount32_y9gs_core_144;
  wire popcount32_y9gs_core_145;
  wire popcount32_y9gs_core_146_not;
  wire popcount32_y9gs_core_148;
  wire popcount32_y9gs_core_150;
  wire popcount32_y9gs_core_151;
  wire popcount32_y9gs_core_152;
  wire popcount32_y9gs_core_157;
  wire popcount32_y9gs_core_159;
  wire popcount32_y9gs_core_160;
  wire popcount32_y9gs_core_162;
  wire popcount32_y9gs_core_163;
  wire popcount32_y9gs_core_165;
  wire popcount32_y9gs_core_168;
  wire popcount32_y9gs_core_169;
  wire popcount32_y9gs_core_172;
  wire popcount32_y9gs_core_173_not;
  wire popcount32_y9gs_core_174;
  wire popcount32_y9gs_core_175;
  wire popcount32_y9gs_core_176;
  wire popcount32_y9gs_core_177;
  wire popcount32_y9gs_core_179;
  wire popcount32_y9gs_core_180;
  wire popcount32_y9gs_core_185;
  wire popcount32_y9gs_core_186;
  wire popcount32_y9gs_core_187;
  wire popcount32_y9gs_core_188;
  wire popcount32_y9gs_core_190;
  wire popcount32_y9gs_core_193;
  wire popcount32_y9gs_core_194;
  wire popcount32_y9gs_core_195;
  wire popcount32_y9gs_core_198;
  wire popcount32_y9gs_core_202;
  wire popcount32_y9gs_core_204;
  wire popcount32_y9gs_core_210;
  wire popcount32_y9gs_core_211;
  wire popcount32_y9gs_core_212;
  wire popcount32_y9gs_core_213;
  wire popcount32_y9gs_core_214_not;
  wire popcount32_y9gs_core_217;
  wire popcount32_y9gs_core_219;
  wire popcount32_y9gs_core_220;
  wire popcount32_y9gs_core_221;
  wire popcount32_y9gs_core_222;
  wire popcount32_y9gs_core_223;
  wire popcount32_y9gs_core_224;
  wire popcount32_y9gs_core_225_not;

  assign popcount32_y9gs_core_034 = input_a[11] ^ input_a[0];
  assign popcount32_y9gs_core_035 = ~input_a[25];
  assign popcount32_y9gs_core_037 = input_a[17] | input_a[7];
  assign popcount32_y9gs_core_038 = ~(input_a[18] ^ input_a[9]);
  assign popcount32_y9gs_core_039 = ~input_a[14];
  assign popcount32_y9gs_core_040 = input_a[28] | input_a[23];
  assign popcount32_y9gs_core_043 = ~(input_a[0] | input_a[18]);
  assign popcount32_y9gs_core_045_not = ~input_a[11];
  assign popcount32_y9gs_core_046_not = ~input_a[19];
  assign popcount32_y9gs_core_048 = ~(input_a[12] ^ input_a[30]);
  assign popcount32_y9gs_core_050 = ~input_a[11];
  assign popcount32_y9gs_core_051 = ~(input_a[14] & input_a[18]);
  assign popcount32_y9gs_core_052 = ~(input_a[8] ^ input_a[24]);
  assign popcount32_y9gs_core_053 = input_a[11] & input_a[26];
  assign popcount32_y9gs_core_054 = ~(input_a[3] ^ input_a[11]);
  assign popcount32_y9gs_core_055 = input_a[2] & input_a[14];
  assign popcount32_y9gs_core_056 = ~(input_a[9] | input_a[7]);
  assign popcount32_y9gs_core_057 = input_a[19] ^ input_a[14];
  assign popcount32_y9gs_core_060 = input_a[8] | input_a[17];
  assign popcount32_y9gs_core_063 = input_a[12] | input_a[25];
  assign popcount32_y9gs_core_065 = input_a[6] ^ input_a[21];
  assign popcount32_y9gs_core_066 = input_a[14] | input_a[15];
  assign popcount32_y9gs_core_067 = input_a[4] & input_a[6];
  assign popcount32_y9gs_core_069 = ~(input_a[22] & input_a[30]);
  assign popcount32_y9gs_core_070 = input_a[21] ^ input_a[25];
  assign popcount32_y9gs_core_071 = ~(input_a[2] ^ input_a[11]);
  assign popcount32_y9gs_core_072 = input_a[31] & input_a[13];
  assign popcount32_y9gs_core_076 = ~(input_a[8] & input_a[31]);
  assign popcount32_y9gs_core_077 = input_a[31] ^ input_a[19];
  assign popcount32_y9gs_core_078 = input_a[1] | input_a[25];
  assign popcount32_y9gs_core_079 = input_a[24] & input_a[19];
  assign popcount32_y9gs_core_080 = input_a[3] ^ input_a[0];
  assign popcount32_y9gs_core_083 = input_a[8] ^ input_a[25];
  assign popcount32_y9gs_core_085 = input_a[14] | input_a[27];
  assign popcount32_y9gs_core_086 = input_a[8] ^ input_a[29];
  assign popcount32_y9gs_core_087 = input_a[10] ^ input_a[13];
  assign popcount32_y9gs_core_090 = input_a[22] | input_a[3];
  assign popcount32_y9gs_core_091 = input_a[0] | input_a[30];
  assign popcount32_y9gs_core_092 = ~input_a[1];
  assign popcount32_y9gs_core_093 = input_a[15] ^ input_a[20];
  assign popcount32_y9gs_core_095 = ~(input_a[23] ^ input_a[0]);
  assign popcount32_y9gs_core_097 = ~(input_a[12] & input_a[6]);
  assign popcount32_y9gs_core_098 = ~(input_a[10] & input_a[31]);
  assign popcount32_y9gs_core_099 = ~(input_a[17] | input_a[23]);
  assign popcount32_y9gs_core_100 = input_a[15] & input_a[17];
  assign popcount32_y9gs_core_101 = input_a[1] ^ input_a[13];
  assign popcount32_y9gs_core_103 = input_a[11] & input_a[27];
  assign popcount32_y9gs_core_106 = ~(input_a[8] & input_a[0]);
  assign popcount32_y9gs_core_107_not = ~input_a[12];
  assign popcount32_y9gs_core_108 = input_a[8] ^ input_a[15];
  assign popcount32_y9gs_core_109 = input_a[2] & input_a[25];
  assign popcount32_y9gs_core_110 = input_a[24] & input_a[18];
  assign popcount32_y9gs_core_111 = input_a[15] & input_a[29];
  assign popcount32_y9gs_core_112 = ~(input_a[30] & input_a[8]);
  assign popcount32_y9gs_core_114 = ~(input_a[24] ^ input_a[20]);
  assign popcount32_y9gs_core_115 = input_a[24] ^ input_a[20];
  assign popcount32_y9gs_core_116 = input_a[20] ^ input_a[21];
  assign popcount32_y9gs_core_118 = input_a[18] & input_a[23];
  assign popcount32_y9gs_core_120 = ~(input_a[30] | input_a[27]);
  assign popcount32_y9gs_core_121 = ~input_a[26];
  assign popcount32_y9gs_core_122 = ~input_a[7];
  assign popcount32_y9gs_core_124 = input_a[10] | input_a[7];
  assign popcount32_y9gs_core_127 = input_a[5] | input_a[13];
  assign popcount32_y9gs_core_129 = input_a[19] ^ input_a[22];
  assign popcount32_y9gs_core_131 = ~(input_a[31] & input_a[0]);
  assign popcount32_y9gs_core_134 = input_a[27] & input_a[2];
  assign popcount32_y9gs_core_135 = ~(input_a[1] ^ input_a[23]);
  assign popcount32_y9gs_core_138 = ~(input_a[1] | input_a[18]);
  assign popcount32_y9gs_core_139 = ~(input_a[28] | input_a[20]);
  assign popcount32_y9gs_core_140 = ~(input_a[25] | input_a[8]);
  assign popcount32_y9gs_core_141 = input_a[10] & input_a[9];
  assign popcount32_y9gs_core_142 = ~(input_a[27] ^ input_a[13]);
  assign popcount32_y9gs_core_143 = ~input_a[18];
  assign popcount32_y9gs_core_144 = input_a[20] ^ input_a[4];
  assign popcount32_y9gs_core_145 = ~(input_a[13] | input_a[16]);
  assign popcount32_y9gs_core_146_not = ~input_a[0];
  assign popcount32_y9gs_core_148 = input_a[11] & input_a[31];
  assign popcount32_y9gs_core_150 = ~input_a[21];
  assign popcount32_y9gs_core_151 = ~(input_a[8] ^ input_a[13]);
  assign popcount32_y9gs_core_152 = ~(input_a[24] & input_a[15]);
  assign popcount32_y9gs_core_157 = ~(input_a[19] & input_a[23]);
  assign popcount32_y9gs_core_159 = input_a[17] & input_a[8];
  assign popcount32_y9gs_core_160 = ~(input_a[17] & input_a[10]);
  assign popcount32_y9gs_core_162 = ~input_a[22];
  assign popcount32_y9gs_core_163 = ~input_a[10];
  assign popcount32_y9gs_core_165 = input_a[10] ^ input_a[18];
  assign popcount32_y9gs_core_168 = ~(input_a[24] & input_a[5]);
  assign popcount32_y9gs_core_169 = ~(input_a[14] ^ input_a[20]);
  assign popcount32_y9gs_core_172 = input_a[6] ^ input_a[29];
  assign popcount32_y9gs_core_173_not = ~input_a[27];
  assign popcount32_y9gs_core_174 = ~(input_a[25] ^ input_a[22]);
  assign popcount32_y9gs_core_175 = input_a[7] | input_a[8];
  assign popcount32_y9gs_core_176 = input_a[26] | input_a[6];
  assign popcount32_y9gs_core_177 = ~(input_a[3] ^ input_a[25]);
  assign popcount32_y9gs_core_179 = ~(input_a[1] ^ input_a[8]);
  assign popcount32_y9gs_core_180 = ~(input_a[15] | input_a[0]);
  assign popcount32_y9gs_core_185 = ~(input_a[8] ^ input_a[27]);
  assign popcount32_y9gs_core_186 = input_a[14] ^ input_a[9];
  assign popcount32_y9gs_core_187 = input_a[27] ^ input_a[29];
  assign popcount32_y9gs_core_188 = input_a[20] | input_a[25];
  assign popcount32_y9gs_core_190 = ~input_a[14];
  assign popcount32_y9gs_core_193 = ~(input_a[6] & input_a[9]);
  assign popcount32_y9gs_core_194 = ~(input_a[29] | input_a[18]);
  assign popcount32_y9gs_core_195 = input_a[19] ^ input_a[4];
  assign popcount32_y9gs_core_198 = ~input_a[8];
  assign popcount32_y9gs_core_202 = input_a[7] ^ input_a[21];
  assign popcount32_y9gs_core_204 = ~(input_a[29] ^ input_a[7]);
  assign popcount32_y9gs_core_210 = ~input_a[0];
  assign popcount32_y9gs_core_211 = input_a[3] | input_a[7];
  assign popcount32_y9gs_core_212 = input_a[22] | input_a[1];
  assign popcount32_y9gs_core_213 = input_a[8] ^ input_a[9];
  assign popcount32_y9gs_core_214_not = ~input_a[21];
  assign popcount32_y9gs_core_217 = input_a[9] ^ input_a[0];
  assign popcount32_y9gs_core_219 = ~(input_a[8] & input_a[31]);
  assign popcount32_y9gs_core_220 = input_a[31] ^ input_a[12];
  assign popcount32_y9gs_core_221 = ~input_a[4];
  assign popcount32_y9gs_core_222 = ~(input_a[29] & input_a[12]);
  assign popcount32_y9gs_core_223 = input_a[2] ^ input_a[28];
  assign popcount32_y9gs_core_224 = ~input_a[26];
  assign popcount32_y9gs_core_225_not = ~input_a[3];

  assign popcount32_y9gs_out[0] = 1'b1;
  assign popcount32_y9gs_out[1] = 1'b1;
  assign popcount32_y9gs_out[2] = input_a[3];
  assign popcount32_y9gs_out[3] = 1'b0;
  assign popcount32_y9gs_out[4] = 1'b0;
  assign popcount32_y9gs_out[5] = input_a[11];
endmodule