// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.59666
// WCE=19.0
// EP=0.962691%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_yfl4(input [28:0] input_a, output [4:0] popcount29_yfl4_out);
  wire popcount29_yfl4_core_031;
  wire popcount29_yfl4_core_034;
  wire popcount29_yfl4_core_035;
  wire popcount29_yfl4_core_037;
  wire popcount29_yfl4_core_038;
  wire popcount29_yfl4_core_042;
  wire popcount29_yfl4_core_043;
  wire popcount29_yfl4_core_044;
  wire popcount29_yfl4_core_047;
  wire popcount29_yfl4_core_048;
  wire popcount29_yfl4_core_049;
  wire popcount29_yfl4_core_051;
  wire popcount29_yfl4_core_052;
  wire popcount29_yfl4_core_054;
  wire popcount29_yfl4_core_055;
  wire popcount29_yfl4_core_056;
  wire popcount29_yfl4_core_057;
  wire popcount29_yfl4_core_059;
  wire popcount29_yfl4_core_060;
  wire popcount29_yfl4_core_061;
  wire popcount29_yfl4_core_062;
  wire popcount29_yfl4_core_063;
  wire popcount29_yfl4_core_064;
  wire popcount29_yfl4_core_065;
  wire popcount29_yfl4_core_067;
  wire popcount29_yfl4_core_068;
  wire popcount29_yfl4_core_072;
  wire popcount29_yfl4_core_074;
  wire popcount29_yfl4_core_076;
  wire popcount29_yfl4_core_079;
  wire popcount29_yfl4_core_081;
  wire popcount29_yfl4_core_082;
  wire popcount29_yfl4_core_084;
  wire popcount29_yfl4_core_085;
  wire popcount29_yfl4_core_086;
  wire popcount29_yfl4_core_087;
  wire popcount29_yfl4_core_088;
  wire popcount29_yfl4_core_089;
  wire popcount29_yfl4_core_090;
  wire popcount29_yfl4_core_091;
  wire popcount29_yfl4_core_095;
  wire popcount29_yfl4_core_097;
  wire popcount29_yfl4_core_099;
  wire popcount29_yfl4_core_101;
  wire popcount29_yfl4_core_102;
  wire popcount29_yfl4_core_103;
  wire popcount29_yfl4_core_104;
  wire popcount29_yfl4_core_107;
  wire popcount29_yfl4_core_108;
  wire popcount29_yfl4_core_110;
  wire popcount29_yfl4_core_112;
  wire popcount29_yfl4_core_115_not;
  wire popcount29_yfl4_core_117;
  wire popcount29_yfl4_core_119;
  wire popcount29_yfl4_core_121;
  wire popcount29_yfl4_core_122;
  wire popcount29_yfl4_core_123;
  wire popcount29_yfl4_core_124_not;
  wire popcount29_yfl4_core_125;
  wire popcount29_yfl4_core_126;
  wire popcount29_yfl4_core_129;
  wire popcount29_yfl4_core_130;
  wire popcount29_yfl4_core_132;
  wire popcount29_yfl4_core_133;
  wire popcount29_yfl4_core_134;
  wire popcount29_yfl4_core_136;
  wire popcount29_yfl4_core_137;
  wire popcount29_yfl4_core_138;
  wire popcount29_yfl4_core_139;
  wire popcount29_yfl4_core_142;
  wire popcount29_yfl4_core_146;
  wire popcount29_yfl4_core_147;
  wire popcount29_yfl4_core_153;
  wire popcount29_yfl4_core_154;
  wire popcount29_yfl4_core_155_not;
  wire popcount29_yfl4_core_157;
  wire popcount29_yfl4_core_158;
  wire popcount29_yfl4_core_159;
  wire popcount29_yfl4_core_160;
  wire popcount29_yfl4_core_161;
  wire popcount29_yfl4_core_162;
  wire popcount29_yfl4_core_163;
  wire popcount29_yfl4_core_164;
  wire popcount29_yfl4_core_166;
  wire popcount29_yfl4_core_169;
  wire popcount29_yfl4_core_170;
  wire popcount29_yfl4_core_174;
  wire popcount29_yfl4_core_175;
  wire popcount29_yfl4_core_177;
  wire popcount29_yfl4_core_178;
  wire popcount29_yfl4_core_181;
  wire popcount29_yfl4_core_183;
  wire popcount29_yfl4_core_184;
  wire popcount29_yfl4_core_185;
  wire popcount29_yfl4_core_186;
  wire popcount29_yfl4_core_187;
  wire popcount29_yfl4_core_188;
  wire popcount29_yfl4_core_189;
  wire popcount29_yfl4_core_191;
  wire popcount29_yfl4_core_193;
  wire popcount29_yfl4_core_194;
  wire popcount29_yfl4_core_195;
  wire popcount29_yfl4_core_196;
  wire popcount29_yfl4_core_197;
  wire popcount29_yfl4_core_198;
  wire popcount29_yfl4_core_199;
  wire popcount29_yfl4_core_200;
  wire popcount29_yfl4_core_204;
  wire popcount29_yfl4_core_206;

  assign popcount29_yfl4_core_031 = ~(input_a[27] | input_a[7]);
  assign popcount29_yfl4_core_034 = ~(input_a[12] & input_a[7]);
  assign popcount29_yfl4_core_035 = ~(input_a[27] | input_a[23]);
  assign popcount29_yfl4_core_037 = input_a[21] & input_a[0];
  assign popcount29_yfl4_core_038 = ~(input_a[27] | input_a[0]);
  assign popcount29_yfl4_core_042 = input_a[0] ^ input_a[24];
  assign popcount29_yfl4_core_043 = ~(input_a[22] ^ input_a[21]);
  assign popcount29_yfl4_core_044 = ~(input_a[23] & input_a[19]);
  assign popcount29_yfl4_core_047 = ~(input_a[11] ^ input_a[15]);
  assign popcount29_yfl4_core_048 = ~(input_a[1] & input_a[23]);
  assign popcount29_yfl4_core_049 = ~(input_a[20] ^ input_a[5]);
  assign popcount29_yfl4_core_051 = input_a[28] | input_a[5];
  assign popcount29_yfl4_core_052 = ~(input_a[4] & input_a[16]);
  assign popcount29_yfl4_core_054 = ~(input_a[28] & input_a[17]);
  assign popcount29_yfl4_core_055 = ~input_a[17];
  assign popcount29_yfl4_core_056 = input_a[22] ^ input_a[21];
  assign popcount29_yfl4_core_057 = ~(input_a[5] ^ input_a[20]);
  assign popcount29_yfl4_core_059 = ~input_a[21];
  assign popcount29_yfl4_core_060 = input_a[14] ^ input_a[3];
  assign popcount29_yfl4_core_061 = input_a[2] ^ input_a[14];
  assign popcount29_yfl4_core_062 = ~(input_a[9] | input_a[5]);
  assign popcount29_yfl4_core_063 = input_a[24] ^ input_a[18];
  assign popcount29_yfl4_core_064 = ~(input_a[18] ^ input_a[28]);
  assign popcount29_yfl4_core_065 = ~(input_a[8] | input_a[17]);
  assign popcount29_yfl4_core_067 = input_a[7] & input_a[28];
  assign popcount29_yfl4_core_068 = ~(input_a[18] & input_a[0]);
  assign popcount29_yfl4_core_072 = input_a[7] & input_a[26];
  assign popcount29_yfl4_core_074 = ~(input_a[25] & input_a[8]);
  assign popcount29_yfl4_core_076 = ~input_a[7];
  assign popcount29_yfl4_core_079 = input_a[12] & input_a[3];
  assign popcount29_yfl4_core_081 = input_a[23] & input_a[13];
  assign popcount29_yfl4_core_082 = ~(input_a[6] & input_a[16]);
  assign popcount29_yfl4_core_084 = ~(input_a[10] ^ input_a[19]);
  assign popcount29_yfl4_core_085 = input_a[11] & input_a[11];
  assign popcount29_yfl4_core_086 = input_a[22] & input_a[8];
  assign popcount29_yfl4_core_087 = input_a[14] | input_a[28];
  assign popcount29_yfl4_core_088 = input_a[4] ^ input_a[24];
  assign popcount29_yfl4_core_089 = input_a[17] ^ input_a[1];
  assign popcount29_yfl4_core_090 = input_a[20] | input_a[20];
  assign popcount29_yfl4_core_091 = ~(input_a[25] ^ input_a[7]);
  assign popcount29_yfl4_core_095 = ~(input_a[4] & input_a[23]);
  assign popcount29_yfl4_core_097 = ~(input_a[22] ^ input_a[4]);
  assign popcount29_yfl4_core_099 = input_a[3] & input_a[2];
  assign popcount29_yfl4_core_101 = ~input_a[11];
  assign popcount29_yfl4_core_102 = ~input_a[11];
  assign popcount29_yfl4_core_103 = input_a[12] | input_a[9];
  assign popcount29_yfl4_core_104 = input_a[11] | input_a[5];
  assign popcount29_yfl4_core_107 = input_a[28] | input_a[14];
  assign popcount29_yfl4_core_108 = ~(input_a[8] ^ input_a[4]);
  assign popcount29_yfl4_core_110 = ~(input_a[1] | input_a[14]);
  assign popcount29_yfl4_core_112 = input_a[26] & input_a[26];
  assign popcount29_yfl4_core_115_not = ~input_a[4];
  assign popcount29_yfl4_core_117 = ~(input_a[23] & input_a[25]);
  assign popcount29_yfl4_core_119 = ~(input_a[24] & input_a[19]);
  assign popcount29_yfl4_core_121 = input_a[25] & input_a[14];
  assign popcount29_yfl4_core_122 = ~(input_a[20] | input_a[16]);
  assign popcount29_yfl4_core_123 = input_a[4] ^ input_a[20];
  assign popcount29_yfl4_core_124_not = ~input_a[28];
  assign popcount29_yfl4_core_125 = input_a[3] ^ input_a[13];
  assign popcount29_yfl4_core_126 = ~(input_a[0] & input_a[10]);
  assign popcount29_yfl4_core_129 = ~(input_a[7] & input_a[23]);
  assign popcount29_yfl4_core_130 = input_a[15] & input_a[9];
  assign popcount29_yfl4_core_132 = ~input_a[28];
  assign popcount29_yfl4_core_133 = input_a[21] | input_a[28];
  assign popcount29_yfl4_core_134 = ~(input_a[10] | input_a[7]);
  assign popcount29_yfl4_core_136 = input_a[10] & input_a[19];
  assign popcount29_yfl4_core_137 = input_a[12] & input_a[28];
  assign popcount29_yfl4_core_138 = input_a[26] & input_a[25];
  assign popcount29_yfl4_core_139 = input_a[23] | input_a[25];
  assign popcount29_yfl4_core_142 = ~(input_a[19] ^ input_a[2]);
  assign popcount29_yfl4_core_146 = ~(input_a[21] & input_a[21]);
  assign popcount29_yfl4_core_147 = ~(input_a[8] | input_a[4]);
  assign popcount29_yfl4_core_153 = ~(input_a[21] | input_a[14]);
  assign popcount29_yfl4_core_154 = input_a[19] ^ input_a[5];
  assign popcount29_yfl4_core_155_not = ~input_a[18];
  assign popcount29_yfl4_core_157 = ~(input_a[19] | input_a[3]);
  assign popcount29_yfl4_core_158 = input_a[9] ^ input_a[5];
  assign popcount29_yfl4_core_159 = input_a[24] ^ input_a[5];
  assign popcount29_yfl4_core_160 = input_a[26] | input_a[27];
  assign popcount29_yfl4_core_161 = ~(input_a[27] & input_a[15]);
  assign popcount29_yfl4_core_162 = ~input_a[14];
  assign popcount29_yfl4_core_163 = ~input_a[8];
  assign popcount29_yfl4_core_164 = ~(input_a[9] ^ input_a[27]);
  assign popcount29_yfl4_core_166 = ~(input_a[13] ^ input_a[18]);
  assign popcount29_yfl4_core_169 = input_a[11] & input_a[6];
  assign popcount29_yfl4_core_170 = input_a[13] & input_a[7];
  assign popcount29_yfl4_core_174 = input_a[24] | input_a[19];
  assign popcount29_yfl4_core_175 = input_a[25] | input_a[10];
  assign popcount29_yfl4_core_177 = input_a[6] | input_a[26];
  assign popcount29_yfl4_core_178 = input_a[20] ^ input_a[25];
  assign popcount29_yfl4_core_181 = ~(input_a[8] | input_a[7]);
  assign popcount29_yfl4_core_183 = input_a[12] & input_a[7];
  assign popcount29_yfl4_core_184 = ~(input_a[0] | input_a[20]);
  assign popcount29_yfl4_core_185 = ~(input_a[6] & input_a[17]);
  assign popcount29_yfl4_core_186 = input_a[17] | input_a[26];
  assign popcount29_yfl4_core_187 = ~(input_a[4] & input_a[2]);
  assign popcount29_yfl4_core_188 = input_a[1] & input_a[8];
  assign popcount29_yfl4_core_189 = ~(input_a[1] | input_a[27]);
  assign popcount29_yfl4_core_191 = ~(input_a[3] & input_a[2]);
  assign popcount29_yfl4_core_193 = ~input_a[16];
  assign popcount29_yfl4_core_194 = ~(input_a[25] & input_a[27]);
  assign popcount29_yfl4_core_195 = input_a[13] | input_a[19];
  assign popcount29_yfl4_core_196 = input_a[21] & input_a[10];
  assign popcount29_yfl4_core_197 = input_a[11] & input_a[19];
  assign popcount29_yfl4_core_198 = ~input_a[26];
  assign popcount29_yfl4_core_199 = input_a[25] ^ input_a[8];
  assign popcount29_yfl4_core_200 = ~input_a[0];
  assign popcount29_yfl4_core_204 = input_a[1] | input_a[8];
  assign popcount29_yfl4_core_206 = ~(input_a[19] ^ input_a[4]);

  assign popcount29_yfl4_out[0] = 1'b1;
  assign popcount29_yfl4_out[1] = input_a[10];
  assign popcount29_yfl4_out[2] = 1'b0;
  assign popcount29_yfl4_out[3] = 1'b1;
  assign popcount29_yfl4_out[4] = 1'b0;
endmodule