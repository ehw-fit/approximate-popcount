// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.13539
// WCE=17.0
// EP=0.926298%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_rprm(input [20:0] input_a, output [4:0] popcount21_rprm_out);
  wire popcount21_rprm_core_023;
  wire popcount21_rprm_core_025;
  wire popcount21_rprm_core_026;
  wire popcount21_rprm_core_027_not;
  wire popcount21_rprm_core_029;
  wire popcount21_rprm_core_030;
  wire popcount21_rprm_core_031;
  wire popcount21_rprm_core_032;
  wire popcount21_rprm_core_034;
  wire popcount21_rprm_core_035;
  wire popcount21_rprm_core_036;
  wire popcount21_rprm_core_037;
  wire popcount21_rprm_core_038;
  wire popcount21_rprm_core_039;
  wire popcount21_rprm_core_044;
  wire popcount21_rprm_core_045;
  wire popcount21_rprm_core_047;
  wire popcount21_rprm_core_048;
  wire popcount21_rprm_core_049;
  wire popcount21_rprm_core_051;
  wire popcount21_rprm_core_052;
  wire popcount21_rprm_core_057;
  wire popcount21_rprm_core_059;
  wire popcount21_rprm_core_061;
  wire popcount21_rprm_core_062;
  wire popcount21_rprm_core_065;
  wire popcount21_rprm_core_066;
  wire popcount21_rprm_core_067;
  wire popcount21_rprm_core_068;
  wire popcount21_rprm_core_069;
  wire popcount21_rprm_core_072;
  wire popcount21_rprm_core_073;
  wire popcount21_rprm_core_074;
  wire popcount21_rprm_core_076;
  wire popcount21_rprm_core_078;
  wire popcount21_rprm_core_080;
  wire popcount21_rprm_core_081;
  wire popcount21_rprm_core_082;
  wire popcount21_rprm_core_086;
  wire popcount21_rprm_core_089;
  wire popcount21_rprm_core_091;
  wire popcount21_rprm_core_093;
  wire popcount21_rprm_core_094;
  wire popcount21_rprm_core_095_not;
  wire popcount21_rprm_core_098;
  wire popcount21_rprm_core_099;
  wire popcount21_rprm_core_100;
  wire popcount21_rprm_core_102_not;
  wire popcount21_rprm_core_104;
  wire popcount21_rprm_core_105;
  wire popcount21_rprm_core_110;
  wire popcount21_rprm_core_111;
  wire popcount21_rprm_core_112;
  wire popcount21_rprm_core_113;
  wire popcount21_rprm_core_114;
  wire popcount21_rprm_core_115;
  wire popcount21_rprm_core_116;
  wire popcount21_rprm_core_117;
  wire popcount21_rprm_core_118;
  wire popcount21_rprm_core_119;
  wire popcount21_rprm_core_121;
  wire popcount21_rprm_core_122;
  wire popcount21_rprm_core_129;
  wire popcount21_rprm_core_130;
  wire popcount21_rprm_core_132;
  wire popcount21_rprm_core_133;
  wire popcount21_rprm_core_135;
  wire popcount21_rprm_core_136;
  wire popcount21_rprm_core_137;
  wire popcount21_rprm_core_138;
  wire popcount21_rprm_core_140;
  wire popcount21_rprm_core_142;
  wire popcount21_rprm_core_144;
  wire popcount21_rprm_core_145;
  wire popcount21_rprm_core_146;
  wire popcount21_rprm_core_147;
  wire popcount21_rprm_core_150;
  wire popcount21_rprm_core_151_not;
  wire popcount21_rprm_core_152;
  wire popcount21_rprm_core_153;

  assign popcount21_rprm_core_023 = ~(input_a[2] ^ input_a[7]);
  assign popcount21_rprm_core_025 = input_a[16] ^ input_a[4];
  assign popcount21_rprm_core_026 = input_a[19] & input_a[17];
  assign popcount21_rprm_core_027_not = ~input_a[6];
  assign popcount21_rprm_core_029 = ~(input_a[1] & input_a[16]);
  assign popcount21_rprm_core_030 = input_a[7] & input_a[9];
  assign popcount21_rprm_core_031 = ~input_a[20];
  assign popcount21_rprm_core_032 = input_a[6] & input_a[0];
  assign popcount21_rprm_core_034 = ~(input_a[13] | input_a[10]);
  assign popcount21_rprm_core_035 = ~(input_a[17] | input_a[7]);
  assign popcount21_rprm_core_036 = ~(input_a[16] ^ input_a[17]);
  assign popcount21_rprm_core_037 = input_a[17] | input_a[3];
  assign popcount21_rprm_core_038 = ~(input_a[9] | input_a[18]);
  assign popcount21_rprm_core_039 = input_a[11] ^ input_a[8];
  assign popcount21_rprm_core_044 = input_a[14] & input_a[10];
  assign popcount21_rprm_core_045 = ~(input_a[20] | input_a[0]);
  assign popcount21_rprm_core_047 = ~(input_a[18] | input_a[4]);
  assign popcount21_rprm_core_048 = input_a[2] ^ input_a[18];
  assign popcount21_rprm_core_049 = ~input_a[8];
  assign popcount21_rprm_core_051 = input_a[16] & input_a[15];
  assign popcount21_rprm_core_052 = ~(input_a[6] & input_a[15]);
  assign popcount21_rprm_core_057 = ~(input_a[16] ^ input_a[8]);
  assign popcount21_rprm_core_059 = input_a[12] | input_a[14];
  assign popcount21_rprm_core_061 = input_a[16] & input_a[5];
  assign popcount21_rprm_core_062 = ~(input_a[11] & input_a[16]);
  assign popcount21_rprm_core_065 = ~input_a[16];
  assign popcount21_rprm_core_066 = ~(input_a[12] | input_a[17]);
  assign popcount21_rprm_core_067 = ~input_a[16];
  assign popcount21_rprm_core_068 = ~input_a[12];
  assign popcount21_rprm_core_069 = ~(input_a[13] | input_a[2]);
  assign popcount21_rprm_core_072 = ~input_a[6];
  assign popcount21_rprm_core_073 = input_a[14] ^ input_a[8];
  assign popcount21_rprm_core_074 = ~input_a[3];
  assign popcount21_rprm_core_076 = input_a[18] & input_a[7];
  assign popcount21_rprm_core_078 = ~input_a[9];
  assign popcount21_rprm_core_080 = ~(input_a[12] & input_a[10]);
  assign popcount21_rprm_core_081 = input_a[9] & input_a[16];
  assign popcount21_rprm_core_082 = ~(input_a[4] | input_a[14]);
  assign popcount21_rprm_core_086 = input_a[15] & input_a[11];
  assign popcount21_rprm_core_089 = ~(input_a[6] & input_a[4]);
  assign popcount21_rprm_core_091 = input_a[13] ^ input_a[17];
  assign popcount21_rprm_core_093 = ~(input_a[18] & input_a[0]);
  assign popcount21_rprm_core_094 = ~(input_a[13] & input_a[12]);
  assign popcount21_rprm_core_095_not = ~input_a[7];
  assign popcount21_rprm_core_098 = ~(input_a[8] | input_a[19]);
  assign popcount21_rprm_core_099 = input_a[19] | input_a[8];
  assign popcount21_rprm_core_100 = ~input_a[10];
  assign popcount21_rprm_core_102_not = ~input_a[17];
  assign popcount21_rprm_core_104 = ~(input_a[7] & input_a[9]);
  assign popcount21_rprm_core_105 = input_a[12] | input_a[10];
  assign popcount21_rprm_core_110 = input_a[14] ^ input_a[3];
  assign popcount21_rprm_core_111 = ~input_a[14];
  assign popcount21_rprm_core_112 = input_a[15] & input_a[19];
  assign popcount21_rprm_core_113 = ~(input_a[6] & input_a[16]);
  assign popcount21_rprm_core_114 = ~input_a[7];
  assign popcount21_rprm_core_115 = input_a[16] & input_a[19];
  assign popcount21_rprm_core_116 = ~input_a[2];
  assign popcount21_rprm_core_117 = ~(input_a[17] | input_a[0]);
  assign popcount21_rprm_core_118 = ~(input_a[14] ^ input_a[19]);
  assign popcount21_rprm_core_119 = input_a[20] & input_a[9];
  assign popcount21_rprm_core_121 = ~(input_a[1] | input_a[18]);
  assign popcount21_rprm_core_122 = input_a[10] & input_a[3];
  assign popcount21_rprm_core_129 = input_a[7] | input_a[4];
  assign popcount21_rprm_core_130 = input_a[9] | input_a[17];
  assign popcount21_rprm_core_132 = ~(input_a[12] & input_a[14]);
  assign popcount21_rprm_core_133 = ~(input_a[2] ^ input_a[11]);
  assign popcount21_rprm_core_135 = ~(input_a[15] & input_a[17]);
  assign popcount21_rprm_core_136 = input_a[14] & input_a[12];
  assign popcount21_rprm_core_137 = ~(input_a[11] | input_a[20]);
  assign popcount21_rprm_core_138 = ~(input_a[3] & input_a[17]);
  assign popcount21_rprm_core_140 = ~(input_a[6] & input_a[4]);
  assign popcount21_rprm_core_142 = ~(input_a[3] | input_a[18]);
  assign popcount21_rprm_core_144 = input_a[12] & input_a[6];
  assign popcount21_rprm_core_145 = ~(input_a[16] | input_a[10]);
  assign popcount21_rprm_core_146 = ~(input_a[2] | input_a[14]);
  assign popcount21_rprm_core_147 = input_a[5] & input_a[0];
  assign popcount21_rprm_core_150 = input_a[18] ^ input_a[12];
  assign popcount21_rprm_core_151_not = ~input_a[19];
  assign popcount21_rprm_core_152 = ~(input_a[12] | input_a[6]);
  assign popcount21_rprm_core_153 = ~(input_a[1] ^ input_a[20]);

  assign popcount21_rprm_out[0] = 1'b0;
  assign popcount21_rprm_out[1] = 1'b1;
  assign popcount21_rprm_out[2] = input_a[6];
  assign popcount21_rprm_out[3] = input_a[5];
  assign popcount21_rprm_out[4] = 1'b0;
endmodule