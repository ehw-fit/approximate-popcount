// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.47244
// WCE=33.0
// EP=0.904025%
// Printed PDK parameters:
//  Area=73475914.0
//  Delay=80990424.0
//  Power=3589500.0

module popcount35_kfnc(input [34:0] input_a, output [5:0] popcount35_kfnc_out);
  wire popcount35_kfnc_core_037;
  wire popcount35_kfnc_core_038;
  wire popcount35_kfnc_core_039;
  wire popcount35_kfnc_core_040;
  wire popcount35_kfnc_core_042;
  wire popcount35_kfnc_core_043;
  wire popcount35_kfnc_core_044;
  wire popcount35_kfnc_core_045;
  wire popcount35_kfnc_core_046;
  wire popcount35_kfnc_core_047;
  wire popcount35_kfnc_core_048;
  wire popcount35_kfnc_core_052;
  wire popcount35_kfnc_core_057;
  wire popcount35_kfnc_core_059_not;
  wire popcount35_kfnc_core_061;
  wire popcount35_kfnc_core_063;
  wire popcount35_kfnc_core_064;
  wire popcount35_kfnc_core_066_not;
  wire popcount35_kfnc_core_068;
  wire popcount35_kfnc_core_069;
  wire popcount35_kfnc_core_070;
  wire popcount35_kfnc_core_071;
  wire popcount35_kfnc_core_073;
  wire popcount35_kfnc_core_074;
  wire popcount35_kfnc_core_075;
  wire popcount35_kfnc_core_076;
  wire popcount35_kfnc_core_077;
  wire popcount35_kfnc_core_078;
  wire popcount35_kfnc_core_079;
  wire popcount35_kfnc_core_080;
  wire popcount35_kfnc_core_081;
  wire popcount35_kfnc_core_082;
  wire popcount35_kfnc_core_083;
  wire popcount35_kfnc_core_084;
  wire popcount35_kfnc_core_086;
  wire popcount35_kfnc_core_088;
  wire popcount35_kfnc_core_089;
  wire popcount35_kfnc_core_090;
  wire popcount35_kfnc_core_091;
  wire popcount35_kfnc_core_092;
  wire popcount35_kfnc_core_093;
  wire popcount35_kfnc_core_095;
  wire popcount35_kfnc_core_096;
  wire popcount35_kfnc_core_098;
  wire popcount35_kfnc_core_099;
  wire popcount35_kfnc_core_100;
  wire popcount35_kfnc_core_103;
  wire popcount35_kfnc_core_104;
  wire popcount35_kfnc_core_106;
  wire popcount35_kfnc_core_107;
  wire popcount35_kfnc_core_108;
  wire popcount35_kfnc_core_109;
  wire popcount35_kfnc_core_114;
  wire popcount35_kfnc_core_115;
  wire popcount35_kfnc_core_116;
  wire popcount35_kfnc_core_117;
  wire popcount35_kfnc_core_118;
  wire popcount35_kfnc_core_119;
  wire popcount35_kfnc_core_120;
  wire popcount35_kfnc_core_121;
  wire popcount35_kfnc_core_122;
  wire popcount35_kfnc_core_123;
  wire popcount35_kfnc_core_124;
  wire popcount35_kfnc_core_125;
  wire popcount35_kfnc_core_126;
  wire popcount35_kfnc_core_127;
  wire popcount35_kfnc_core_128;
  wire popcount35_kfnc_core_129;
  wire popcount35_kfnc_core_132;
  wire popcount35_kfnc_core_133;
  wire popcount35_kfnc_core_135;
  wire popcount35_kfnc_core_138;
  wire popcount35_kfnc_core_139;
  wire popcount35_kfnc_core_143;
  wire popcount35_kfnc_core_144;
  wire popcount35_kfnc_core_145;
  wire popcount35_kfnc_core_146;
  wire popcount35_kfnc_core_147;
  wire popcount35_kfnc_core_149;
  wire popcount35_kfnc_core_150;
  wire popcount35_kfnc_core_151;
  wire popcount35_kfnc_core_153;
  wire popcount35_kfnc_core_161;
  wire popcount35_kfnc_core_162_not;
  wire popcount35_kfnc_core_164;
  wire popcount35_kfnc_core_165;
  wire popcount35_kfnc_core_166;
  wire popcount35_kfnc_core_167;
  wire popcount35_kfnc_core_169;
  wire popcount35_kfnc_core_170;
  wire popcount35_kfnc_core_174;
  wire popcount35_kfnc_core_175;
  wire popcount35_kfnc_core_176;
  wire popcount35_kfnc_core_177;
  wire popcount35_kfnc_core_178;
  wire popcount35_kfnc_core_179;
  wire popcount35_kfnc_core_180;
  wire popcount35_kfnc_core_181;
  wire popcount35_kfnc_core_182;
  wire popcount35_kfnc_core_183;
  wire popcount35_kfnc_core_184;
  wire popcount35_kfnc_core_185;
  wire popcount35_kfnc_core_187;
  wire popcount35_kfnc_core_188;
  wire popcount35_kfnc_core_189;
  wire popcount35_kfnc_core_190;
  wire popcount35_kfnc_core_191;
  wire popcount35_kfnc_core_192;
  wire popcount35_kfnc_core_193;
  wire popcount35_kfnc_core_194;
  wire popcount35_kfnc_core_197;
  wire popcount35_kfnc_core_198;
  wire popcount35_kfnc_core_200;
  wire popcount35_kfnc_core_201;
  wire popcount35_kfnc_core_202;
  wire popcount35_kfnc_core_203;
  wire popcount35_kfnc_core_204;
  wire popcount35_kfnc_core_205;
  wire popcount35_kfnc_core_206;
  wire popcount35_kfnc_core_207;
  wire popcount35_kfnc_core_208;
  wire popcount35_kfnc_core_209;
  wire popcount35_kfnc_core_210;
  wire popcount35_kfnc_core_211;
  wire popcount35_kfnc_core_212;
  wire popcount35_kfnc_core_213;
  wire popcount35_kfnc_core_214;
  wire popcount35_kfnc_core_215;
  wire popcount35_kfnc_core_216;
  wire popcount35_kfnc_core_217;
  wire popcount35_kfnc_core_218;
  wire popcount35_kfnc_core_219;
  wire popcount35_kfnc_core_220;
  wire popcount35_kfnc_core_221;
  wire popcount35_kfnc_core_222;
  wire popcount35_kfnc_core_223;
  wire popcount35_kfnc_core_224;
  wire popcount35_kfnc_core_225;
  wire popcount35_kfnc_core_226;
  wire popcount35_kfnc_core_227;
  wire popcount35_kfnc_core_228;
  wire popcount35_kfnc_core_229;
  wire popcount35_kfnc_core_230;
  wire popcount35_kfnc_core_231;
  wire popcount35_kfnc_core_232;
  wire popcount35_kfnc_core_234;
  wire popcount35_kfnc_core_235;
  wire popcount35_kfnc_core_236;
  wire popcount35_kfnc_core_237;
  wire popcount35_kfnc_core_238;
  wire popcount35_kfnc_core_239;
  wire popcount35_kfnc_core_241;
  wire popcount35_kfnc_core_242;
  wire popcount35_kfnc_core_243;
  wire popcount35_kfnc_core_244;
  wire popcount35_kfnc_core_245;
  wire popcount35_kfnc_core_246;
  wire popcount35_kfnc_core_247;
  wire popcount35_kfnc_core_248;
  wire popcount35_kfnc_core_249;
  wire popcount35_kfnc_core_250;
  wire popcount35_kfnc_core_251;
  wire popcount35_kfnc_core_252;
  wire popcount35_kfnc_core_253;
  wire popcount35_kfnc_core_254;
  wire popcount35_kfnc_core_257;
  wire popcount35_kfnc_core_258;
  wire popcount35_kfnc_core_261_not;
  wire popcount35_kfnc_core_262;
  wire popcount35_kfnc_core_263;
  wire popcount35_kfnc_core_264;

  assign popcount35_kfnc_core_037 = input_a[0] ^ input_a[1];
  assign popcount35_kfnc_core_038 = input_a[0] & input_a[1];
  assign popcount35_kfnc_core_039 = input_a[2] ^ input_a[3];
  assign popcount35_kfnc_core_040 = input_a[2] & input_a[3];
  assign popcount35_kfnc_core_042 = popcount35_kfnc_core_037 & popcount35_kfnc_core_039;
  assign popcount35_kfnc_core_043 = popcount35_kfnc_core_038 ^ popcount35_kfnc_core_040;
  assign popcount35_kfnc_core_044 = popcount35_kfnc_core_038 & popcount35_kfnc_core_040;
  assign popcount35_kfnc_core_045 = ~popcount35_kfnc_core_043;
  assign popcount35_kfnc_core_046 = popcount35_kfnc_core_043 & popcount35_kfnc_core_042;
  assign popcount35_kfnc_core_047 = popcount35_kfnc_core_044 | popcount35_kfnc_core_046;
  assign popcount35_kfnc_core_048 = input_a[4] ^ input_a[5];
  assign popcount35_kfnc_core_052 = popcount35_kfnc_core_048 ^ input_a[10];
  assign popcount35_kfnc_core_057 = input_a[4] & input_a[26];
  assign popcount35_kfnc_core_059_not = ~popcount35_kfnc_core_052;
  assign popcount35_kfnc_core_061 = popcount35_kfnc_core_045 ^ input_a[14];
  assign popcount35_kfnc_core_063 = popcount35_kfnc_core_061 ^ popcount35_kfnc_core_052;
  assign popcount35_kfnc_core_064 = popcount35_kfnc_core_061 & popcount35_kfnc_core_052;
  assign popcount35_kfnc_core_066_not = ~popcount35_kfnc_core_047;
  assign popcount35_kfnc_core_068 = popcount35_kfnc_core_066_not ^ popcount35_kfnc_core_064;
  assign popcount35_kfnc_core_069 = popcount35_kfnc_core_066_not & popcount35_kfnc_core_064;
  assign popcount35_kfnc_core_070 = popcount35_kfnc_core_047 | popcount35_kfnc_core_069;
  assign popcount35_kfnc_core_071 = input_a[8] ^ input_a[9];
  assign popcount35_kfnc_core_073 = input_a[10] ^ input_a[11];
  assign popcount35_kfnc_core_074 = input_a[10] & input_a[11];
  assign popcount35_kfnc_core_075 = ~popcount35_kfnc_core_071;
  assign popcount35_kfnc_core_076 = input_a[13] & popcount35_kfnc_core_073;
  assign popcount35_kfnc_core_077 = input_a[8] ^ popcount35_kfnc_core_074;
  assign popcount35_kfnc_core_078 = input_a[8] & popcount35_kfnc_core_074;
  assign popcount35_kfnc_core_079 = popcount35_kfnc_core_077 ^ popcount35_kfnc_core_076;
  assign popcount35_kfnc_core_080 = popcount35_kfnc_core_077 & popcount35_kfnc_core_076;
  assign popcount35_kfnc_core_081 = popcount35_kfnc_core_078 | popcount35_kfnc_core_080;
  assign popcount35_kfnc_core_082 = ~(input_a[29] & input_a[6]);
  assign popcount35_kfnc_core_083 = input_a[21] & input_a[13];
  assign popcount35_kfnc_core_084 = input_a[24] ^ input_a[16];
  assign popcount35_kfnc_core_086 = input_a[14] & input_a[32];
  assign popcount35_kfnc_core_088 = ~(input_a[15] & input_a[2]);
  assign popcount35_kfnc_core_089 = input_a[15] & input_a[2];
  assign popcount35_kfnc_core_090 = input_a[17] ^ input_a[24];
  assign popcount35_kfnc_core_091 = popcount35_kfnc_core_082 & input_a[22];
  assign popcount35_kfnc_core_092 = ~(input_a[34] | popcount35_kfnc_core_088);
  assign popcount35_kfnc_core_093 = input_a[22] & popcount35_kfnc_core_088;
  assign popcount35_kfnc_core_095 = input_a[11] & input_a[31];
  assign popcount35_kfnc_core_096 = input_a[15] | popcount35_kfnc_core_095;
  assign popcount35_kfnc_core_098 = popcount35_kfnc_core_089 & popcount35_kfnc_core_096;
  assign popcount35_kfnc_core_099 = ~(popcount35_kfnc_core_075 & popcount35_kfnc_core_090);
  assign popcount35_kfnc_core_100 = popcount35_kfnc_core_075 & popcount35_kfnc_core_090;
  assign popcount35_kfnc_core_103 = popcount35_kfnc_core_079 ^ popcount35_kfnc_core_100;
  assign popcount35_kfnc_core_104 = popcount35_kfnc_core_079 & popcount35_kfnc_core_100;
  assign popcount35_kfnc_core_106 = popcount35_kfnc_core_081 ^ popcount35_kfnc_core_089;
  assign popcount35_kfnc_core_107 = popcount35_kfnc_core_081 & popcount35_kfnc_core_089;
  assign popcount35_kfnc_core_108 = popcount35_kfnc_core_106 ^ popcount35_kfnc_core_104;
  assign popcount35_kfnc_core_109 = popcount35_kfnc_core_106 & popcount35_kfnc_core_104;
  assign popcount35_kfnc_core_114 = popcount35_kfnc_core_059_not & popcount35_kfnc_core_099;
  assign popcount35_kfnc_core_115 = popcount35_kfnc_core_063 ^ popcount35_kfnc_core_103;
  assign popcount35_kfnc_core_116 = popcount35_kfnc_core_063 & popcount35_kfnc_core_103;
  assign popcount35_kfnc_core_117 = popcount35_kfnc_core_115 ^ popcount35_kfnc_core_114;
  assign popcount35_kfnc_core_118 = popcount35_kfnc_core_115 & popcount35_kfnc_core_114;
  assign popcount35_kfnc_core_119 = popcount35_kfnc_core_116 | popcount35_kfnc_core_118;
  assign popcount35_kfnc_core_120 = popcount35_kfnc_core_068 ^ popcount35_kfnc_core_108;
  assign popcount35_kfnc_core_121 = popcount35_kfnc_core_068 & popcount35_kfnc_core_108;
  assign popcount35_kfnc_core_122 = popcount35_kfnc_core_120 ^ popcount35_kfnc_core_119;
  assign popcount35_kfnc_core_123 = popcount35_kfnc_core_120 & popcount35_kfnc_core_119;
  assign popcount35_kfnc_core_124 = popcount35_kfnc_core_121 | popcount35_kfnc_core_123;
  assign popcount35_kfnc_core_125 = popcount35_kfnc_core_070 ^ popcount35_kfnc_core_098;
  assign popcount35_kfnc_core_126 = input_a[15] & input_a[16];
  assign popcount35_kfnc_core_127 = popcount35_kfnc_core_125 ^ popcount35_kfnc_core_124;
  assign popcount35_kfnc_core_128 = input_a[25] & popcount35_kfnc_core_124;
  assign popcount35_kfnc_core_129 = popcount35_kfnc_core_126 | popcount35_kfnc_core_128;
  assign popcount35_kfnc_core_132 = ~input_a[17];
  assign popcount35_kfnc_core_133 = input_a[17] & input_a[28];
  assign popcount35_kfnc_core_135 = input_a[19] & input_a[18];
  assign popcount35_kfnc_core_138 = popcount35_kfnc_core_133 ^ popcount35_kfnc_core_135;
  assign popcount35_kfnc_core_139 = popcount35_kfnc_core_133 & popcount35_kfnc_core_135;
  assign popcount35_kfnc_core_143 = input_a[21] & input_a[22];
  assign popcount35_kfnc_core_144 = input_a[21] & input_a[22];
  assign popcount35_kfnc_core_145 = input_a[3] ^ input_a[13];
  assign popcount35_kfnc_core_146 = input_a[24] & input_a[21];
  assign popcount35_kfnc_core_147 = input_a[19] ^ popcount35_kfnc_core_145;
  assign popcount35_kfnc_core_149 = popcount35_kfnc_core_146 ^ input_a[12];
  assign popcount35_kfnc_core_150 = popcount35_kfnc_core_146 & input_a[12];
  assign popcount35_kfnc_core_151 = ~input_a[26];
  assign popcount35_kfnc_core_153 = input_a[13] ^ popcount35_kfnc_core_149;
  assign popcount35_kfnc_core_161 = input_a[16] & input_a[16];
  assign popcount35_kfnc_core_162_not = ~popcount35_kfnc_core_138;
  assign popcount35_kfnc_core_164 = popcount35_kfnc_core_162_not ^ popcount35_kfnc_core_161;
  assign popcount35_kfnc_core_165 = popcount35_kfnc_core_162_not & popcount35_kfnc_core_161;
  assign popcount35_kfnc_core_166 = popcount35_kfnc_core_138 | popcount35_kfnc_core_165;
  assign popcount35_kfnc_core_167 = popcount35_kfnc_core_139 ^ popcount35_kfnc_core_150;
  assign popcount35_kfnc_core_169 = popcount35_kfnc_core_167 ^ popcount35_kfnc_core_166;
  assign popcount35_kfnc_core_170 = popcount35_kfnc_core_167 & popcount35_kfnc_core_166;
  assign popcount35_kfnc_core_174 = input_a[26] ^ input_a[20];
  assign popcount35_kfnc_core_175 = input_a[25] & input_a[27];
  assign popcount35_kfnc_core_176 = ~input_a[28];
  assign popcount35_kfnc_core_177 = input_a[28] & input_a[20];
  assign popcount35_kfnc_core_178 = input_a[17] ^ popcount35_kfnc_core_176;
  assign popcount35_kfnc_core_179 = input_a[27] & popcount35_kfnc_core_176;
  assign popcount35_kfnc_core_180 = popcount35_kfnc_core_175 ^ popcount35_kfnc_core_177;
  assign popcount35_kfnc_core_181 = popcount35_kfnc_core_175 & input_a[15];
  assign popcount35_kfnc_core_182 = popcount35_kfnc_core_180 ^ input_a[9];
  assign popcount35_kfnc_core_183 = popcount35_kfnc_core_180 & input_a[15];
  assign popcount35_kfnc_core_184 = popcount35_kfnc_core_181 | popcount35_kfnc_core_183;
  assign popcount35_kfnc_core_185 = input_a[22] ^ input_a[31];
  assign popcount35_kfnc_core_187 = input_a[33] ^ input_a[34];
  assign popcount35_kfnc_core_188 = input_a[33] & input_a[34];
  assign popcount35_kfnc_core_189 = input_a[32] ^ input_a[0];
  assign popcount35_kfnc_core_190 = input_a[32] & popcount35_kfnc_core_187;
  assign popcount35_kfnc_core_191 = popcount35_kfnc_core_188 ^ popcount35_kfnc_core_190;
  assign popcount35_kfnc_core_192 = popcount35_kfnc_core_188 & popcount35_kfnc_core_190;
  assign popcount35_kfnc_core_193 = popcount35_kfnc_core_185 ^ popcount35_kfnc_core_189;
  assign popcount35_kfnc_core_194 = popcount35_kfnc_core_185 & popcount35_kfnc_core_189;
  assign popcount35_kfnc_core_197 = popcount35_kfnc_core_191 ^ popcount35_kfnc_core_194;
  assign popcount35_kfnc_core_198 = popcount35_kfnc_core_191 & popcount35_kfnc_core_194;
  assign popcount35_kfnc_core_200 = popcount35_kfnc_core_192 ^ popcount35_kfnc_core_198;
  assign popcount35_kfnc_core_201 = popcount35_kfnc_core_192 & input_a[11];
  assign popcount35_kfnc_core_202 = ~(popcount35_kfnc_core_178 & input_a[0]);
  assign popcount35_kfnc_core_203 = popcount35_kfnc_core_178 & popcount35_kfnc_core_193;
  assign popcount35_kfnc_core_204 = popcount35_kfnc_core_182 ^ popcount35_kfnc_core_197;
  assign popcount35_kfnc_core_205 = popcount35_kfnc_core_182 & popcount35_kfnc_core_197;
  assign popcount35_kfnc_core_206 = popcount35_kfnc_core_204 ^ popcount35_kfnc_core_203;
  assign popcount35_kfnc_core_207 = popcount35_kfnc_core_204 & popcount35_kfnc_core_203;
  assign popcount35_kfnc_core_208 = popcount35_kfnc_core_205 | popcount35_kfnc_core_207;
  assign popcount35_kfnc_core_209 = popcount35_kfnc_core_184 | popcount35_kfnc_core_200;
  assign popcount35_kfnc_core_210 = popcount35_kfnc_core_184 & popcount35_kfnc_core_200;
  assign popcount35_kfnc_core_211 = popcount35_kfnc_core_209 ^ popcount35_kfnc_core_208;
  assign popcount35_kfnc_core_212 = popcount35_kfnc_core_209 & popcount35_kfnc_core_208;
  assign popcount35_kfnc_core_213 = popcount35_kfnc_core_210 & input_a[3];
  assign popcount35_kfnc_core_214 = popcount35_kfnc_core_201 ^ popcount35_kfnc_core_213;
  assign popcount35_kfnc_core_215 = popcount35_kfnc_core_201 & input_a[8];
  assign popcount35_kfnc_core_216 = ~input_a[23];
  assign popcount35_kfnc_core_217 = input_a[0] & popcount35_kfnc_core_202;
  assign popcount35_kfnc_core_218 = popcount35_kfnc_core_164 ^ popcount35_kfnc_core_206;
  assign popcount35_kfnc_core_219 = popcount35_kfnc_core_164 & popcount35_kfnc_core_206;
  assign popcount35_kfnc_core_220 = popcount35_kfnc_core_218 ^ input_a[24];
  assign popcount35_kfnc_core_221 = popcount35_kfnc_core_218 & popcount35_kfnc_core_217;
  assign popcount35_kfnc_core_222 = popcount35_kfnc_core_219 | popcount35_kfnc_core_221;
  assign popcount35_kfnc_core_223 = popcount35_kfnc_core_169 ^ popcount35_kfnc_core_211;
  assign popcount35_kfnc_core_224 = popcount35_kfnc_core_169 & popcount35_kfnc_core_211;
  assign popcount35_kfnc_core_225 = popcount35_kfnc_core_223 ^ popcount35_kfnc_core_222;
  assign popcount35_kfnc_core_226 = popcount35_kfnc_core_223 & popcount35_kfnc_core_222;
  assign popcount35_kfnc_core_227 = popcount35_kfnc_core_224 | popcount35_kfnc_core_226;
  assign popcount35_kfnc_core_228 = popcount35_kfnc_core_170 ^ popcount35_kfnc_core_214;
  assign popcount35_kfnc_core_229 = input_a[2] & popcount35_kfnc_core_214;
  assign popcount35_kfnc_core_230 = popcount35_kfnc_core_228 ^ popcount35_kfnc_core_227;
  assign popcount35_kfnc_core_231 = popcount35_kfnc_core_228 & popcount35_kfnc_core_227;
  assign popcount35_kfnc_core_232 = popcount35_kfnc_core_229 | popcount35_kfnc_core_231;
  assign popcount35_kfnc_core_234 = input_a[16] & popcount35_kfnc_core_215;
  assign popcount35_kfnc_core_235 = popcount35_kfnc_core_215 ^ popcount35_kfnc_core_232;
  assign popcount35_kfnc_core_236 = popcount35_kfnc_core_215 & popcount35_kfnc_core_232;
  assign popcount35_kfnc_core_237 = popcount35_kfnc_core_234 | popcount35_kfnc_core_236;
  assign popcount35_kfnc_core_238 = ~(input_a[10] ^ input_a[30]);
  assign popcount35_kfnc_core_239 = input_a[10] & input_a[27];
  assign popcount35_kfnc_core_241 = popcount35_kfnc_core_117 & input_a[5];
  assign popcount35_kfnc_core_242 = input_a[7] ^ popcount35_kfnc_core_239;
  assign popcount35_kfnc_core_243 = input_a[7] & popcount35_kfnc_core_239;
  assign popcount35_kfnc_core_244 = popcount35_kfnc_core_241 | popcount35_kfnc_core_243;
  assign popcount35_kfnc_core_245 = popcount35_kfnc_core_122 ^ popcount35_kfnc_core_225;
  assign popcount35_kfnc_core_246 = popcount35_kfnc_core_122 & popcount35_kfnc_core_225;
  assign popcount35_kfnc_core_247 = popcount35_kfnc_core_245 ^ popcount35_kfnc_core_244;
  assign popcount35_kfnc_core_248 = popcount35_kfnc_core_245 & popcount35_kfnc_core_244;
  assign popcount35_kfnc_core_249 = popcount35_kfnc_core_246 | popcount35_kfnc_core_248;
  assign popcount35_kfnc_core_250 = popcount35_kfnc_core_127 ^ popcount35_kfnc_core_230;
  assign popcount35_kfnc_core_251 = popcount35_kfnc_core_127 & popcount35_kfnc_core_230;
  assign popcount35_kfnc_core_252 = popcount35_kfnc_core_250 ^ popcount35_kfnc_core_249;
  assign popcount35_kfnc_core_253 = popcount35_kfnc_core_250 & popcount35_kfnc_core_249;
  assign popcount35_kfnc_core_254 = popcount35_kfnc_core_251 | popcount35_kfnc_core_253;
  assign popcount35_kfnc_core_257 = popcount35_kfnc_core_235 ^ popcount35_kfnc_core_254;
  assign popcount35_kfnc_core_258 = popcount35_kfnc_core_235 & popcount35_kfnc_core_254;
  assign popcount35_kfnc_core_261_not = ~popcount35_kfnc_core_237;
  assign popcount35_kfnc_core_262 = popcount35_kfnc_core_237 | popcount35_kfnc_core_258;
  assign popcount35_kfnc_core_263 = popcount35_kfnc_core_237 & input_a[22];
  assign popcount35_kfnc_core_264 = input_a[10] | input_a[34];

  assign popcount35_kfnc_out[0] = popcount35_kfnc_core_170;
  assign popcount35_kfnc_out[1] = popcount35_kfnc_core_242;
  assign popcount35_kfnc_out[2] = popcount35_kfnc_core_247;
  assign popcount35_kfnc_out[3] = popcount35_kfnc_core_252;
  assign popcount35_kfnc_out[4] = popcount35_kfnc_core_257;
  assign popcount35_kfnc_out[5] = popcount35_kfnc_core_262;
endmodule