// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.12171
// WCE=30.0
// EP=0.972364%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_vmye(input [35:0] input_a, output [5:0] popcount36_vmye_out);
  wire popcount36_vmye_core_038;
  wire popcount36_vmye_core_039;
  wire popcount36_vmye_core_040;
  wire popcount36_vmye_core_041;
  wire popcount36_vmye_core_042;
  wire popcount36_vmye_core_043;
  wire popcount36_vmye_core_044;
  wire popcount36_vmye_core_045;
  wire popcount36_vmye_core_046;
  wire popcount36_vmye_core_047;
  wire popcount36_vmye_core_049;
  wire popcount36_vmye_core_050;
  wire popcount36_vmye_core_051;
  wire popcount36_vmye_core_052;
  wire popcount36_vmye_core_053;
  wire popcount36_vmye_core_054;
  wire popcount36_vmye_core_055;
  wire popcount36_vmye_core_056;
  wire popcount36_vmye_core_057;
  wire popcount36_vmye_core_061;
  wire popcount36_vmye_core_062;
  wire popcount36_vmye_core_065;
  wire popcount36_vmye_core_066;
  wire popcount36_vmye_core_067;
  wire popcount36_vmye_core_068;
  wire popcount36_vmye_core_070;
  wire popcount36_vmye_core_072;
  wire popcount36_vmye_core_073_not;
  wire popcount36_vmye_core_075;
  wire popcount36_vmye_core_077;
  wire popcount36_vmye_core_078;
  wire popcount36_vmye_core_080;
  wire popcount36_vmye_core_081;
  wire popcount36_vmye_core_083;
  wire popcount36_vmye_core_084;
  wire popcount36_vmye_core_086;
  wire popcount36_vmye_core_087;
  wire popcount36_vmye_core_088;
  wire popcount36_vmye_core_090;
  wire popcount36_vmye_core_091;
  wire popcount36_vmye_core_092;
  wire popcount36_vmye_core_093;
  wire popcount36_vmye_core_094;
  wire popcount36_vmye_core_095;
  wire popcount36_vmye_core_096;
  wire popcount36_vmye_core_099;
  wire popcount36_vmye_core_100;
  wire popcount36_vmye_core_103;
  wire popcount36_vmye_core_104;
  wire popcount36_vmye_core_107;
  wire popcount36_vmye_core_108;
  wire popcount36_vmye_core_109;
  wire popcount36_vmye_core_110;
  wire popcount36_vmye_core_111;
  wire popcount36_vmye_core_112;
  wire popcount36_vmye_core_114;
  wire popcount36_vmye_core_115;
  wire popcount36_vmye_core_116;
  wire popcount36_vmye_core_117;
  wire popcount36_vmye_core_118;
  wire popcount36_vmye_core_120;
  wire popcount36_vmye_core_123;
  wire popcount36_vmye_core_125;
  wire popcount36_vmye_core_128;
  wire popcount36_vmye_core_129;
  wire popcount36_vmye_core_130;
  wire popcount36_vmye_core_132;
  wire popcount36_vmye_core_133;
  wire popcount36_vmye_core_135;
  wire popcount36_vmye_core_139;
  wire popcount36_vmye_core_143;
  wire popcount36_vmye_core_144;
  wire popcount36_vmye_core_145;
  wire popcount36_vmye_core_147;
  wire popcount36_vmye_core_148;
  wire popcount36_vmye_core_149;
  wire popcount36_vmye_core_150;
  wire popcount36_vmye_core_151;
  wire popcount36_vmye_core_154;
  wire popcount36_vmye_core_157;
  wire popcount36_vmye_core_158;
  wire popcount36_vmye_core_160;
  wire popcount36_vmye_core_161;
  wire popcount36_vmye_core_162;
  wire popcount36_vmye_core_164;
  wire popcount36_vmye_core_166;
  wire popcount36_vmye_core_167_not;
  wire popcount36_vmye_core_168;
  wire popcount36_vmye_core_169;
  wire popcount36_vmye_core_171;
  wire popcount36_vmye_core_172;
  wire popcount36_vmye_core_173;
  wire popcount36_vmye_core_175;
  wire popcount36_vmye_core_176;
  wire popcount36_vmye_core_177;
  wire popcount36_vmye_core_178_not;
  wire popcount36_vmye_core_179;
  wire popcount36_vmye_core_180;
  wire popcount36_vmye_core_183;
  wire popcount36_vmye_core_186;
  wire popcount36_vmye_core_188;
  wire popcount36_vmye_core_190;
  wire popcount36_vmye_core_191;
  wire popcount36_vmye_core_192;
  wire popcount36_vmye_core_193;
  wire popcount36_vmye_core_194;
  wire popcount36_vmye_core_195;
  wire popcount36_vmye_core_196;
  wire popcount36_vmye_core_199;
  wire popcount36_vmye_core_202;
  wire popcount36_vmye_core_203;
  wire popcount36_vmye_core_207;
  wire popcount36_vmye_core_208;
  wire popcount36_vmye_core_211;
  wire popcount36_vmye_core_212;
  wire popcount36_vmye_core_214;
  wire popcount36_vmye_core_215;
  wire popcount36_vmye_core_216;
  wire popcount36_vmye_core_217;
  wire popcount36_vmye_core_218;
  wire popcount36_vmye_core_219;
  wire popcount36_vmye_core_222;
  wire popcount36_vmye_core_223;
  wire popcount36_vmye_core_224;
  wire popcount36_vmye_core_225;
  wire popcount36_vmye_core_226;
  wire popcount36_vmye_core_228;
  wire popcount36_vmye_core_229;
  wire popcount36_vmye_core_230;
  wire popcount36_vmye_core_231;
  wire popcount36_vmye_core_233;
  wire popcount36_vmye_core_235;
  wire popcount36_vmye_core_236;
  wire popcount36_vmye_core_237;
  wire popcount36_vmye_core_238;
  wire popcount36_vmye_core_241;
  wire popcount36_vmye_core_242;
  wire popcount36_vmye_core_244;
  wire popcount36_vmye_core_245;
  wire popcount36_vmye_core_246;
  wire popcount36_vmye_core_249;
  wire popcount36_vmye_core_251;
  wire popcount36_vmye_core_252;
  wire popcount36_vmye_core_253;
  wire popcount36_vmye_core_254_not;
  wire popcount36_vmye_core_255;
  wire popcount36_vmye_core_256;
  wire popcount36_vmye_core_257;
  wire popcount36_vmye_core_258;
  wire popcount36_vmye_core_260;
  wire popcount36_vmye_core_261;
  wire popcount36_vmye_core_262;
  wire popcount36_vmye_core_263;
  wire popcount36_vmye_core_265;
  wire popcount36_vmye_core_266;
  wire popcount36_vmye_core_267;
  wire popcount36_vmye_core_268;
  wire popcount36_vmye_core_270;
  wire popcount36_vmye_core_272;
  wire popcount36_vmye_core_274;
  wire popcount36_vmye_core_275;
  wire popcount36_vmye_core_276;

  assign popcount36_vmye_core_038 = input_a[5] & input_a[15];
  assign popcount36_vmye_core_039 = input_a[7] ^ input_a[0];
  assign popcount36_vmye_core_040 = ~(input_a[11] ^ input_a[20]);
  assign popcount36_vmye_core_041 = input_a[35] ^ input_a[15];
  assign popcount36_vmye_core_042 = ~(input_a[19] & input_a[9]);
  assign popcount36_vmye_core_043 = input_a[6] | input_a[5];
  assign popcount36_vmye_core_044 = ~(input_a[30] | input_a[2]);
  assign popcount36_vmye_core_045 = ~(input_a[1] ^ input_a[34]);
  assign popcount36_vmye_core_046 = ~(input_a[15] & input_a[4]);
  assign popcount36_vmye_core_047 = ~(input_a[15] ^ input_a[2]);
  assign popcount36_vmye_core_049 = input_a[3] ^ input_a[10];
  assign popcount36_vmye_core_050 = input_a[31] & input_a[9];
  assign popcount36_vmye_core_051 = ~(input_a[8] ^ input_a[26]);
  assign popcount36_vmye_core_052 = ~input_a[35];
  assign popcount36_vmye_core_053 = ~input_a[30];
  assign popcount36_vmye_core_054 = ~(input_a[6] & input_a[0]);
  assign popcount36_vmye_core_055 = ~(input_a[19] ^ input_a[35]);
  assign popcount36_vmye_core_056 = input_a[29] & input_a[35];
  assign popcount36_vmye_core_057 = input_a[12] | input_a[4];
  assign popcount36_vmye_core_061 = input_a[10] ^ input_a[17];
  assign popcount36_vmye_core_062 = ~(input_a[13] & input_a[29]);
  assign popcount36_vmye_core_065 = ~(input_a[26] & input_a[20]);
  assign popcount36_vmye_core_066 = input_a[17] & input_a[35];
  assign popcount36_vmye_core_067 = input_a[26] ^ input_a[22];
  assign popcount36_vmye_core_068 = input_a[2] | input_a[7];
  assign popcount36_vmye_core_070 = ~(input_a[14] ^ input_a[12]);
  assign popcount36_vmye_core_072 = ~input_a[23];
  assign popcount36_vmye_core_073_not = ~input_a[18];
  assign popcount36_vmye_core_075 = input_a[33] ^ input_a[9];
  assign popcount36_vmye_core_077 = input_a[24] ^ input_a[34];
  assign popcount36_vmye_core_078 = ~(input_a[24] ^ input_a[4]);
  assign popcount36_vmye_core_080 = ~input_a[16];
  assign popcount36_vmye_core_081 = input_a[24] ^ input_a[34];
  assign popcount36_vmye_core_083 = ~input_a[7];
  assign popcount36_vmye_core_084 = input_a[28] | input_a[1];
  assign popcount36_vmye_core_086 = ~(input_a[2] ^ input_a[32]);
  assign popcount36_vmye_core_087 = ~input_a[7];
  assign popcount36_vmye_core_088 = input_a[35] | input_a[14];
  assign popcount36_vmye_core_090 = ~(input_a[16] | input_a[15]);
  assign popcount36_vmye_core_091 = ~input_a[21];
  assign popcount36_vmye_core_092 = ~input_a[11];
  assign popcount36_vmye_core_093 = input_a[24] ^ input_a[14];
  assign popcount36_vmye_core_094 = ~(input_a[26] | input_a[19]);
  assign popcount36_vmye_core_095 = ~(input_a[21] & input_a[22]);
  assign popcount36_vmye_core_096 = ~(input_a[29] | input_a[31]);
  assign popcount36_vmye_core_099 = ~(input_a[28] | input_a[13]);
  assign popcount36_vmye_core_100 = ~(input_a[9] | input_a[17]);
  assign popcount36_vmye_core_103 = input_a[0] | input_a[2];
  assign popcount36_vmye_core_104 = input_a[21] & input_a[20];
  assign popcount36_vmye_core_107 = ~(input_a[13] | input_a[11]);
  assign popcount36_vmye_core_108 = input_a[24] ^ input_a[9];
  assign popcount36_vmye_core_109 = ~(input_a[20] | input_a[30]);
  assign popcount36_vmye_core_110 = input_a[24] ^ input_a[11];
  assign popcount36_vmye_core_111 = ~(input_a[14] | input_a[6]);
  assign popcount36_vmye_core_112 = ~(input_a[16] ^ input_a[8]);
  assign popcount36_vmye_core_114 = input_a[34] ^ input_a[5];
  assign popcount36_vmye_core_115 = input_a[14] ^ input_a[16];
  assign popcount36_vmye_core_116 = ~(input_a[33] & input_a[29]);
  assign popcount36_vmye_core_117 = ~(input_a[19] | input_a[26]);
  assign popcount36_vmye_core_118 = ~(input_a[35] & input_a[28]);
  assign popcount36_vmye_core_120 = input_a[11] ^ input_a[20];
  assign popcount36_vmye_core_123 = input_a[18] & input_a[9];
  assign popcount36_vmye_core_125 = ~(input_a[1] ^ input_a[17]);
  assign popcount36_vmye_core_128 = ~(input_a[13] ^ input_a[17]);
  assign popcount36_vmye_core_129 = input_a[24] ^ input_a[34];
  assign popcount36_vmye_core_130 = ~(input_a[17] | input_a[24]);
  assign popcount36_vmye_core_132 = input_a[25] | input_a[7];
  assign popcount36_vmye_core_133 = input_a[27] | input_a[33];
  assign popcount36_vmye_core_135 = ~(input_a[22] & input_a[11]);
  assign popcount36_vmye_core_139 = ~(input_a[3] ^ input_a[7]);
  assign popcount36_vmye_core_143 = input_a[9] ^ input_a[13];
  assign popcount36_vmye_core_144 = ~input_a[3];
  assign popcount36_vmye_core_145 = ~input_a[8];
  assign popcount36_vmye_core_147 = input_a[33] | input_a[1];
  assign popcount36_vmye_core_148 = input_a[11] & input_a[22];
  assign popcount36_vmye_core_149 = ~input_a[9];
  assign popcount36_vmye_core_150 = ~(input_a[23] & input_a[4]);
  assign popcount36_vmye_core_151 = ~(input_a[17] & input_a[26]);
  assign popcount36_vmye_core_154 = ~(input_a[35] | input_a[29]);
  assign popcount36_vmye_core_157 = input_a[10] | input_a[25];
  assign popcount36_vmye_core_158 = ~input_a[35];
  assign popcount36_vmye_core_160 = ~(input_a[19] & input_a[17]);
  assign popcount36_vmye_core_161 = input_a[27] & input_a[16];
  assign popcount36_vmye_core_162 = ~(input_a[17] | input_a[32]);
  assign popcount36_vmye_core_164 = ~(input_a[9] | input_a[27]);
  assign popcount36_vmye_core_166 = ~(input_a[14] & input_a[34]);
  assign popcount36_vmye_core_167_not = ~input_a[24];
  assign popcount36_vmye_core_168 = ~(input_a[19] | input_a[26]);
  assign popcount36_vmye_core_169 = ~(input_a[5] | input_a[32]);
  assign popcount36_vmye_core_171 = input_a[23] | input_a[13];
  assign popcount36_vmye_core_172 = input_a[3] ^ input_a[8];
  assign popcount36_vmye_core_173 = input_a[25] | input_a[19];
  assign popcount36_vmye_core_175 = ~(input_a[14] ^ input_a[29]);
  assign popcount36_vmye_core_176 = ~input_a[34];
  assign popcount36_vmye_core_177 = input_a[5] | input_a[26];
  assign popcount36_vmye_core_178_not = ~input_a[0];
  assign popcount36_vmye_core_179 = ~(input_a[17] ^ input_a[23]);
  assign popcount36_vmye_core_180 = ~(input_a[12] ^ input_a[17]);
  assign popcount36_vmye_core_183 = ~(input_a[5] | input_a[16]);
  assign popcount36_vmye_core_186 = ~input_a[0];
  assign popcount36_vmye_core_188 = ~input_a[6];
  assign popcount36_vmye_core_190 = ~(input_a[35] & input_a[3]);
  assign popcount36_vmye_core_191 = input_a[23] | input_a[29];
  assign popcount36_vmye_core_192 = ~(input_a[16] ^ input_a[32]);
  assign popcount36_vmye_core_193 = input_a[28] ^ input_a[8];
  assign popcount36_vmye_core_194 = ~(input_a[8] & input_a[21]);
  assign popcount36_vmye_core_195 = input_a[10] & input_a[34];
  assign popcount36_vmye_core_196 = ~(input_a[7] | input_a[12]);
  assign popcount36_vmye_core_199 = ~(input_a[32] & input_a[25]);
  assign popcount36_vmye_core_202 = ~(input_a[18] | input_a[27]);
  assign popcount36_vmye_core_203 = input_a[30] ^ input_a[24];
  assign popcount36_vmye_core_207 = ~(input_a[22] & input_a[12]);
  assign popcount36_vmye_core_208 = ~(input_a[12] | input_a[9]);
  assign popcount36_vmye_core_211 = ~(input_a[12] | input_a[8]);
  assign popcount36_vmye_core_212 = ~input_a[20];
  assign popcount36_vmye_core_214 = input_a[14] | input_a[6];
  assign popcount36_vmye_core_215 = input_a[22] & input_a[14];
  assign popcount36_vmye_core_216 = input_a[17] & input_a[6];
  assign popcount36_vmye_core_217 = ~(input_a[10] ^ input_a[2]);
  assign popcount36_vmye_core_218 = input_a[15] ^ input_a[1];
  assign popcount36_vmye_core_219 = input_a[26] ^ input_a[19];
  assign popcount36_vmye_core_222 = input_a[33] | input_a[17];
  assign popcount36_vmye_core_223 = input_a[4] | input_a[30];
  assign popcount36_vmye_core_224 = input_a[31] | input_a[6];
  assign popcount36_vmye_core_225 = ~(input_a[28] & input_a[14]);
  assign popcount36_vmye_core_226 = ~input_a[13];
  assign popcount36_vmye_core_228 = ~(input_a[29] ^ input_a[21]);
  assign popcount36_vmye_core_229 = ~(input_a[14] ^ input_a[10]);
  assign popcount36_vmye_core_230 = input_a[33] | input_a[10];
  assign popcount36_vmye_core_231 = ~(input_a[23] & input_a[16]);
  assign popcount36_vmye_core_233 = ~(input_a[26] | input_a[31]);
  assign popcount36_vmye_core_235 = ~(input_a[4] | input_a[2]);
  assign popcount36_vmye_core_236 = input_a[20] ^ input_a[19];
  assign popcount36_vmye_core_237 = ~(input_a[32] & input_a[11]);
  assign popcount36_vmye_core_238 = ~(input_a[15] & input_a[11]);
  assign popcount36_vmye_core_241 = ~(input_a[1] ^ input_a[25]);
  assign popcount36_vmye_core_242 = input_a[4] & input_a[11];
  assign popcount36_vmye_core_244 = input_a[17] & input_a[30];
  assign popcount36_vmye_core_245 = ~(input_a[21] & input_a[1]);
  assign popcount36_vmye_core_246 = ~input_a[7];
  assign popcount36_vmye_core_249 = ~(input_a[5] | input_a[0]);
  assign popcount36_vmye_core_251 = ~(input_a[25] ^ input_a[25]);
  assign popcount36_vmye_core_252 = input_a[14] ^ input_a[30];
  assign popcount36_vmye_core_253 = ~(input_a[3] | input_a[28]);
  assign popcount36_vmye_core_254_not = ~input_a[2];
  assign popcount36_vmye_core_255 = ~(input_a[17] ^ input_a[0]);
  assign popcount36_vmye_core_256 = ~(input_a[27] ^ input_a[35]);
  assign popcount36_vmye_core_257 = input_a[34] ^ input_a[23];
  assign popcount36_vmye_core_258 = ~(input_a[9] ^ input_a[20]);
  assign popcount36_vmye_core_260 = input_a[0] | input_a[29];
  assign popcount36_vmye_core_261 = ~(input_a[5] ^ input_a[23]);
  assign popcount36_vmye_core_262 = input_a[32] & input_a[11];
  assign popcount36_vmye_core_263 = input_a[2] & input_a[31];
  assign popcount36_vmye_core_265 = ~(input_a[15] ^ input_a[12]);
  assign popcount36_vmye_core_266 = ~input_a[22];
  assign popcount36_vmye_core_267 = ~(input_a[11] & input_a[0]);
  assign popcount36_vmye_core_268 = ~(input_a[20] | input_a[32]);
  assign popcount36_vmye_core_270 = input_a[14] ^ input_a[28];
  assign popcount36_vmye_core_272 = input_a[22] | input_a[17];
  assign popcount36_vmye_core_274 = ~(input_a[20] | input_a[8]);
  assign popcount36_vmye_core_275 = ~(input_a[22] & input_a[17]);
  assign popcount36_vmye_core_276 = ~input_a[11];

  assign popcount36_vmye_out[0] = 1'b1;
  assign popcount36_vmye_out[1] = input_a[25];
  assign popcount36_vmye_out[2] = 1'b1;
  assign popcount36_vmye_out[3] = 1'b1;
  assign popcount36_vmye_out[4] = 1'b1;
  assign popcount36_vmye_out[5] = 1'b0;
endmodule