// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.55489
// WCE=22.0
// EP=0.977469%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_h8wc(input [33:0] input_a, output [5:0] popcount34_h8wc_out);
  wire popcount34_h8wc_core_036;
  wire popcount34_h8wc_core_040;
  wire popcount34_h8wc_core_041;
  wire popcount34_h8wc_core_043;
  wire popcount34_h8wc_core_045;
  wire popcount34_h8wc_core_046;
  wire popcount34_h8wc_core_048;
  wire popcount34_h8wc_core_049;
  wire popcount34_h8wc_core_052;
  wire popcount34_h8wc_core_053;
  wire popcount34_h8wc_core_054;
  wire popcount34_h8wc_core_055;
  wire popcount34_h8wc_core_056;
  wire popcount34_h8wc_core_057;
  wire popcount34_h8wc_core_058;
  wire popcount34_h8wc_core_059;
  wire popcount34_h8wc_core_061;
  wire popcount34_h8wc_core_062;
  wire popcount34_h8wc_core_063;
  wire popcount34_h8wc_core_064;
  wire popcount34_h8wc_core_066;
  wire popcount34_h8wc_core_068;
  wire popcount34_h8wc_core_069;
  wire popcount34_h8wc_core_070;
  wire popcount34_h8wc_core_071;
  wire popcount34_h8wc_core_072;
  wire popcount34_h8wc_core_073;
  wire popcount34_h8wc_core_074;
  wire popcount34_h8wc_core_077;
  wire popcount34_h8wc_core_079;
  wire popcount34_h8wc_core_080;
  wire popcount34_h8wc_core_081;
  wire popcount34_h8wc_core_082;
  wire popcount34_h8wc_core_084;
  wire popcount34_h8wc_core_085;
  wire popcount34_h8wc_core_086;
  wire popcount34_h8wc_core_087;
  wire popcount34_h8wc_core_088;
  wire popcount34_h8wc_core_089;
  wire popcount34_h8wc_core_090;
  wire popcount34_h8wc_core_092;
  wire popcount34_h8wc_core_094;
  wire popcount34_h8wc_core_095;
  wire popcount34_h8wc_core_096;
  wire popcount34_h8wc_core_099;
  wire popcount34_h8wc_core_101;
  wire popcount34_h8wc_core_103;
  wire popcount34_h8wc_core_104;
  wire popcount34_h8wc_core_105;
  wire popcount34_h8wc_core_107;
  wire popcount34_h8wc_core_109;
  wire popcount34_h8wc_core_110;
  wire popcount34_h8wc_core_111;
  wire popcount34_h8wc_core_112;
  wire popcount34_h8wc_core_117;
  wire popcount34_h8wc_core_118;
  wire popcount34_h8wc_core_120;
  wire popcount34_h8wc_core_121;
  wire popcount34_h8wc_core_122;
  wire popcount34_h8wc_core_124;
  wire popcount34_h8wc_core_125;
  wire popcount34_h8wc_core_126;
  wire popcount34_h8wc_core_127;
  wire popcount34_h8wc_core_128;
  wire popcount34_h8wc_core_130;
  wire popcount34_h8wc_core_132;
  wire popcount34_h8wc_core_135;
  wire popcount34_h8wc_core_136;
  wire popcount34_h8wc_core_139;
  wire popcount34_h8wc_core_140;
  wire popcount34_h8wc_core_142;
  wire popcount34_h8wc_core_144;
  wire popcount34_h8wc_core_146;
  wire popcount34_h8wc_core_150;
  wire popcount34_h8wc_core_154;
  wire popcount34_h8wc_core_155;
  wire popcount34_h8wc_core_156;
  wire popcount34_h8wc_core_157;
  wire popcount34_h8wc_core_158;
  wire popcount34_h8wc_core_159_not;
  wire popcount34_h8wc_core_162;
  wire popcount34_h8wc_core_164;
  wire popcount34_h8wc_core_165;
  wire popcount34_h8wc_core_166;
  wire popcount34_h8wc_core_168;
  wire popcount34_h8wc_core_169;
  wire popcount34_h8wc_core_171;
  wire popcount34_h8wc_core_173;
  wire popcount34_h8wc_core_175;
  wire popcount34_h8wc_core_176;
  wire popcount34_h8wc_core_178;
  wire popcount34_h8wc_core_179;
  wire popcount34_h8wc_core_180;
  wire popcount34_h8wc_core_181;
  wire popcount34_h8wc_core_183_not;
  wire popcount34_h8wc_core_185;
  wire popcount34_h8wc_core_186;
  wire popcount34_h8wc_core_189;
  wire popcount34_h8wc_core_190;
  wire popcount34_h8wc_core_191;
  wire popcount34_h8wc_core_194;
  wire popcount34_h8wc_core_196;
  wire popcount34_h8wc_core_197;
  wire popcount34_h8wc_core_198;
  wire popcount34_h8wc_core_202;
  wire popcount34_h8wc_core_203;
  wire popcount34_h8wc_core_204;
  wire popcount34_h8wc_core_205;
  wire popcount34_h8wc_core_207;
  wire popcount34_h8wc_core_208;
  wire popcount34_h8wc_core_210;
  wire popcount34_h8wc_core_213;
  wire popcount34_h8wc_core_217;
  wire popcount34_h8wc_core_218;
  wire popcount34_h8wc_core_220;
  wire popcount34_h8wc_core_221;
  wire popcount34_h8wc_core_222;
  wire popcount34_h8wc_core_223;
  wire popcount34_h8wc_core_224;
  wire popcount34_h8wc_core_225;
  wire popcount34_h8wc_core_226;
  wire popcount34_h8wc_core_230;
  wire popcount34_h8wc_core_231;
  wire popcount34_h8wc_core_232;
  wire popcount34_h8wc_core_233;
  wire popcount34_h8wc_core_237;
  wire popcount34_h8wc_core_238;
  wire popcount34_h8wc_core_240;
  wire popcount34_h8wc_core_242;
  wire popcount34_h8wc_core_243;
  wire popcount34_h8wc_core_250;
  wire popcount34_h8wc_core_251;
  wire popcount34_h8wc_core_252;

  assign popcount34_h8wc_core_036 = input_a[9] | input_a[8];
  assign popcount34_h8wc_core_040 = ~input_a[12];
  assign popcount34_h8wc_core_041 = input_a[5] & input_a[32];
  assign popcount34_h8wc_core_043 = input_a[21] | input_a[3];
  assign popcount34_h8wc_core_045 = input_a[26] ^ input_a[5];
  assign popcount34_h8wc_core_046 = input_a[24] | input_a[1];
  assign popcount34_h8wc_core_048 = input_a[29] & input_a[28];
  assign popcount34_h8wc_core_049 = ~(input_a[1] | input_a[19]);
  assign popcount34_h8wc_core_052 = ~(input_a[21] & input_a[26]);
  assign popcount34_h8wc_core_053 = ~(input_a[4] & input_a[7]);
  assign popcount34_h8wc_core_054 = input_a[23] | input_a[8];
  assign popcount34_h8wc_core_055 = ~input_a[32];
  assign popcount34_h8wc_core_056 = ~(input_a[8] ^ input_a[0]);
  assign popcount34_h8wc_core_057 = ~(input_a[25] ^ input_a[17]);
  assign popcount34_h8wc_core_058 = input_a[14] & input_a[21];
  assign popcount34_h8wc_core_059 = input_a[1] | input_a[10];
  assign popcount34_h8wc_core_061 = ~(input_a[16] | input_a[12]);
  assign popcount34_h8wc_core_062 = ~(input_a[21] | input_a[27]);
  assign popcount34_h8wc_core_063 = input_a[3] & input_a[16];
  assign popcount34_h8wc_core_064 = ~(input_a[3] ^ input_a[26]);
  assign popcount34_h8wc_core_066 = ~(input_a[21] | input_a[20]);
  assign popcount34_h8wc_core_068 = ~(input_a[5] ^ input_a[25]);
  assign popcount34_h8wc_core_069 = input_a[6] & input_a[2];
  assign popcount34_h8wc_core_070 = ~(input_a[15] & input_a[24]);
  assign popcount34_h8wc_core_071 = input_a[9] | input_a[31];
  assign popcount34_h8wc_core_072 = ~(input_a[10] ^ input_a[26]);
  assign popcount34_h8wc_core_073 = ~(input_a[24] ^ input_a[24]);
  assign popcount34_h8wc_core_074 = input_a[5] & input_a[0];
  assign popcount34_h8wc_core_077 = ~(input_a[27] | input_a[20]);
  assign popcount34_h8wc_core_079 = input_a[8] | input_a[13];
  assign popcount34_h8wc_core_080 = ~(input_a[16] ^ input_a[18]);
  assign popcount34_h8wc_core_081 = ~input_a[13];
  assign popcount34_h8wc_core_082 = ~(input_a[5] & input_a[23]);
  assign popcount34_h8wc_core_084 = ~input_a[19];
  assign popcount34_h8wc_core_085 = input_a[33] & input_a[18];
  assign popcount34_h8wc_core_086 = ~input_a[18];
  assign popcount34_h8wc_core_087 = ~(input_a[27] & input_a[17]);
  assign popcount34_h8wc_core_088 = ~input_a[12];
  assign popcount34_h8wc_core_089 = ~input_a[17];
  assign popcount34_h8wc_core_090 = ~(input_a[18] ^ input_a[33]);
  assign popcount34_h8wc_core_092 = input_a[13] & input_a[10];
  assign popcount34_h8wc_core_094 = ~(input_a[26] ^ input_a[16]);
  assign popcount34_h8wc_core_095 = input_a[8] & input_a[12];
  assign popcount34_h8wc_core_096 = input_a[13] & input_a[18];
  assign popcount34_h8wc_core_099 = input_a[26] & input_a[6];
  assign popcount34_h8wc_core_101 = ~(input_a[19] | input_a[12]);
  assign popcount34_h8wc_core_103 = ~(input_a[0] & input_a[11]);
  assign popcount34_h8wc_core_104 = ~(input_a[5] & input_a[20]);
  assign popcount34_h8wc_core_105 = ~(input_a[17] | input_a[15]);
  assign popcount34_h8wc_core_107 = input_a[0] | input_a[29];
  assign popcount34_h8wc_core_109 = ~(input_a[15] & input_a[4]);
  assign popcount34_h8wc_core_110 = ~input_a[12];
  assign popcount34_h8wc_core_111 = ~(input_a[28] & input_a[19]);
  assign popcount34_h8wc_core_112 = ~(input_a[8] | input_a[10]);
  assign popcount34_h8wc_core_117 = input_a[26] ^ input_a[29];
  assign popcount34_h8wc_core_118 = ~input_a[23];
  assign popcount34_h8wc_core_120 = ~(input_a[25] ^ input_a[25]);
  assign popcount34_h8wc_core_121 = input_a[31] ^ input_a[28];
  assign popcount34_h8wc_core_122 = input_a[8] ^ input_a[16];
  assign popcount34_h8wc_core_124 = input_a[31] & input_a[10];
  assign popcount34_h8wc_core_125 = ~(input_a[1] ^ input_a[16]);
  assign popcount34_h8wc_core_126 = ~(input_a[18] ^ input_a[13]);
  assign popcount34_h8wc_core_127 = input_a[4] & input_a[26];
  assign popcount34_h8wc_core_128 = input_a[23] | input_a[32];
  assign popcount34_h8wc_core_130 = ~(input_a[15] & input_a[0]);
  assign popcount34_h8wc_core_132 = ~(input_a[0] ^ input_a[23]);
  assign popcount34_h8wc_core_135 = input_a[20] ^ input_a[5];
  assign popcount34_h8wc_core_136 = input_a[26] | input_a[11];
  assign popcount34_h8wc_core_139 = input_a[4] | input_a[8];
  assign popcount34_h8wc_core_140 = input_a[30] & input_a[8];
  assign popcount34_h8wc_core_142 = ~(input_a[3] & input_a[18]);
  assign popcount34_h8wc_core_144 = ~(input_a[27] & input_a[29]);
  assign popcount34_h8wc_core_146 = ~input_a[14];
  assign popcount34_h8wc_core_150 = input_a[27] ^ input_a[1];
  assign popcount34_h8wc_core_154 = ~(input_a[12] | input_a[13]);
  assign popcount34_h8wc_core_155 = ~(input_a[3] | input_a[17]);
  assign popcount34_h8wc_core_156 = input_a[0] | input_a[25];
  assign popcount34_h8wc_core_157 = ~(input_a[18] & input_a[27]);
  assign popcount34_h8wc_core_158 = ~(input_a[22] ^ input_a[21]);
  assign popcount34_h8wc_core_159_not = ~input_a[28];
  assign popcount34_h8wc_core_162 = ~(input_a[2] | input_a[25]);
  assign popcount34_h8wc_core_164 = input_a[31] ^ input_a[22];
  assign popcount34_h8wc_core_165 = ~(input_a[27] | input_a[21]);
  assign popcount34_h8wc_core_166 = ~(input_a[1] & input_a[1]);
  assign popcount34_h8wc_core_168 = input_a[0] | input_a[12];
  assign popcount34_h8wc_core_169 = input_a[24] & input_a[17];
  assign popcount34_h8wc_core_171 = input_a[10] & input_a[15];
  assign popcount34_h8wc_core_173 = input_a[29] | input_a[3];
  assign popcount34_h8wc_core_175 = input_a[1] & input_a[3];
  assign popcount34_h8wc_core_176 = ~(input_a[28] & input_a[20]);
  assign popcount34_h8wc_core_178 = ~(input_a[20] | input_a[14]);
  assign popcount34_h8wc_core_179 = ~(input_a[27] & input_a[17]);
  assign popcount34_h8wc_core_180 = ~(input_a[27] | input_a[7]);
  assign popcount34_h8wc_core_181 = ~input_a[1];
  assign popcount34_h8wc_core_183_not = ~input_a[9];
  assign popcount34_h8wc_core_185 = input_a[2] ^ input_a[21];
  assign popcount34_h8wc_core_186 = input_a[14] & input_a[3];
  assign popcount34_h8wc_core_189 = ~input_a[6];
  assign popcount34_h8wc_core_190 = input_a[9] | input_a[16];
  assign popcount34_h8wc_core_191 = ~(input_a[25] | input_a[15]);
  assign popcount34_h8wc_core_194 = ~(input_a[15] & input_a[33]);
  assign popcount34_h8wc_core_196 = input_a[24] | input_a[9];
  assign popcount34_h8wc_core_197 = ~input_a[3];
  assign popcount34_h8wc_core_198 = ~input_a[1];
  assign popcount34_h8wc_core_202 = ~input_a[26];
  assign popcount34_h8wc_core_203 = ~(input_a[27] | input_a[17]);
  assign popcount34_h8wc_core_204 = input_a[23] | input_a[3];
  assign popcount34_h8wc_core_205 = input_a[20] & input_a[10];
  assign popcount34_h8wc_core_207 = ~(input_a[13] | input_a[0]);
  assign popcount34_h8wc_core_208 = input_a[31] & input_a[8];
  assign popcount34_h8wc_core_210 = input_a[16] & input_a[25];
  assign popcount34_h8wc_core_213 = ~(input_a[26] | input_a[23]);
  assign popcount34_h8wc_core_217 = input_a[13] | input_a[25];
  assign popcount34_h8wc_core_218 = ~input_a[19];
  assign popcount34_h8wc_core_220 = input_a[26] | input_a[14];
  assign popcount34_h8wc_core_221 = ~(input_a[25] ^ input_a[21]);
  assign popcount34_h8wc_core_222 = input_a[8] & input_a[32];
  assign popcount34_h8wc_core_223 = ~(input_a[33] ^ input_a[16]);
  assign popcount34_h8wc_core_224 = ~(input_a[22] & input_a[7]);
  assign popcount34_h8wc_core_225 = input_a[14] | input_a[17];
  assign popcount34_h8wc_core_226 = input_a[20] ^ input_a[1];
  assign popcount34_h8wc_core_230 = input_a[9] | input_a[25];
  assign popcount34_h8wc_core_231 = input_a[26] | input_a[29];
  assign popcount34_h8wc_core_232 = ~(input_a[22] | input_a[2]);
  assign popcount34_h8wc_core_233 = ~input_a[18];
  assign popcount34_h8wc_core_237 = ~(input_a[3] & input_a[31]);
  assign popcount34_h8wc_core_238 = input_a[19] ^ input_a[3];
  assign popcount34_h8wc_core_240 = input_a[8] ^ input_a[29];
  assign popcount34_h8wc_core_242 = ~(input_a[31] & input_a[29]);
  assign popcount34_h8wc_core_243 = ~input_a[21];
  assign popcount34_h8wc_core_250 = ~(input_a[26] & input_a[1]);
  assign popcount34_h8wc_core_251 = ~input_a[33];
  assign popcount34_h8wc_core_252 = input_a[5] | input_a[24];

  assign popcount34_h8wc_out[0] = input_a[17];
  assign popcount34_h8wc_out[1] = 1'b1;
  assign popcount34_h8wc_out[2] = 1'b1;
  assign popcount34_h8wc_out[3] = 1'b0;
  assign popcount34_h8wc_out[4] = 1'b1;
  assign popcount34_h8wc_out[5] = 1'b0;
endmodule