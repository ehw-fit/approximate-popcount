// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.59654
// WCE=11.0
// EP=0.805715%
// Printed PDK parameters:
//  Area=32714223.0
//  Delay=61172684.0
//  Power=1906800.0

module popcount32_lqzk(input [31:0] input_a, output [5:0] popcount32_lqzk_out);
  wire popcount32_lqzk_core_034;
  wire popcount32_lqzk_core_035;
  wire popcount32_lqzk_core_037;
  wire popcount32_lqzk_core_038;
  wire popcount32_lqzk_core_039;
  wire popcount32_lqzk_core_040;
  wire popcount32_lqzk_core_042;
  wire popcount32_lqzk_core_043;
  wire popcount32_lqzk_core_044;
  wire popcount32_lqzk_core_045;
  wire popcount32_lqzk_core_047;
  wire popcount32_lqzk_core_048;
  wire popcount32_lqzk_core_051;
  wire popcount32_lqzk_core_053;
  wire popcount32_lqzk_core_054;
  wire popcount32_lqzk_core_055;
  wire popcount32_lqzk_core_056;
  wire popcount32_lqzk_core_057;
  wire popcount32_lqzk_core_058;
  wire popcount32_lqzk_core_061;
  wire popcount32_lqzk_core_064;
  wire popcount32_lqzk_core_066;
  wire popcount32_lqzk_core_068;
  wire popcount32_lqzk_core_071;
  wire popcount32_lqzk_core_072;
  wire popcount32_lqzk_core_073;
  wire popcount32_lqzk_core_074;
  wire popcount32_lqzk_core_075;
  wire popcount32_lqzk_core_076;
  wire popcount32_lqzk_core_078;
  wire popcount32_lqzk_core_082;
  wire popcount32_lqzk_core_083;
  wire popcount32_lqzk_core_084;
  wire popcount32_lqzk_core_085;
  wire popcount32_lqzk_core_087;
  wire popcount32_lqzk_core_088;
  wire popcount32_lqzk_core_089_not;
  wire popcount32_lqzk_core_090;
  wire popcount32_lqzk_core_092;
  wire popcount32_lqzk_core_093;
  wire popcount32_lqzk_core_095;
  wire popcount32_lqzk_core_098;
  wire popcount32_lqzk_core_100;
  wire popcount32_lqzk_core_101;
  wire popcount32_lqzk_core_102;
  wire popcount32_lqzk_core_104;
  wire popcount32_lqzk_core_106;
  wire popcount32_lqzk_core_108;
  wire popcount32_lqzk_core_109;
  wire popcount32_lqzk_core_111;
  wire popcount32_lqzk_core_113;
  wire popcount32_lqzk_core_117_not;
  wire popcount32_lqzk_core_118;
  wire popcount32_lqzk_core_121;
  wire popcount32_lqzk_core_122;
  wire popcount32_lqzk_core_125;
  wire popcount32_lqzk_core_126;
  wire popcount32_lqzk_core_128;
  wire popcount32_lqzk_core_130;
  wire popcount32_lqzk_core_131;
  wire popcount32_lqzk_core_132;
  wire popcount32_lqzk_core_133;
  wire popcount32_lqzk_core_135;
  wire popcount32_lqzk_core_136;
  wire popcount32_lqzk_core_138;
  wire popcount32_lqzk_core_139;
  wire popcount32_lqzk_core_142;
  wire popcount32_lqzk_core_143;
  wire popcount32_lqzk_core_144;
  wire popcount32_lqzk_core_145;
  wire popcount32_lqzk_core_146;
  wire popcount32_lqzk_core_147;
  wire popcount32_lqzk_core_149;
  wire popcount32_lqzk_core_150;
  wire popcount32_lqzk_core_151;
  wire popcount32_lqzk_core_153;
  wire popcount32_lqzk_core_154;
  wire popcount32_lqzk_core_155;
  wire popcount32_lqzk_core_156;
  wire popcount32_lqzk_core_157_not;
  wire popcount32_lqzk_core_158;
  wire popcount32_lqzk_core_159;
  wire popcount32_lqzk_core_161;
  wire popcount32_lqzk_core_162;
  wire popcount32_lqzk_core_164;
  wire popcount32_lqzk_core_165;
  wire popcount32_lqzk_core_167;
  wire popcount32_lqzk_core_169;
  wire popcount32_lqzk_core_171;
  wire popcount32_lqzk_core_172;
  wire popcount32_lqzk_core_173;
  wire popcount32_lqzk_core_176;
  wire popcount32_lqzk_core_177;
  wire popcount32_lqzk_core_178;
  wire popcount32_lqzk_core_180;
  wire popcount32_lqzk_core_183;
  wire popcount32_lqzk_core_185_not;
  wire popcount32_lqzk_core_186;
  wire popcount32_lqzk_core_188;
  wire popcount32_lqzk_core_189;
  wire popcount32_lqzk_core_190;
  wire popcount32_lqzk_core_191;
  wire popcount32_lqzk_core_192;
  wire popcount32_lqzk_core_193;
  wire popcount32_lqzk_core_194;
  wire popcount32_lqzk_core_195;
  wire popcount32_lqzk_core_196;
  wire popcount32_lqzk_core_197;
  wire popcount32_lqzk_core_198;
  wire popcount32_lqzk_core_200;
  wire popcount32_lqzk_core_202;
  wire popcount32_lqzk_core_203;
  wire popcount32_lqzk_core_204;
  wire popcount32_lqzk_core_205;
  wire popcount32_lqzk_core_206;
  wire popcount32_lqzk_core_207;
  wire popcount32_lqzk_core_208;
  wire popcount32_lqzk_core_209;
  wire popcount32_lqzk_core_210;
  wire popcount32_lqzk_core_211;
  wire popcount32_lqzk_core_212;
  wire popcount32_lqzk_core_213;
  wire popcount32_lqzk_core_214;
  wire popcount32_lqzk_core_215;
  wire popcount32_lqzk_core_216;
  wire popcount32_lqzk_core_217;
  wire popcount32_lqzk_core_218;
  wire popcount32_lqzk_core_219;
  wire popcount32_lqzk_core_220;
  wire popcount32_lqzk_core_221;
  wire popcount32_lqzk_core_223;
  wire popcount32_lqzk_core_225;

  assign popcount32_lqzk_core_034 = ~(input_a[7] | input_a[14]);
  assign popcount32_lqzk_core_035 = input_a[25] & input_a[1];
  assign popcount32_lqzk_core_037 = input_a[27] & input_a[21];
  assign popcount32_lqzk_core_038 = input_a[13] & input_a[4];
  assign popcount32_lqzk_core_039 = input_a[11] & input_a[20];
  assign popcount32_lqzk_core_040 = popcount32_lqzk_core_035 | popcount32_lqzk_core_037;
  assign popcount32_lqzk_core_042 = popcount32_lqzk_core_040 | popcount32_lqzk_core_039;
  assign popcount32_lqzk_core_043 = ~input_a[19];
  assign popcount32_lqzk_core_044 = ~input_a[26];
  assign popcount32_lqzk_core_045 = input_a[30] ^ input_a[21];
  assign popcount32_lqzk_core_047 = input_a[3] ^ input_a[24];
  assign popcount32_lqzk_core_048 = ~(input_a[11] | input_a[28]);
  assign popcount32_lqzk_core_051 = ~(input_a[15] & input_a[29]);
  assign popcount32_lqzk_core_053 = input_a[28] & input_a[16];
  assign popcount32_lqzk_core_054 = ~input_a[20];
  assign popcount32_lqzk_core_055 = ~input_a[19];
  assign popcount32_lqzk_core_056 = ~(input_a[18] & input_a[18]);
  assign popcount32_lqzk_core_057 = input_a[26] ^ input_a[7];
  assign popcount32_lqzk_core_058 = ~popcount32_lqzk_core_042;
  assign popcount32_lqzk_core_061 = input_a[14] & input_a[5];
  assign popcount32_lqzk_core_064 = input_a[16] | input_a[11];
  assign popcount32_lqzk_core_066 = ~(input_a[4] & input_a[22]);
  assign popcount32_lqzk_core_068 = ~(input_a[1] | input_a[30]);
  assign popcount32_lqzk_core_071 = input_a[26] & input_a[8];
  assign popcount32_lqzk_core_072 = input_a[23] ^ input_a[21];
  assign popcount32_lqzk_core_073 = input_a[23] ^ input_a[7];
  assign popcount32_lqzk_core_074 = input_a[23] | popcount32_lqzk_core_071;
  assign popcount32_lqzk_core_075 = input_a[21] & input_a[19];
  assign popcount32_lqzk_core_076 = popcount32_lqzk_core_074 | input_a[15];
  assign popcount32_lqzk_core_078 = input_a[26] ^ input_a[23];
  assign popcount32_lqzk_core_082 = ~(input_a[6] & input_a[24]);
  assign popcount32_lqzk_core_083 = ~input_a[8];
  assign popcount32_lqzk_core_084 = input_a[21] | input_a[8];
  assign popcount32_lqzk_core_085 = input_a[5] ^ input_a[27];
  assign popcount32_lqzk_core_087 = input_a[13] | input_a[30];
  assign popcount32_lqzk_core_088 = input_a[30] & input_a[9];
  assign popcount32_lqzk_core_089_not = ~input_a[22];
  assign popcount32_lqzk_core_090 = ~(input_a[11] | input_a[2]);
  assign popcount32_lqzk_core_092 = ~(popcount32_lqzk_core_076 & popcount32_lqzk_core_087);
  assign popcount32_lqzk_core_093 = popcount32_lqzk_core_076 & popcount32_lqzk_core_087;
  assign popcount32_lqzk_core_095 = input_a[23] ^ input_a[31];
  assign popcount32_lqzk_core_098 = input_a[18] ^ input_a[3];
  assign popcount32_lqzk_core_100 = ~(input_a[19] ^ input_a[11]);
  assign popcount32_lqzk_core_101 = ~(input_a[26] & input_a[5]);
  assign popcount32_lqzk_core_102 = input_a[9] ^ input_a[11];
  assign popcount32_lqzk_core_104 = popcount32_lqzk_core_058 ^ popcount32_lqzk_core_092;
  assign popcount32_lqzk_core_106 = ~popcount32_lqzk_core_104;
  assign popcount32_lqzk_core_108 = popcount32_lqzk_core_058 | popcount32_lqzk_core_104;
  assign popcount32_lqzk_core_109 = popcount32_lqzk_core_042 ^ popcount32_lqzk_core_093;
  assign popcount32_lqzk_core_111 = popcount32_lqzk_core_109 ^ popcount32_lqzk_core_108;
  assign popcount32_lqzk_core_113 = popcount32_lqzk_core_042 | popcount32_lqzk_core_109;
  assign popcount32_lqzk_core_117_not = ~input_a[23];
  assign popcount32_lqzk_core_118 = input_a[15] & input_a[9];
  assign popcount32_lqzk_core_121 = input_a[30] & input_a[4];
  assign popcount32_lqzk_core_122 = input_a[22] & input_a[18];
  assign popcount32_lqzk_core_125 = input_a[19] ^ popcount32_lqzk_core_122;
  assign popcount32_lqzk_core_126 = input_a[20] ^ input_a[17];
  assign popcount32_lqzk_core_128 = input_a[28] & input_a[2];
  assign popcount32_lqzk_core_130 = ~(input_a[20] ^ input_a[20]);
  assign popcount32_lqzk_core_131 = input_a[16] & input_a[31];
  assign popcount32_lqzk_core_132 = input_a[18] | input_a[25];
  assign popcount32_lqzk_core_133 = input_a[6] & input_a[4];
  assign popcount32_lqzk_core_135 = input_a[14] & input_a[13];
  assign popcount32_lqzk_core_136 = popcount32_lqzk_core_131 | popcount32_lqzk_core_133;
  assign popcount32_lqzk_core_138 = popcount32_lqzk_core_136 ^ input_a[18];
  assign popcount32_lqzk_core_139 = popcount32_lqzk_core_136 & input_a[18];
  assign popcount32_lqzk_core_142 = ~(input_a[7] & input_a[2]);
  assign popcount32_lqzk_core_143 = popcount32_lqzk_core_125 ^ popcount32_lqzk_core_138;
  assign popcount32_lqzk_core_144 = input_a[19] & popcount32_lqzk_core_138;
  assign popcount32_lqzk_core_145 = popcount32_lqzk_core_143 ^ input_a[22];
  assign popcount32_lqzk_core_146 = popcount32_lqzk_core_143 & input_a[22];
  assign popcount32_lqzk_core_147 = popcount32_lqzk_core_144 | popcount32_lqzk_core_146;
  assign popcount32_lqzk_core_149 = input_a[16] ^ input_a[29];
  assign popcount32_lqzk_core_150 = popcount32_lqzk_core_139 | popcount32_lqzk_core_147;
  assign popcount32_lqzk_core_151 = ~(input_a[17] ^ input_a[15]);
  assign popcount32_lqzk_core_153 = input_a[23] | input_a[10];
  assign popcount32_lqzk_core_154 = input_a[24] & input_a[17];
  assign popcount32_lqzk_core_155 = ~(input_a[27] | input_a[10]);
  assign popcount32_lqzk_core_156 = input_a[5] & input_a[7];
  assign popcount32_lqzk_core_157_not = ~input_a[2];
  assign popcount32_lqzk_core_158 = input_a[26] & input_a[10];
  assign popcount32_lqzk_core_159 = popcount32_lqzk_core_154 | popcount32_lqzk_core_156;
  assign popcount32_lqzk_core_161 = popcount32_lqzk_core_159 | popcount32_lqzk_core_158;
  assign popcount32_lqzk_core_162 = input_a[20] ^ input_a[10];
  assign popcount32_lqzk_core_164 = ~(input_a[10] & input_a[13]);
  assign popcount32_lqzk_core_165 = ~(input_a[15] ^ input_a[12]);
  assign popcount32_lqzk_core_167 = ~(input_a[31] ^ input_a[2]);
  assign popcount32_lqzk_core_169 = input_a[16] & input_a[17];
  assign popcount32_lqzk_core_171 = input_a[25] | input_a[13];
  assign popcount32_lqzk_core_172 = input_a[2] | input_a[29];
  assign popcount32_lqzk_core_173 = input_a[14] ^ input_a[1];
  assign popcount32_lqzk_core_176 = input_a[12] | input_a[2];
  assign popcount32_lqzk_core_177 = popcount32_lqzk_core_161 ^ popcount32_lqzk_core_172;
  assign popcount32_lqzk_core_178 = popcount32_lqzk_core_161 & popcount32_lqzk_core_172;
  assign popcount32_lqzk_core_180 = input_a[4] ^ input_a[18];
  assign popcount32_lqzk_core_183 = ~(input_a[23] ^ input_a[2]);
  assign popcount32_lqzk_core_185_not = ~input_a[23];
  assign popcount32_lqzk_core_186 = ~(input_a[3] & input_a[22]);
  assign popcount32_lqzk_core_188 = input_a[0] & input_a[12];
  assign popcount32_lqzk_core_189 = popcount32_lqzk_core_145 ^ popcount32_lqzk_core_177;
  assign popcount32_lqzk_core_190 = popcount32_lqzk_core_145 & popcount32_lqzk_core_177;
  assign popcount32_lqzk_core_191 = popcount32_lqzk_core_189 ^ popcount32_lqzk_core_188;
  assign popcount32_lqzk_core_192 = popcount32_lqzk_core_189 & popcount32_lqzk_core_188;
  assign popcount32_lqzk_core_193 = popcount32_lqzk_core_190 | popcount32_lqzk_core_192;
  assign popcount32_lqzk_core_194 = popcount32_lqzk_core_150 ^ popcount32_lqzk_core_178;
  assign popcount32_lqzk_core_195 = popcount32_lqzk_core_150 & popcount32_lqzk_core_178;
  assign popcount32_lqzk_core_196 = popcount32_lqzk_core_194 ^ popcount32_lqzk_core_193;
  assign popcount32_lqzk_core_197 = popcount32_lqzk_core_194 & popcount32_lqzk_core_193;
  assign popcount32_lqzk_core_198 = popcount32_lqzk_core_195 | popcount32_lqzk_core_197;
  assign popcount32_lqzk_core_200 = ~input_a[8];
  assign popcount32_lqzk_core_202 = ~(input_a[10] & input_a[23]);
  assign popcount32_lqzk_core_203 = input_a[17] & input_a[23];
  assign popcount32_lqzk_core_204 = input_a[14] | input_a[15];
  assign popcount32_lqzk_core_205 = input_a[28] & input_a[9];
  assign popcount32_lqzk_core_206 = popcount32_lqzk_core_106 ^ popcount32_lqzk_core_191;
  assign popcount32_lqzk_core_207 = popcount32_lqzk_core_106 & popcount32_lqzk_core_191;
  assign popcount32_lqzk_core_208 = popcount32_lqzk_core_206 ^ popcount32_lqzk_core_205;
  assign popcount32_lqzk_core_209 = popcount32_lqzk_core_206 & popcount32_lqzk_core_205;
  assign popcount32_lqzk_core_210 = popcount32_lqzk_core_207 | popcount32_lqzk_core_209;
  assign popcount32_lqzk_core_211 = popcount32_lqzk_core_111 ^ popcount32_lqzk_core_196;
  assign popcount32_lqzk_core_212 = popcount32_lqzk_core_111 & popcount32_lqzk_core_196;
  assign popcount32_lqzk_core_213 = popcount32_lqzk_core_211 ^ popcount32_lqzk_core_210;
  assign popcount32_lqzk_core_214 = popcount32_lqzk_core_211 & popcount32_lqzk_core_210;
  assign popcount32_lqzk_core_215 = popcount32_lqzk_core_212 | popcount32_lqzk_core_214;
  assign popcount32_lqzk_core_216 = popcount32_lqzk_core_113 ^ popcount32_lqzk_core_198;
  assign popcount32_lqzk_core_217 = popcount32_lqzk_core_113 & popcount32_lqzk_core_198;
  assign popcount32_lqzk_core_218 = popcount32_lqzk_core_216 ^ popcount32_lqzk_core_215;
  assign popcount32_lqzk_core_219 = popcount32_lqzk_core_216 & popcount32_lqzk_core_215;
  assign popcount32_lqzk_core_220 = popcount32_lqzk_core_217 | popcount32_lqzk_core_219;
  assign popcount32_lqzk_core_221 = ~(input_a[12] ^ input_a[21]);
  assign popcount32_lqzk_core_223 = ~input_a[24];
  assign popcount32_lqzk_core_225 = input_a[3] | input_a[12];

  assign popcount32_lqzk_out[0] = popcount32_lqzk_core_218;
  assign popcount32_lqzk_out[1] = popcount32_lqzk_core_208;
  assign popcount32_lqzk_out[2] = popcount32_lqzk_core_213;
  assign popcount32_lqzk_out[3] = popcount32_lqzk_core_218;
  assign popcount32_lqzk_out[4] = popcount32_lqzk_core_220;
  assign popcount32_lqzk_out[5] = 1'b0;
endmodule