// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5091
// WCE=46.0
// EP=0.996364%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount47_oyl3(input [46:0] input_a, output [5:0] popcount47_oyl3_out);
  wire popcount47_oyl3_core_049;
  wire popcount47_oyl3_core_051;
  wire popcount47_oyl3_core_054;
  wire popcount47_oyl3_core_055;
  wire popcount47_oyl3_core_056;
  wire popcount47_oyl3_core_058;
  wire popcount47_oyl3_core_059;
  wire popcount47_oyl3_core_062;
  wire popcount47_oyl3_core_065;
  wire popcount47_oyl3_core_067;
  wire popcount47_oyl3_core_068;
  wire popcount47_oyl3_core_069;
  wire popcount47_oyl3_core_071;
  wire popcount47_oyl3_core_072;
  wire popcount47_oyl3_core_074;
  wire popcount47_oyl3_core_075;
  wire popcount47_oyl3_core_077;
  wire popcount47_oyl3_core_078;
  wire popcount47_oyl3_core_079;
  wire popcount47_oyl3_core_080;
  wire popcount47_oyl3_core_081;
  wire popcount47_oyl3_core_084;
  wire popcount47_oyl3_core_085;
  wire popcount47_oyl3_core_086;
  wire popcount47_oyl3_core_087;
  wire popcount47_oyl3_core_088;
  wire popcount47_oyl3_core_090;
  wire popcount47_oyl3_core_091;
  wire popcount47_oyl3_core_092;
  wire popcount47_oyl3_core_093;
  wire popcount47_oyl3_core_097;
  wire popcount47_oyl3_core_100;
  wire popcount47_oyl3_core_101;
  wire popcount47_oyl3_core_102;
  wire popcount47_oyl3_core_103;
  wire popcount47_oyl3_core_106;
  wire popcount47_oyl3_core_108;
  wire popcount47_oyl3_core_109;
  wire popcount47_oyl3_core_110;
  wire popcount47_oyl3_core_111;
  wire popcount47_oyl3_core_112;
  wire popcount47_oyl3_core_113;
  wire popcount47_oyl3_core_114;
  wire popcount47_oyl3_core_115;
  wire popcount47_oyl3_core_116;
  wire popcount47_oyl3_core_117;
  wire popcount47_oyl3_core_119;
  wire popcount47_oyl3_core_120;
  wire popcount47_oyl3_core_121;
  wire popcount47_oyl3_core_122;
  wire popcount47_oyl3_core_123;
  wire popcount47_oyl3_core_124;
  wire popcount47_oyl3_core_125;
  wire popcount47_oyl3_core_127;
  wire popcount47_oyl3_core_129;
  wire popcount47_oyl3_core_130;
  wire popcount47_oyl3_core_131;
  wire popcount47_oyl3_core_132;
  wire popcount47_oyl3_core_133;
  wire popcount47_oyl3_core_134;
  wire popcount47_oyl3_core_135;
  wire popcount47_oyl3_core_137;
  wire popcount47_oyl3_core_138;
  wire popcount47_oyl3_core_139;
  wire popcount47_oyl3_core_140;
  wire popcount47_oyl3_core_142;
  wire popcount47_oyl3_core_143;
  wire popcount47_oyl3_core_144;
  wire popcount47_oyl3_core_145;
  wire popcount47_oyl3_core_147;
  wire popcount47_oyl3_core_148;
  wire popcount47_oyl3_core_150;
  wire popcount47_oyl3_core_151;
  wire popcount47_oyl3_core_155;
  wire popcount47_oyl3_core_158;
  wire popcount47_oyl3_core_159_not;
  wire popcount47_oyl3_core_160;
  wire popcount47_oyl3_core_162;
  wire popcount47_oyl3_core_164;
  wire popcount47_oyl3_core_165;
  wire popcount47_oyl3_core_167;
  wire popcount47_oyl3_core_168;
  wire popcount47_oyl3_core_169;
  wire popcount47_oyl3_core_171;
  wire popcount47_oyl3_core_173;
  wire popcount47_oyl3_core_174;
  wire popcount47_oyl3_core_176;
  wire popcount47_oyl3_core_177;
  wire popcount47_oyl3_core_178;
  wire popcount47_oyl3_core_179;
  wire popcount47_oyl3_core_180;
  wire popcount47_oyl3_core_181;
  wire popcount47_oyl3_core_183;
  wire popcount47_oyl3_core_184;
  wire popcount47_oyl3_core_185;
  wire popcount47_oyl3_core_186;
  wire popcount47_oyl3_core_187;
  wire popcount47_oyl3_core_191;
  wire popcount47_oyl3_core_192;
  wire popcount47_oyl3_core_193;
  wire popcount47_oyl3_core_194;
  wire popcount47_oyl3_core_198;
  wire popcount47_oyl3_core_199;
  wire popcount47_oyl3_core_200;
  wire popcount47_oyl3_core_201;
  wire popcount47_oyl3_core_204;
  wire popcount47_oyl3_core_205;
  wire popcount47_oyl3_core_207;
  wire popcount47_oyl3_core_213;
  wire popcount47_oyl3_core_215;
  wire popcount47_oyl3_core_217;
  wire popcount47_oyl3_core_218;
  wire popcount47_oyl3_core_219;
  wire popcount47_oyl3_core_220;
  wire popcount47_oyl3_core_222;
  wire popcount47_oyl3_core_224;
  wire popcount47_oyl3_core_226;
  wire popcount47_oyl3_core_227;
  wire popcount47_oyl3_core_228;
  wire popcount47_oyl3_core_229;
  wire popcount47_oyl3_core_231;
  wire popcount47_oyl3_core_234_not;
  wire popcount47_oyl3_core_235;
  wire popcount47_oyl3_core_236;
  wire popcount47_oyl3_core_237;
  wire popcount47_oyl3_core_238;
  wire popcount47_oyl3_core_239;
  wire popcount47_oyl3_core_242;
  wire popcount47_oyl3_core_244;
  wire popcount47_oyl3_core_245;
  wire popcount47_oyl3_core_246;
  wire popcount47_oyl3_core_250;
  wire popcount47_oyl3_core_252;
  wire popcount47_oyl3_core_253;
  wire popcount47_oyl3_core_254;
  wire popcount47_oyl3_core_255;
  wire popcount47_oyl3_core_256;
  wire popcount47_oyl3_core_257;
  wire popcount47_oyl3_core_258;
  wire popcount47_oyl3_core_260;
  wire popcount47_oyl3_core_261;
  wire popcount47_oyl3_core_262;
  wire popcount47_oyl3_core_263;
  wire popcount47_oyl3_core_264;
  wire popcount47_oyl3_core_265;
  wire popcount47_oyl3_core_266;
  wire popcount47_oyl3_core_267;
  wire popcount47_oyl3_core_268;
  wire popcount47_oyl3_core_270;
  wire popcount47_oyl3_core_276;
  wire popcount47_oyl3_core_277;
  wire popcount47_oyl3_core_278_not;
  wire popcount47_oyl3_core_279;
  wire popcount47_oyl3_core_281;
  wire popcount47_oyl3_core_283;
  wire popcount47_oyl3_core_284;
  wire popcount47_oyl3_core_285;
  wire popcount47_oyl3_core_286;
  wire popcount47_oyl3_core_289_not;
  wire popcount47_oyl3_core_290;
  wire popcount47_oyl3_core_291;
  wire popcount47_oyl3_core_292;
  wire popcount47_oyl3_core_293;
  wire popcount47_oyl3_core_294;
  wire popcount47_oyl3_core_295;
  wire popcount47_oyl3_core_296;
  wire popcount47_oyl3_core_297;
  wire popcount47_oyl3_core_298;
  wire popcount47_oyl3_core_299;
  wire popcount47_oyl3_core_300;
  wire popcount47_oyl3_core_302;
  wire popcount47_oyl3_core_303;
  wire popcount47_oyl3_core_305;
  wire popcount47_oyl3_core_307;
  wire popcount47_oyl3_core_308;
  wire popcount47_oyl3_core_310;
  wire popcount47_oyl3_core_313_not;
  wire popcount47_oyl3_core_315;
  wire popcount47_oyl3_core_316;
  wire popcount47_oyl3_core_317;
  wire popcount47_oyl3_core_318;
  wire popcount47_oyl3_core_321;
  wire popcount47_oyl3_core_322;
  wire popcount47_oyl3_core_323;
  wire popcount47_oyl3_core_324;
  wire popcount47_oyl3_core_325;
  wire popcount47_oyl3_core_326;
  wire popcount47_oyl3_core_328;
  wire popcount47_oyl3_core_330;
  wire popcount47_oyl3_core_333;
  wire popcount47_oyl3_core_334;
  wire popcount47_oyl3_core_336;
  wire popcount47_oyl3_core_337;
  wire popcount47_oyl3_core_345;
  wire popcount47_oyl3_core_347;
  wire popcount47_oyl3_core_349;
  wire popcount47_oyl3_core_350;
  wire popcount47_oyl3_core_352;
  wire popcount47_oyl3_core_353;
  wire popcount47_oyl3_core_354;
  wire popcount47_oyl3_core_355;
  wire popcount47_oyl3_core_356;
  wire popcount47_oyl3_core_359;
  wire popcount47_oyl3_core_360;
  wire popcount47_oyl3_core_362;
  wire popcount47_oyl3_core_363;
  wire popcount47_oyl3_core_364;
  wire popcount47_oyl3_core_365;
  wire popcount47_oyl3_core_366;
  wire popcount47_oyl3_core_367;
  wire popcount47_oyl3_core_368;
  wire popcount47_oyl3_core_370;
  wire popcount47_oyl3_core_372;

  assign popcount47_oyl3_core_049 = ~(input_a[29] | input_a[16]);
  assign popcount47_oyl3_core_051 = ~(input_a[26] | input_a[1]);
  assign popcount47_oyl3_core_054 = ~input_a[41];
  assign popcount47_oyl3_core_055 = ~input_a[37];
  assign popcount47_oyl3_core_056 = input_a[36] | input_a[5];
  assign popcount47_oyl3_core_058 = input_a[19] ^ input_a[29];
  assign popcount47_oyl3_core_059 = input_a[13] & input_a[3];
  assign popcount47_oyl3_core_062 = input_a[38] | input_a[6];
  assign popcount47_oyl3_core_065 = input_a[35] & input_a[41];
  assign popcount47_oyl3_core_067 = input_a[46] | input_a[15];
  assign popcount47_oyl3_core_068 = input_a[46] | input_a[17];
  assign popcount47_oyl3_core_069 = input_a[20] ^ input_a[4];
  assign popcount47_oyl3_core_071 = input_a[1] & input_a[11];
  assign popcount47_oyl3_core_072 = ~input_a[8];
  assign popcount47_oyl3_core_074 = input_a[36] & input_a[17];
  assign popcount47_oyl3_core_075 = ~(input_a[18] | input_a[1]);
  assign popcount47_oyl3_core_077 = ~input_a[4];
  assign popcount47_oyl3_core_078 = ~(input_a[1] ^ input_a[14]);
  assign popcount47_oyl3_core_079 = ~(input_a[10] & input_a[2]);
  assign popcount47_oyl3_core_080 = ~(input_a[2] ^ input_a[2]);
  assign popcount47_oyl3_core_081 = ~(input_a[37] ^ input_a[17]);
  assign popcount47_oyl3_core_084 = input_a[16] & input_a[4];
  assign popcount47_oyl3_core_085 = ~(input_a[9] & input_a[35]);
  assign popcount47_oyl3_core_086 = input_a[29] | input_a[35];
  assign popcount47_oyl3_core_087 = ~input_a[9];
  assign popcount47_oyl3_core_088 = ~input_a[31];
  assign popcount47_oyl3_core_090 = ~input_a[1];
  assign popcount47_oyl3_core_091 = ~(input_a[31] ^ input_a[24]);
  assign popcount47_oyl3_core_092 = input_a[36] & input_a[39];
  assign popcount47_oyl3_core_093 = ~(input_a[8] | input_a[39]);
  assign popcount47_oyl3_core_097 = ~(input_a[6] | input_a[32]);
  assign popcount47_oyl3_core_100 = ~(input_a[21] | input_a[6]);
  assign popcount47_oyl3_core_101 = ~input_a[26];
  assign popcount47_oyl3_core_102 = ~(input_a[11] | input_a[35]);
  assign popcount47_oyl3_core_103 = input_a[39] & input_a[26];
  assign popcount47_oyl3_core_106 = ~(input_a[43] & input_a[31]);
  assign popcount47_oyl3_core_108 = input_a[42] | input_a[11];
  assign popcount47_oyl3_core_109 = ~input_a[23];
  assign popcount47_oyl3_core_110 = ~input_a[14];
  assign popcount47_oyl3_core_111 = input_a[0] | input_a[33];
  assign popcount47_oyl3_core_112 = ~input_a[17];
  assign popcount47_oyl3_core_113 = ~(input_a[38] & input_a[18]);
  assign popcount47_oyl3_core_114 = ~input_a[34];
  assign popcount47_oyl3_core_115 = ~input_a[19];
  assign popcount47_oyl3_core_116 = input_a[9] | input_a[44];
  assign popcount47_oyl3_core_117 = ~input_a[30];
  assign popcount47_oyl3_core_119 = ~input_a[17];
  assign popcount47_oyl3_core_120 = input_a[11] ^ input_a[18];
  assign popcount47_oyl3_core_121 = ~(input_a[18] & input_a[44]);
  assign popcount47_oyl3_core_122 = ~(input_a[32] ^ input_a[4]);
  assign popcount47_oyl3_core_123 = ~(input_a[34] | input_a[29]);
  assign popcount47_oyl3_core_124 = ~(input_a[30] | input_a[31]);
  assign popcount47_oyl3_core_125 = input_a[45] ^ input_a[1];
  assign popcount47_oyl3_core_127 = input_a[44] & input_a[2];
  assign popcount47_oyl3_core_129 = input_a[45] ^ input_a[43];
  assign popcount47_oyl3_core_130 = input_a[22] & input_a[6];
  assign popcount47_oyl3_core_131 = input_a[41] ^ input_a[14];
  assign popcount47_oyl3_core_132 = ~input_a[16];
  assign popcount47_oyl3_core_133 = ~(input_a[29] & input_a[5]);
  assign popcount47_oyl3_core_134 = input_a[35] ^ input_a[23];
  assign popcount47_oyl3_core_135 = ~(input_a[6] ^ input_a[37]);
  assign popcount47_oyl3_core_137 = ~(input_a[28] ^ input_a[1]);
  assign popcount47_oyl3_core_138 = ~(input_a[27] | input_a[1]);
  assign popcount47_oyl3_core_139 = input_a[5] ^ input_a[27];
  assign popcount47_oyl3_core_140 = input_a[13] ^ input_a[44];
  assign popcount47_oyl3_core_142 = ~(input_a[29] & input_a[5]);
  assign popcount47_oyl3_core_143 = ~(input_a[24] ^ input_a[12]);
  assign popcount47_oyl3_core_144 = ~(input_a[7] | input_a[17]);
  assign popcount47_oyl3_core_145 = input_a[36] | input_a[35];
  assign popcount47_oyl3_core_147 = ~(input_a[32] & input_a[1]);
  assign popcount47_oyl3_core_148 = input_a[21] & input_a[15];
  assign popcount47_oyl3_core_150 = input_a[23] & input_a[23];
  assign popcount47_oyl3_core_151 = ~(input_a[18] ^ input_a[45]);
  assign popcount47_oyl3_core_155 = ~(input_a[29] ^ input_a[1]);
  assign popcount47_oyl3_core_158 = input_a[35] & input_a[26];
  assign popcount47_oyl3_core_159_not = ~input_a[15];
  assign popcount47_oyl3_core_160 = ~(input_a[13] | input_a[14]);
  assign popcount47_oyl3_core_162 = ~input_a[9];
  assign popcount47_oyl3_core_164 = input_a[26] | input_a[2];
  assign popcount47_oyl3_core_165 = input_a[32] & input_a[30];
  assign popcount47_oyl3_core_167 = ~(input_a[13] & input_a[24]);
  assign popcount47_oyl3_core_168 = ~input_a[0];
  assign popcount47_oyl3_core_169 = ~(input_a[8] ^ input_a[45]);
  assign popcount47_oyl3_core_171 = ~(input_a[11] | input_a[18]);
  assign popcount47_oyl3_core_173 = input_a[14] ^ input_a[43];
  assign popcount47_oyl3_core_174 = input_a[9] & input_a[11];
  assign popcount47_oyl3_core_176 = input_a[7] & input_a[43];
  assign popcount47_oyl3_core_177 = input_a[11] & input_a[13];
  assign popcount47_oyl3_core_178 = ~(input_a[7] | input_a[2]);
  assign popcount47_oyl3_core_179 = input_a[8] | input_a[11];
  assign popcount47_oyl3_core_180 = ~(input_a[34] | input_a[5]);
  assign popcount47_oyl3_core_181 = input_a[10] & input_a[37];
  assign popcount47_oyl3_core_183 = input_a[9] & input_a[15];
  assign popcount47_oyl3_core_184 = ~(input_a[30] ^ input_a[28]);
  assign popcount47_oyl3_core_185 = ~input_a[12];
  assign popcount47_oyl3_core_186 = ~(input_a[13] & input_a[45]);
  assign popcount47_oyl3_core_187 = ~(input_a[9] ^ input_a[16]);
  assign popcount47_oyl3_core_191 = ~input_a[32];
  assign popcount47_oyl3_core_192 = ~input_a[5];
  assign popcount47_oyl3_core_193 = input_a[12] | input_a[3];
  assign popcount47_oyl3_core_194 = input_a[34] & input_a[13];
  assign popcount47_oyl3_core_198 = ~input_a[24];
  assign popcount47_oyl3_core_199 = input_a[24] & input_a[26];
  assign popcount47_oyl3_core_200 = input_a[32] | input_a[27];
  assign popcount47_oyl3_core_201 = input_a[19] & input_a[10];
  assign popcount47_oyl3_core_204 = ~input_a[28];
  assign popcount47_oyl3_core_205 = input_a[14] & input_a[0];
  assign popcount47_oyl3_core_207 = ~(input_a[33] & input_a[12]);
  assign popcount47_oyl3_core_213 = ~(input_a[34] | input_a[41]);
  assign popcount47_oyl3_core_215 = ~(input_a[45] ^ input_a[2]);
  assign popcount47_oyl3_core_217 = input_a[29] | input_a[13];
  assign popcount47_oyl3_core_218 = input_a[44] | input_a[38];
  assign popcount47_oyl3_core_219 = ~(input_a[24] & input_a[18]);
  assign popcount47_oyl3_core_220 = ~(input_a[8] ^ input_a[10]);
  assign popcount47_oyl3_core_222 = ~(input_a[22] & input_a[4]);
  assign popcount47_oyl3_core_224 = ~(input_a[16] & input_a[21]);
  assign popcount47_oyl3_core_226 = ~(input_a[26] & input_a[24]);
  assign popcount47_oyl3_core_227 = input_a[5] | input_a[42];
  assign popcount47_oyl3_core_228 = ~(input_a[37] ^ input_a[29]);
  assign popcount47_oyl3_core_229 = input_a[17] ^ input_a[28];
  assign popcount47_oyl3_core_231 = input_a[15] & input_a[43];
  assign popcount47_oyl3_core_234_not = ~input_a[12];
  assign popcount47_oyl3_core_235 = ~(input_a[29] & input_a[5]);
  assign popcount47_oyl3_core_236 = ~(input_a[45] & input_a[32]);
  assign popcount47_oyl3_core_237 = input_a[16] & input_a[2];
  assign popcount47_oyl3_core_238 = ~(input_a[6] & input_a[38]);
  assign popcount47_oyl3_core_239 = ~input_a[6];
  assign popcount47_oyl3_core_242 = ~(input_a[19] & input_a[44]);
  assign popcount47_oyl3_core_244 = ~input_a[10];
  assign popcount47_oyl3_core_245 = input_a[6] & input_a[14];
  assign popcount47_oyl3_core_246 = input_a[39] ^ input_a[45];
  assign popcount47_oyl3_core_250 = input_a[24] | input_a[28];
  assign popcount47_oyl3_core_252 = input_a[40] ^ input_a[1];
  assign popcount47_oyl3_core_253 = ~(input_a[32] ^ input_a[24]);
  assign popcount47_oyl3_core_254 = input_a[43] | input_a[12];
  assign popcount47_oyl3_core_255 = ~(input_a[41] | input_a[42]);
  assign popcount47_oyl3_core_256 = input_a[5] & input_a[12];
  assign popcount47_oyl3_core_257 = ~input_a[22];
  assign popcount47_oyl3_core_258 = input_a[4] | input_a[8];
  assign popcount47_oyl3_core_260 = ~input_a[41];
  assign popcount47_oyl3_core_261 = ~(input_a[33] ^ input_a[14]);
  assign popcount47_oyl3_core_262 = ~input_a[32];
  assign popcount47_oyl3_core_263 = input_a[9] ^ input_a[5];
  assign popcount47_oyl3_core_264 = ~(input_a[34] | input_a[43]);
  assign popcount47_oyl3_core_265 = input_a[23] | input_a[13];
  assign popcount47_oyl3_core_266 = ~(input_a[34] & input_a[25]);
  assign popcount47_oyl3_core_267 = input_a[17] | input_a[12];
  assign popcount47_oyl3_core_268 = input_a[27] & input_a[44];
  assign popcount47_oyl3_core_270 = ~(input_a[19] & input_a[28]);
  assign popcount47_oyl3_core_276 = input_a[19] | input_a[18];
  assign popcount47_oyl3_core_277 = ~(input_a[29] | input_a[29]);
  assign popcount47_oyl3_core_278_not = ~input_a[13];
  assign popcount47_oyl3_core_279 = ~(input_a[5] ^ input_a[20]);
  assign popcount47_oyl3_core_281 = ~input_a[15];
  assign popcount47_oyl3_core_283 = input_a[12] | input_a[23];
  assign popcount47_oyl3_core_284 = input_a[31] | input_a[34];
  assign popcount47_oyl3_core_285 = ~(input_a[34] & input_a[28]);
  assign popcount47_oyl3_core_286 = input_a[46] ^ input_a[16];
  assign popcount47_oyl3_core_289_not = ~input_a[40];
  assign popcount47_oyl3_core_290 = input_a[23] | input_a[30];
  assign popcount47_oyl3_core_291 = ~(input_a[32] ^ input_a[46]);
  assign popcount47_oyl3_core_292 = input_a[20] & input_a[39];
  assign popcount47_oyl3_core_293 = ~(input_a[10] ^ input_a[4]);
  assign popcount47_oyl3_core_294 = ~(input_a[25] | input_a[1]);
  assign popcount47_oyl3_core_295 = ~(input_a[36] | input_a[13]);
  assign popcount47_oyl3_core_296 = ~(input_a[24] & input_a[15]);
  assign popcount47_oyl3_core_297 = ~(input_a[44] | input_a[21]);
  assign popcount47_oyl3_core_298 = ~(input_a[16] ^ input_a[14]);
  assign popcount47_oyl3_core_299 = ~(input_a[26] ^ input_a[40]);
  assign popcount47_oyl3_core_300 = input_a[43] & input_a[8];
  assign popcount47_oyl3_core_302 = input_a[35] & input_a[41];
  assign popcount47_oyl3_core_303 = ~(input_a[22] | input_a[15]);
  assign popcount47_oyl3_core_305 = ~(input_a[34] ^ input_a[14]);
  assign popcount47_oyl3_core_307 = ~(input_a[15] | input_a[24]);
  assign popcount47_oyl3_core_308 = ~input_a[14];
  assign popcount47_oyl3_core_310 = ~(input_a[27] ^ input_a[6]);
  assign popcount47_oyl3_core_313_not = ~input_a[7];
  assign popcount47_oyl3_core_315 = ~input_a[32];
  assign popcount47_oyl3_core_316 = input_a[2] & input_a[16];
  assign popcount47_oyl3_core_317 = ~(input_a[44] & input_a[36]);
  assign popcount47_oyl3_core_318 = ~(input_a[17] ^ input_a[45]);
  assign popcount47_oyl3_core_321 = ~input_a[25];
  assign popcount47_oyl3_core_322 = ~input_a[20];
  assign popcount47_oyl3_core_323 = input_a[18] & input_a[40];
  assign popcount47_oyl3_core_324 = input_a[13] & input_a[4];
  assign popcount47_oyl3_core_325 = input_a[36] & input_a[6];
  assign popcount47_oyl3_core_326 = input_a[39] | input_a[26];
  assign popcount47_oyl3_core_328 = input_a[17] & input_a[44];
  assign popcount47_oyl3_core_330 = input_a[41] & input_a[9];
  assign popcount47_oyl3_core_333 = input_a[25] | input_a[2];
  assign popcount47_oyl3_core_334 = input_a[5] & input_a[37];
  assign popcount47_oyl3_core_336 = ~(input_a[14] ^ input_a[23]);
  assign popcount47_oyl3_core_337 = ~(input_a[8] | input_a[41]);
  assign popcount47_oyl3_core_345 = ~(input_a[4] ^ input_a[16]);
  assign popcount47_oyl3_core_347 = ~(input_a[0] | input_a[36]);
  assign popcount47_oyl3_core_349 = input_a[2] ^ input_a[33];
  assign popcount47_oyl3_core_350 = ~(input_a[12] & input_a[13]);
  assign popcount47_oyl3_core_352 = input_a[28] & input_a[43];
  assign popcount47_oyl3_core_353 = input_a[22] ^ input_a[29];
  assign popcount47_oyl3_core_354 = input_a[15] & input_a[40];
  assign popcount47_oyl3_core_355 = ~input_a[32];
  assign popcount47_oyl3_core_356 = ~(input_a[38] | input_a[0]);
  assign popcount47_oyl3_core_359 = ~input_a[35];
  assign popcount47_oyl3_core_360 = ~(input_a[15] ^ input_a[36]);
  assign popcount47_oyl3_core_362 = ~input_a[12];
  assign popcount47_oyl3_core_363 = input_a[27] ^ input_a[16];
  assign popcount47_oyl3_core_364 = input_a[39] ^ input_a[3];
  assign popcount47_oyl3_core_365 = ~(input_a[44] | input_a[37]);
  assign popcount47_oyl3_core_366 = input_a[6] | input_a[28];
  assign popcount47_oyl3_core_367 = ~(input_a[41] | input_a[1]);
  assign popcount47_oyl3_core_368 = ~input_a[15];
  assign popcount47_oyl3_core_370 = input_a[4] | input_a[5];
  assign popcount47_oyl3_core_372 = ~(input_a[27] & input_a[23]);

  assign popcount47_oyl3_out[0] = 1'b0;
  assign popcount47_oyl3_out[1] = 1'b0;
  assign popcount47_oyl3_out[2] = 1'b0;
  assign popcount47_oyl3_out[3] = 1'b0;
  assign popcount47_oyl3_out[4] = input_a[36];
  assign popcount47_oyl3_out[5] = input_a[23];
endmodule