// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.44912
// WCE=17.0
// EP=0.872399%
// Printed PDK parameters:
//  Area=627920.0
//  Delay=2618200.0
//  Power=30372.0

module popcount34_q4e0(input [33:0] input_a, output [5:0] popcount34_q4e0_out);
  wire popcount34_q4e0_core_036;
  wire popcount34_q4e0_core_037;
  wire popcount34_q4e0_core_038;
  wire popcount34_q4e0_core_039;
  wire popcount34_q4e0_core_040;
  wire popcount34_q4e0_core_041;
  wire popcount34_q4e0_core_042;
  wire popcount34_q4e0_core_044;
  wire popcount34_q4e0_core_045;
  wire popcount34_q4e0_core_049;
  wire popcount34_q4e0_core_050;
  wire popcount34_q4e0_core_052;
  wire popcount34_q4e0_core_055;
  wire popcount34_q4e0_core_057;
  wire popcount34_q4e0_core_058;
  wire popcount34_q4e0_core_061;
  wire popcount34_q4e0_core_062;
  wire popcount34_q4e0_core_064;
  wire popcount34_q4e0_core_066;
  wire popcount34_q4e0_core_067;
  wire popcount34_q4e0_core_068;
  wire popcount34_q4e0_core_070;
  wire popcount34_q4e0_core_071;
  wire popcount34_q4e0_core_074;
  wire popcount34_q4e0_core_075;
  wire popcount34_q4e0_core_077;
  wire popcount34_q4e0_core_078;
  wire popcount34_q4e0_core_079_not;
  wire popcount34_q4e0_core_080;
  wire popcount34_q4e0_core_081;
  wire popcount34_q4e0_core_083_not;
  wire popcount34_q4e0_core_084;
  wire popcount34_q4e0_core_085;
  wire popcount34_q4e0_core_087;
  wire popcount34_q4e0_core_089;
  wire popcount34_q4e0_core_092;
  wire popcount34_q4e0_core_094_not;
  wire popcount34_q4e0_core_096;
  wire popcount34_q4e0_core_097;
  wire popcount34_q4e0_core_098;
  wire popcount34_q4e0_core_101;
  wire popcount34_q4e0_core_102;
  wire popcount34_q4e0_core_103;
  wire popcount34_q4e0_core_104;
  wire popcount34_q4e0_core_105;
  wire popcount34_q4e0_core_106;
  wire popcount34_q4e0_core_107;
  wire popcount34_q4e0_core_109;
  wire popcount34_q4e0_core_111;
  wire popcount34_q4e0_core_112;
  wire popcount34_q4e0_core_114;
  wire popcount34_q4e0_core_115;
  wire popcount34_q4e0_core_116;
  wire popcount34_q4e0_core_117;
  wire popcount34_q4e0_core_119;
  wire popcount34_q4e0_core_121;
  wire popcount34_q4e0_core_122;
  wire popcount34_q4e0_core_125;
  wire popcount34_q4e0_core_127;
  wire popcount34_q4e0_core_128;
  wire popcount34_q4e0_core_130;
  wire popcount34_q4e0_core_132;
  wire popcount34_q4e0_core_133;
  wire popcount34_q4e0_core_139;
  wire popcount34_q4e0_core_140_not;
  wire popcount34_q4e0_core_141;
  wire popcount34_q4e0_core_144;
  wire popcount34_q4e0_core_145;
  wire popcount34_q4e0_core_146;
  wire popcount34_q4e0_core_147;
  wire popcount34_q4e0_core_148;
  wire popcount34_q4e0_core_149_not;
  wire popcount34_q4e0_core_150;
  wire popcount34_q4e0_core_151;
  wire popcount34_q4e0_core_152;
  wire popcount34_q4e0_core_154;
  wire popcount34_q4e0_core_155;
  wire popcount34_q4e0_core_157;
  wire popcount34_q4e0_core_159;
  wire popcount34_q4e0_core_160;
  wire popcount34_q4e0_core_162;
  wire popcount34_q4e0_core_163;
  wire popcount34_q4e0_core_164_not;
  wire popcount34_q4e0_core_166;
  wire popcount34_q4e0_core_167;
  wire popcount34_q4e0_core_168;
  wire popcount34_q4e0_core_169;
  wire popcount34_q4e0_core_170;
  wire popcount34_q4e0_core_172;
  wire popcount34_q4e0_core_173;
  wire popcount34_q4e0_core_174;
  wire popcount34_q4e0_core_176;
  wire popcount34_q4e0_core_177;
  wire popcount34_q4e0_core_178;
  wire popcount34_q4e0_core_180;
  wire popcount34_q4e0_core_181;
  wire popcount34_q4e0_core_182;
  wire popcount34_q4e0_core_185;
  wire popcount34_q4e0_core_186;
  wire popcount34_q4e0_core_187;
  wire popcount34_q4e0_core_189;
  wire popcount34_q4e0_core_191;
  wire popcount34_q4e0_core_192;
  wire popcount34_q4e0_core_193;
  wire popcount34_q4e0_core_194;
  wire popcount34_q4e0_core_195;
  wire popcount34_q4e0_core_196;
  wire popcount34_q4e0_core_200;
  wire popcount34_q4e0_core_202;
  wire popcount34_q4e0_core_203;
  wire popcount34_q4e0_core_204;
  wire popcount34_q4e0_core_205;
  wire popcount34_q4e0_core_209;
  wire popcount34_q4e0_core_210;
  wire popcount34_q4e0_core_211;
  wire popcount34_q4e0_core_212;
  wire popcount34_q4e0_core_214;
  wire popcount34_q4e0_core_215;
  wire popcount34_q4e0_core_216;
  wire popcount34_q4e0_core_218;
  wire popcount34_q4e0_core_219;
  wire popcount34_q4e0_core_220;
  wire popcount34_q4e0_core_224;
  wire popcount34_q4e0_core_225;
  wire popcount34_q4e0_core_227_not;
  wire popcount34_q4e0_core_229;
  wire popcount34_q4e0_core_231;
  wire popcount34_q4e0_core_232;
  wire popcount34_q4e0_core_234;
  wire popcount34_q4e0_core_235;
  wire popcount34_q4e0_core_236_not;
  wire popcount34_q4e0_core_238;
  wire popcount34_q4e0_core_239;
  wire popcount34_q4e0_core_240;
  wire popcount34_q4e0_core_241;
  wire popcount34_q4e0_core_242;
  wire popcount34_q4e0_core_243;
  wire popcount34_q4e0_core_244;
  wire popcount34_q4e0_core_246;
  wire popcount34_q4e0_core_247;
  wire popcount34_q4e0_core_249;
  wire popcount34_q4e0_core_250;
  wire popcount34_q4e0_core_252;

  assign popcount34_q4e0_core_036 = ~input_a[27];
  assign popcount34_q4e0_core_037 = input_a[16] | input_a[29];
  assign popcount34_q4e0_core_038 = ~(input_a[26] | input_a[16]);
  assign popcount34_q4e0_core_039 = ~(input_a[24] ^ input_a[25]);
  assign popcount34_q4e0_core_040 = ~(input_a[24] & input_a[21]);
  assign popcount34_q4e0_core_041 = input_a[6] & input_a[27];
  assign popcount34_q4e0_core_042 = ~input_a[4];
  assign popcount34_q4e0_core_044 = input_a[10] ^ input_a[31];
  assign popcount34_q4e0_core_045 = ~(input_a[5] & input_a[30]);
  assign popcount34_q4e0_core_049 = ~input_a[10];
  assign popcount34_q4e0_core_050 = input_a[28] | input_a[3];
  assign popcount34_q4e0_core_052 = ~input_a[26];
  assign popcount34_q4e0_core_055 = ~(input_a[20] | input_a[30]);
  assign popcount34_q4e0_core_057 = input_a[22] | input_a[25];
  assign popcount34_q4e0_core_058 = ~(input_a[14] | input_a[4]);
  assign popcount34_q4e0_core_061 = ~(input_a[32] | input_a[20]);
  assign popcount34_q4e0_core_062 = ~input_a[12];
  assign popcount34_q4e0_core_064 = ~(input_a[1] ^ input_a[21]);
  assign popcount34_q4e0_core_066 = input_a[25] & input_a[23];
  assign popcount34_q4e0_core_067 = ~input_a[22];
  assign popcount34_q4e0_core_068 = input_a[31] & input_a[1];
  assign popcount34_q4e0_core_070 = input_a[16] | input_a[27];
  assign popcount34_q4e0_core_071 = input_a[32] & input_a[10];
  assign popcount34_q4e0_core_074 = ~(input_a[12] ^ input_a[24]);
  assign popcount34_q4e0_core_075 = ~(input_a[8] | input_a[13]);
  assign popcount34_q4e0_core_077 = ~input_a[11];
  assign popcount34_q4e0_core_078 = ~(input_a[7] | input_a[31]);
  assign popcount34_q4e0_core_079_not = ~input_a[33];
  assign popcount34_q4e0_core_080 = input_a[31] & input_a[26];
  assign popcount34_q4e0_core_081 = input_a[5] & input_a[0];
  assign popcount34_q4e0_core_083_not = ~input_a[11];
  assign popcount34_q4e0_core_084 = input_a[9] | input_a[15];
  assign popcount34_q4e0_core_085 = input_a[8] & input_a[4];
  assign popcount34_q4e0_core_087 = ~(input_a[8] | input_a[17]);
  assign popcount34_q4e0_core_089 = ~(input_a[1] ^ input_a[1]);
  assign popcount34_q4e0_core_092 = ~input_a[32];
  assign popcount34_q4e0_core_094_not = ~input_a[1];
  assign popcount34_q4e0_core_096 = ~(input_a[24] | input_a[13]);
  assign popcount34_q4e0_core_097 = input_a[8] | input_a[4];
  assign popcount34_q4e0_core_098 = ~(input_a[0] ^ input_a[27]);
  assign popcount34_q4e0_core_101 = input_a[7] ^ input_a[5];
  assign popcount34_q4e0_core_102 = input_a[12] & input_a[17];
  assign popcount34_q4e0_core_103 = ~input_a[6];
  assign popcount34_q4e0_core_104 = ~input_a[26];
  assign popcount34_q4e0_core_105 = ~(input_a[32] ^ input_a[15]);
  assign popcount34_q4e0_core_106 = ~input_a[2];
  assign popcount34_q4e0_core_107 = ~input_a[23];
  assign popcount34_q4e0_core_109 = ~input_a[9];
  assign popcount34_q4e0_core_111 = ~input_a[9];
  assign popcount34_q4e0_core_112 = ~input_a[16];
  assign popcount34_q4e0_core_114 = ~(input_a[13] & input_a[15]);
  assign popcount34_q4e0_core_115 = ~(input_a[13] ^ input_a[2]);
  assign popcount34_q4e0_core_116 = ~(input_a[5] & input_a[23]);
  assign popcount34_q4e0_core_117 = ~(input_a[23] & input_a[6]);
  assign popcount34_q4e0_core_119 = input_a[20] & input_a[0];
  assign popcount34_q4e0_core_121 = ~input_a[7];
  assign popcount34_q4e0_core_122 = ~input_a[27];
  assign popcount34_q4e0_core_125 = ~(input_a[20] ^ input_a[7]);
  assign popcount34_q4e0_core_127 = ~(input_a[4] | input_a[29]);
  assign popcount34_q4e0_core_128 = ~(input_a[25] ^ input_a[31]);
  assign popcount34_q4e0_core_130 = ~(input_a[31] ^ input_a[25]);
  assign popcount34_q4e0_core_132 = ~input_a[28];
  assign popcount34_q4e0_core_133 = ~input_a[28];
  assign popcount34_q4e0_core_139 = ~(input_a[21] & input_a[15]);
  assign popcount34_q4e0_core_140_not = ~input_a[12];
  assign popcount34_q4e0_core_141 = input_a[0] | input_a[0];
  assign popcount34_q4e0_core_144 = ~input_a[10];
  assign popcount34_q4e0_core_145 = input_a[7] | input_a[15];
  assign popcount34_q4e0_core_146 = ~(input_a[4] ^ input_a[7]);
  assign popcount34_q4e0_core_147 = ~(input_a[15] | input_a[31]);
  assign popcount34_q4e0_core_148 = ~(input_a[31] ^ input_a[1]);
  assign popcount34_q4e0_core_149_not = ~input_a[16];
  assign popcount34_q4e0_core_150 = input_a[5] ^ input_a[15];
  assign popcount34_q4e0_core_151 = input_a[16] | input_a[19];
  assign popcount34_q4e0_core_152 = input_a[19] | input_a[33];
  assign popcount34_q4e0_core_154 = ~input_a[11];
  assign popcount34_q4e0_core_155 = ~input_a[8];
  assign popcount34_q4e0_core_157 = ~(input_a[17] & input_a[0]);
  assign popcount34_q4e0_core_159 = ~input_a[32];
  assign popcount34_q4e0_core_160 = ~(input_a[33] & input_a[4]);
  assign popcount34_q4e0_core_162 = input_a[32] | input_a[30];
  assign popcount34_q4e0_core_163 = ~(input_a[4] & input_a[18]);
  assign popcount34_q4e0_core_164_not = ~input_a[30];
  assign popcount34_q4e0_core_166 = ~(input_a[8] & input_a[27]);
  assign popcount34_q4e0_core_167 = input_a[14] | input_a[9];
  assign popcount34_q4e0_core_168 = input_a[15] & input_a[19];
  assign popcount34_q4e0_core_169 = input_a[12] ^ input_a[10];
  assign popcount34_q4e0_core_170 = input_a[20] | input_a[31];
  assign popcount34_q4e0_core_172 = input_a[7] | input_a[2];
  assign popcount34_q4e0_core_173 = input_a[24] | input_a[24];
  assign popcount34_q4e0_core_174 = ~input_a[7];
  assign popcount34_q4e0_core_176 = input_a[26] & input_a[18];
  assign popcount34_q4e0_core_177 = ~(input_a[24] | input_a[26]);
  assign popcount34_q4e0_core_178 = input_a[27] ^ input_a[9];
  assign popcount34_q4e0_core_180 = ~(input_a[21] ^ input_a[14]);
  assign popcount34_q4e0_core_181 = input_a[28] & input_a[13];
  assign popcount34_q4e0_core_182 = ~(input_a[13] | input_a[0]);
  assign popcount34_q4e0_core_185 = input_a[19] & input_a[21];
  assign popcount34_q4e0_core_186 = input_a[10] & input_a[33];
  assign popcount34_q4e0_core_187 = ~(input_a[21] ^ input_a[12]);
  assign popcount34_q4e0_core_189 = ~(input_a[21] & input_a[7]);
  assign popcount34_q4e0_core_191 = input_a[21] | input_a[22];
  assign popcount34_q4e0_core_192 = input_a[13] ^ input_a[26];
  assign popcount34_q4e0_core_193 = input_a[13] ^ input_a[27];
  assign popcount34_q4e0_core_194 = ~(input_a[25] | input_a[2]);
  assign popcount34_q4e0_core_195 = ~input_a[30];
  assign popcount34_q4e0_core_196 = input_a[15] | input_a[2];
  assign popcount34_q4e0_core_200 = input_a[33] | input_a[2];
  assign popcount34_q4e0_core_202 = input_a[16] ^ input_a[12];
  assign popcount34_q4e0_core_203 = ~input_a[5];
  assign popcount34_q4e0_core_204 = input_a[25] & input_a[24];
  assign popcount34_q4e0_core_205 = ~(input_a[27] & input_a[29]);
  assign popcount34_q4e0_core_209 = ~(input_a[20] | input_a[6]);
  assign popcount34_q4e0_core_210 = input_a[18] | input_a[29];
  assign popcount34_q4e0_core_211 = input_a[11] & input_a[17];
  assign popcount34_q4e0_core_212 = ~(input_a[20] & input_a[22]);
  assign popcount34_q4e0_core_214 = input_a[15] ^ input_a[25];
  assign popcount34_q4e0_core_215 = ~(input_a[12] & input_a[11]);
  assign popcount34_q4e0_core_216 = ~input_a[8];
  assign popcount34_q4e0_core_218 = input_a[8] | input_a[17];
  assign popcount34_q4e0_core_219 = input_a[8] | input_a[6];
  assign popcount34_q4e0_core_220 = input_a[28] ^ input_a[10];
  assign popcount34_q4e0_core_224 = ~input_a[17];
  assign popcount34_q4e0_core_225 = ~(input_a[21] & input_a[16]);
  assign popcount34_q4e0_core_227_not = ~input_a[4];
  assign popcount34_q4e0_core_229 = ~(input_a[13] & input_a[22]);
  assign popcount34_q4e0_core_231 = ~input_a[21];
  assign popcount34_q4e0_core_232 = ~input_a[25];
  assign popcount34_q4e0_core_234 = input_a[19] & popcount34_q4e0_core_216;
  assign popcount34_q4e0_core_235 = ~(input_a[0] ^ input_a[5]);
  assign popcount34_q4e0_core_236_not = ~input_a[3];
  assign popcount34_q4e0_core_238 = ~input_a[8];
  assign popcount34_q4e0_core_239 = ~(input_a[16] & input_a[2]);
  assign popcount34_q4e0_core_240 = popcount34_q4e0_core_238 ^ popcount34_q4e0_core_234;
  assign popcount34_q4e0_core_241 = input_a[10] ^ input_a[13];
  assign popcount34_q4e0_core_242 = input_a[8] | input_a[19];
  assign popcount34_q4e0_core_243 = input_a[18] | input_a[32];
  assign popcount34_q4e0_core_244 = input_a[33] ^ input_a[2];
  assign popcount34_q4e0_core_246 = ~(input_a[9] ^ input_a[22]);
  assign popcount34_q4e0_core_247 = input_a[11] | input_a[19];
  assign popcount34_q4e0_core_249 = ~(input_a[8] ^ input_a[2]);
  assign popcount34_q4e0_core_250 = ~input_a[2];
  assign popcount34_q4e0_core_252 = ~input_a[24];

  assign popcount34_q4e0_out[0] = input_a[0];
  assign popcount34_q4e0_out[1] = 1'b1;
  assign popcount34_q4e0_out[2] = popcount34_q4e0_core_240;
  assign popcount34_q4e0_out[3] = popcount34_q4e0_core_240;
  assign popcount34_q4e0_out[4] = popcount34_q4e0_core_242;
  assign popcount34_q4e0_out[5] = 1'b0;
endmodule