// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.01475
// WCE=13.0
// EP=0.845019%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_ikmp(input [24:0] input_a, output [4:0] popcount25_ikmp_out);
  wire popcount25_ikmp_core_027;
  wire popcount25_ikmp_core_028;
  wire popcount25_ikmp_core_030;
  wire popcount25_ikmp_core_032;
  wire popcount25_ikmp_core_033;
  wire popcount25_ikmp_core_036;
  wire popcount25_ikmp_core_037;
  wire popcount25_ikmp_core_038;
  wire popcount25_ikmp_core_039;
  wire popcount25_ikmp_core_040_not;
  wire popcount25_ikmp_core_044;
  wire popcount25_ikmp_core_046;
  wire popcount25_ikmp_core_048;
  wire popcount25_ikmp_core_049;
  wire popcount25_ikmp_core_052;
  wire popcount25_ikmp_core_053;
  wire popcount25_ikmp_core_056;
  wire popcount25_ikmp_core_057;
  wire popcount25_ikmp_core_058_not;
  wire popcount25_ikmp_core_059;
  wire popcount25_ikmp_core_061;
  wire popcount25_ikmp_core_062;
  wire popcount25_ikmp_core_064;
  wire popcount25_ikmp_core_066;
  wire popcount25_ikmp_core_067;
  wire popcount25_ikmp_core_068;
  wire popcount25_ikmp_core_070;
  wire popcount25_ikmp_core_071;
  wire popcount25_ikmp_core_072;
  wire popcount25_ikmp_core_073;
  wire popcount25_ikmp_core_075;
  wire popcount25_ikmp_core_076;
  wire popcount25_ikmp_core_077;
  wire popcount25_ikmp_core_078;
  wire popcount25_ikmp_core_079;
  wire popcount25_ikmp_core_080;
  wire popcount25_ikmp_core_082;
  wire popcount25_ikmp_core_083_not;
  wire popcount25_ikmp_core_089;
  wire popcount25_ikmp_core_093;
  wire popcount25_ikmp_core_094;
  wire popcount25_ikmp_core_095;
  wire popcount25_ikmp_core_096;
  wire popcount25_ikmp_core_097;
  wire popcount25_ikmp_core_098;
  wire popcount25_ikmp_core_099_not;
  wire popcount25_ikmp_core_100;
  wire popcount25_ikmp_core_102;
  wire popcount25_ikmp_core_105;
  wire popcount25_ikmp_core_108;
  wire popcount25_ikmp_core_111;
  wire popcount25_ikmp_core_114;
  wire popcount25_ikmp_core_117;
  wire popcount25_ikmp_core_118;
  wire popcount25_ikmp_core_119;
  wire popcount25_ikmp_core_121;
  wire popcount25_ikmp_core_123;
  wire popcount25_ikmp_core_126;
  wire popcount25_ikmp_core_127;
  wire popcount25_ikmp_core_129;
  wire popcount25_ikmp_core_130;
  wire popcount25_ikmp_core_131;
  wire popcount25_ikmp_core_132;
  wire popcount25_ikmp_core_133;
  wire popcount25_ikmp_core_135;
  wire popcount25_ikmp_core_137;
  wire popcount25_ikmp_core_138;
  wire popcount25_ikmp_core_140_not;
  wire popcount25_ikmp_core_141;
  wire popcount25_ikmp_core_143;
  wire popcount25_ikmp_core_144;
  wire popcount25_ikmp_core_146;
  wire popcount25_ikmp_core_149;
  wire popcount25_ikmp_core_150;
  wire popcount25_ikmp_core_151;
  wire popcount25_ikmp_core_153;
  wire popcount25_ikmp_core_155;
  wire popcount25_ikmp_core_156;
  wire popcount25_ikmp_core_157;
  wire popcount25_ikmp_core_158;
  wire popcount25_ikmp_core_161;
  wire popcount25_ikmp_core_162_not;
  wire popcount25_ikmp_core_163;
  wire popcount25_ikmp_core_165;
  wire popcount25_ikmp_core_167;
  wire popcount25_ikmp_core_169_not;
  wire popcount25_ikmp_core_171;
  wire popcount25_ikmp_core_173;
  wire popcount25_ikmp_core_174;
  wire popcount25_ikmp_core_175;
  wire popcount25_ikmp_core_176;
  wire popcount25_ikmp_core_178;
  wire popcount25_ikmp_core_179;
  wire popcount25_ikmp_core_180;
  wire popcount25_ikmp_core_182;

  assign popcount25_ikmp_core_027 = input_a[8] ^ input_a[15];
  assign popcount25_ikmp_core_028 = input_a[14] ^ input_a[6];
  assign popcount25_ikmp_core_030 = ~(input_a[12] & input_a[9]);
  assign popcount25_ikmp_core_032 = ~(input_a[19] ^ input_a[7]);
  assign popcount25_ikmp_core_033 = input_a[3] & input_a[21];
  assign popcount25_ikmp_core_036 = ~(input_a[15] ^ input_a[6]);
  assign popcount25_ikmp_core_037 = ~(input_a[11] ^ input_a[9]);
  assign popcount25_ikmp_core_038 = ~(input_a[12] & input_a[15]);
  assign popcount25_ikmp_core_039 = ~(input_a[18] ^ input_a[14]);
  assign popcount25_ikmp_core_040_not = ~input_a[9];
  assign popcount25_ikmp_core_044 = input_a[23] ^ input_a[12];
  assign popcount25_ikmp_core_046 = input_a[4] & input_a[10];
  assign popcount25_ikmp_core_048 = input_a[19] ^ input_a[3];
  assign popcount25_ikmp_core_049 = ~(input_a[1] ^ input_a[7]);
  assign popcount25_ikmp_core_052 = ~input_a[23];
  assign popcount25_ikmp_core_053 = input_a[20] | input_a[4];
  assign popcount25_ikmp_core_056 = ~(input_a[1] ^ input_a[3]);
  assign popcount25_ikmp_core_057 = input_a[6] | input_a[5];
  assign popcount25_ikmp_core_058_not = ~input_a[23];
  assign popcount25_ikmp_core_059 = input_a[9] | input_a[22];
  assign popcount25_ikmp_core_061 = input_a[21] | input_a[15];
  assign popcount25_ikmp_core_062 = ~(input_a[1] ^ input_a[12]);
  assign popcount25_ikmp_core_064 = ~(input_a[6] & input_a[23]);
  assign popcount25_ikmp_core_066 = ~(input_a[16] ^ input_a[13]);
  assign popcount25_ikmp_core_067 = input_a[10] ^ input_a[3];
  assign popcount25_ikmp_core_068 = ~(input_a[15] & input_a[22]);
  assign popcount25_ikmp_core_070 = ~input_a[8];
  assign popcount25_ikmp_core_071 = input_a[0] & input_a[21];
  assign popcount25_ikmp_core_072 = input_a[21] | input_a[23];
  assign popcount25_ikmp_core_073 = ~(input_a[8] & input_a[7]);
  assign popcount25_ikmp_core_075 = ~(input_a[2] | input_a[0]);
  assign popcount25_ikmp_core_076 = input_a[6] | input_a[11];
  assign popcount25_ikmp_core_077 = ~input_a[4];
  assign popcount25_ikmp_core_078 = input_a[12] ^ input_a[22];
  assign popcount25_ikmp_core_079 = ~(input_a[7] & input_a[12]);
  assign popcount25_ikmp_core_080 = ~(input_a[21] ^ input_a[14]);
  assign popcount25_ikmp_core_082 = input_a[12] | input_a[2];
  assign popcount25_ikmp_core_083_not = ~input_a[16];
  assign popcount25_ikmp_core_089 = ~input_a[0];
  assign popcount25_ikmp_core_093 = ~(input_a[1] & input_a[15]);
  assign popcount25_ikmp_core_094 = ~(input_a[2] ^ input_a[5]);
  assign popcount25_ikmp_core_095 = input_a[21] ^ input_a[2];
  assign popcount25_ikmp_core_096 = ~input_a[20];
  assign popcount25_ikmp_core_097 = ~(input_a[22] ^ input_a[8]);
  assign popcount25_ikmp_core_098 = ~(input_a[15] & input_a[8]);
  assign popcount25_ikmp_core_099_not = ~input_a[14];
  assign popcount25_ikmp_core_100 = input_a[12] ^ input_a[9];
  assign popcount25_ikmp_core_102 = ~input_a[0];
  assign popcount25_ikmp_core_105 = input_a[5] & input_a[21];
  assign popcount25_ikmp_core_108 = input_a[11] | input_a[14];
  assign popcount25_ikmp_core_111 = input_a[12] ^ input_a[13];
  assign popcount25_ikmp_core_114 = ~(input_a[1] & input_a[22]);
  assign popcount25_ikmp_core_117 = input_a[13] | input_a[22];
  assign popcount25_ikmp_core_118 = input_a[1] ^ input_a[18];
  assign popcount25_ikmp_core_119 = ~(input_a[23] & input_a[12]);
  assign popcount25_ikmp_core_121 = ~input_a[16];
  assign popcount25_ikmp_core_123 = ~(input_a[8] ^ input_a[8]);
  assign popcount25_ikmp_core_126 = ~(input_a[16] & input_a[12]);
  assign popcount25_ikmp_core_127 = ~input_a[15];
  assign popcount25_ikmp_core_129 = input_a[16] ^ input_a[20];
  assign popcount25_ikmp_core_130 = ~input_a[3];
  assign popcount25_ikmp_core_131 = ~(input_a[13] & input_a[11]);
  assign popcount25_ikmp_core_132 = input_a[17] ^ input_a[2];
  assign popcount25_ikmp_core_133 = input_a[12] ^ input_a[22];
  assign popcount25_ikmp_core_135 = input_a[10] | input_a[0];
  assign popcount25_ikmp_core_137 = ~input_a[20];
  assign popcount25_ikmp_core_138 = ~(input_a[16] & input_a[11]);
  assign popcount25_ikmp_core_140_not = ~input_a[2];
  assign popcount25_ikmp_core_141 = ~input_a[12];
  assign popcount25_ikmp_core_143 = input_a[11] | input_a[24];
  assign popcount25_ikmp_core_144 = ~(input_a[20] | input_a[8]);
  assign popcount25_ikmp_core_146 = ~input_a[1];
  assign popcount25_ikmp_core_149 = ~(input_a[2] ^ input_a[12]);
  assign popcount25_ikmp_core_150 = input_a[23] ^ input_a[13];
  assign popcount25_ikmp_core_151 = ~(input_a[23] | input_a[10]);
  assign popcount25_ikmp_core_153 = ~(input_a[15] | input_a[15]);
  assign popcount25_ikmp_core_155 = input_a[9] | input_a[4];
  assign popcount25_ikmp_core_156 = ~input_a[21];
  assign popcount25_ikmp_core_157 = ~input_a[17];
  assign popcount25_ikmp_core_158 = ~(input_a[7] ^ input_a[0]);
  assign popcount25_ikmp_core_161 = input_a[24] ^ input_a[8];
  assign popcount25_ikmp_core_162_not = ~input_a[15];
  assign popcount25_ikmp_core_163 = ~(input_a[5] ^ input_a[16]);
  assign popcount25_ikmp_core_165 = ~(input_a[15] | input_a[11]);
  assign popcount25_ikmp_core_167 = ~(input_a[11] | input_a[12]);
  assign popcount25_ikmp_core_169_not = ~input_a[7];
  assign popcount25_ikmp_core_171 = input_a[0] | input_a[7];
  assign popcount25_ikmp_core_173 = input_a[18] ^ input_a[20];
  assign popcount25_ikmp_core_174 = input_a[21] ^ input_a[22];
  assign popcount25_ikmp_core_175 = input_a[3] ^ input_a[5];
  assign popcount25_ikmp_core_176 = ~(input_a[9] ^ input_a[16]);
  assign popcount25_ikmp_core_178 = input_a[23] ^ input_a[4];
  assign popcount25_ikmp_core_179 = input_a[12] & input_a[1];
  assign popcount25_ikmp_core_180 = input_a[13] ^ input_a[6];
  assign popcount25_ikmp_core_182 = ~(input_a[0] ^ input_a[21]);

  assign popcount25_ikmp_out[0] = 1'b0;
  assign popcount25_ikmp_out[1] = 1'b0;
  assign popcount25_ikmp_out[2] = 1'b1;
  assign popcount25_ikmp_out[3] = 1'b1;
  assign popcount25_ikmp_out[4] = 1'b0;
endmodule