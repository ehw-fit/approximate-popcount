// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.9187
// WCE=46.0
// EP=0.945984%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_2pl6(input [34:0] input_a, output [5:0] popcount35_2pl6_out);
  wire popcount35_2pl6_core_037_not;
  wire popcount35_2pl6_core_038;
  wire popcount35_2pl6_core_041;
  wire popcount35_2pl6_core_042;
  wire popcount35_2pl6_core_044;
  wire popcount35_2pl6_core_045;
  wire popcount35_2pl6_core_047;
  wire popcount35_2pl6_core_048;
  wire popcount35_2pl6_core_050;
  wire popcount35_2pl6_core_051;
  wire popcount35_2pl6_core_052;
  wire popcount35_2pl6_core_053_not;
  wire popcount35_2pl6_core_056;
  wire popcount35_2pl6_core_058;
  wire popcount35_2pl6_core_060;
  wire popcount35_2pl6_core_063;
  wire popcount35_2pl6_core_065;
  wire popcount35_2pl6_core_066;
  wire popcount35_2pl6_core_067;
  wire popcount35_2pl6_core_068;
  wire popcount35_2pl6_core_069;
  wire popcount35_2pl6_core_070;
  wire popcount35_2pl6_core_071;
  wire popcount35_2pl6_core_072;
  wire popcount35_2pl6_core_073;
  wire popcount35_2pl6_core_074;
  wire popcount35_2pl6_core_075;
  wire popcount35_2pl6_core_077;
  wire popcount35_2pl6_core_078;
  wire popcount35_2pl6_core_082;
  wire popcount35_2pl6_core_083;
  wire popcount35_2pl6_core_086;
  wire popcount35_2pl6_core_087;
  wire popcount35_2pl6_core_088;
  wire popcount35_2pl6_core_089;
  wire popcount35_2pl6_core_090;
  wire popcount35_2pl6_core_091;
  wire popcount35_2pl6_core_094;
  wire popcount35_2pl6_core_097;
  wire popcount35_2pl6_core_100;
  wire popcount35_2pl6_core_101;
  wire popcount35_2pl6_core_103;
  wire popcount35_2pl6_core_105;
  wire popcount35_2pl6_core_107;
  wire popcount35_2pl6_core_108;
  wire popcount35_2pl6_core_110;
  wire popcount35_2pl6_core_111;
  wire popcount35_2pl6_core_112;
  wire popcount35_2pl6_core_113;
  wire popcount35_2pl6_core_114;
  wire popcount35_2pl6_core_115;
  wire popcount35_2pl6_core_116;
  wire popcount35_2pl6_core_117;
  wire popcount35_2pl6_core_119;
  wire popcount35_2pl6_core_123;
  wire popcount35_2pl6_core_126;
  wire popcount35_2pl6_core_127;
  wire popcount35_2pl6_core_128;
  wire popcount35_2pl6_core_129;
  wire popcount35_2pl6_core_130;
  wire popcount35_2pl6_core_131;
  wire popcount35_2pl6_core_134;
  wire popcount35_2pl6_core_135;
  wire popcount35_2pl6_core_136;
  wire popcount35_2pl6_core_137;
  wire popcount35_2pl6_core_138;
  wire popcount35_2pl6_core_139;
  wire popcount35_2pl6_core_142;
  wire popcount35_2pl6_core_144;
  wire popcount35_2pl6_core_146;
  wire popcount35_2pl6_core_147;
  wire popcount35_2pl6_core_150;
  wire popcount35_2pl6_core_152;
  wire popcount35_2pl6_core_153;
  wire popcount35_2pl6_core_155_not;
  wire popcount35_2pl6_core_156;
  wire popcount35_2pl6_core_159;
  wire popcount35_2pl6_core_160;
  wire popcount35_2pl6_core_161;
  wire popcount35_2pl6_core_162;
  wire popcount35_2pl6_core_165;
  wire popcount35_2pl6_core_166;
  wire popcount35_2pl6_core_169;
  wire popcount35_2pl6_core_171;
  wire popcount35_2pl6_core_174;
  wire popcount35_2pl6_core_175;
  wire popcount35_2pl6_core_178;
  wire popcount35_2pl6_core_179;
  wire popcount35_2pl6_core_180;
  wire popcount35_2pl6_core_182;
  wire popcount35_2pl6_core_185;
  wire popcount35_2pl6_core_187;
  wire popcount35_2pl6_core_188;
  wire popcount35_2pl6_core_190;
  wire popcount35_2pl6_core_191;
  wire popcount35_2pl6_core_192;
  wire popcount35_2pl6_core_194;
  wire popcount35_2pl6_core_195;
  wire popcount35_2pl6_core_196;
  wire popcount35_2pl6_core_197;
  wire popcount35_2pl6_core_198;
  wire popcount35_2pl6_core_199;
  wire popcount35_2pl6_core_201;
  wire popcount35_2pl6_core_202;
  wire popcount35_2pl6_core_203;
  wire popcount35_2pl6_core_204;
  wire popcount35_2pl6_core_207;
  wire popcount35_2pl6_core_208;
  wire popcount35_2pl6_core_209;
  wire popcount35_2pl6_core_212;
  wire popcount35_2pl6_core_213;
  wire popcount35_2pl6_core_214;
  wire popcount35_2pl6_core_218;
  wire popcount35_2pl6_core_219;
  wire popcount35_2pl6_core_220;
  wire popcount35_2pl6_core_221;
  wire popcount35_2pl6_core_225;
  wire popcount35_2pl6_core_226;
  wire popcount35_2pl6_core_227;
  wire popcount35_2pl6_core_229;
  wire popcount35_2pl6_core_230;
  wire popcount35_2pl6_core_231;
  wire popcount35_2pl6_core_233;
  wire popcount35_2pl6_core_234;
  wire popcount35_2pl6_core_235;
  wire popcount35_2pl6_core_238;
  wire popcount35_2pl6_core_244_not;
  wire popcount35_2pl6_core_248;
  wire popcount35_2pl6_core_249;
  wire popcount35_2pl6_core_250;
  wire popcount35_2pl6_core_251;
  wire popcount35_2pl6_core_252;
  wire popcount35_2pl6_core_253;
  wire popcount35_2pl6_core_254;
  wire popcount35_2pl6_core_255;
  wire popcount35_2pl6_core_256;
  wire popcount35_2pl6_core_257_not;
  wire popcount35_2pl6_core_260;
  wire popcount35_2pl6_core_262;

  assign popcount35_2pl6_core_037_not = ~input_a[20];
  assign popcount35_2pl6_core_038 = ~(input_a[16] & input_a[17]);
  assign popcount35_2pl6_core_041 = ~(input_a[0] & input_a[4]);
  assign popcount35_2pl6_core_042 = ~input_a[26];
  assign popcount35_2pl6_core_044 = input_a[34] | input_a[27];
  assign popcount35_2pl6_core_045 = ~(input_a[32] & input_a[13]);
  assign popcount35_2pl6_core_047 = ~(input_a[29] | input_a[5]);
  assign popcount35_2pl6_core_048 = ~(input_a[26] | input_a[25]);
  assign popcount35_2pl6_core_050 = input_a[25] | input_a[27];
  assign popcount35_2pl6_core_051 = ~(input_a[7] & input_a[34]);
  assign popcount35_2pl6_core_052 = ~(input_a[5] ^ input_a[31]);
  assign popcount35_2pl6_core_053_not = ~input_a[2];
  assign popcount35_2pl6_core_056 = input_a[23] ^ input_a[27];
  assign popcount35_2pl6_core_058 = ~(input_a[22] ^ input_a[12]);
  assign popcount35_2pl6_core_060 = ~(input_a[31] | input_a[20]);
  assign popcount35_2pl6_core_063 = ~(input_a[11] ^ input_a[6]);
  assign popcount35_2pl6_core_065 = input_a[28] & input_a[22];
  assign popcount35_2pl6_core_066 = ~(input_a[20] ^ input_a[10]);
  assign popcount35_2pl6_core_067 = input_a[30] & input_a[24];
  assign popcount35_2pl6_core_068 = input_a[3] & input_a[13];
  assign popcount35_2pl6_core_069 = input_a[15] & input_a[31];
  assign popcount35_2pl6_core_070 = ~(input_a[1] & input_a[1]);
  assign popcount35_2pl6_core_071 = ~(input_a[4] & input_a[34]);
  assign popcount35_2pl6_core_072 = ~(input_a[12] | input_a[26]);
  assign popcount35_2pl6_core_073 = input_a[16] ^ input_a[27];
  assign popcount35_2pl6_core_074 = ~(input_a[2] ^ input_a[27]);
  assign popcount35_2pl6_core_075 = input_a[29] ^ input_a[9];
  assign popcount35_2pl6_core_077 = input_a[32] & input_a[27];
  assign popcount35_2pl6_core_078 = ~(input_a[13] ^ input_a[32]);
  assign popcount35_2pl6_core_082 = ~(input_a[25] & input_a[13]);
  assign popcount35_2pl6_core_083 = input_a[9] & input_a[6];
  assign popcount35_2pl6_core_086 = input_a[22] & input_a[5];
  assign popcount35_2pl6_core_087 = ~(input_a[14] | input_a[10]);
  assign popcount35_2pl6_core_088 = ~(input_a[9] | input_a[7]);
  assign popcount35_2pl6_core_089 = ~(input_a[20] | input_a[4]);
  assign popcount35_2pl6_core_090 = ~input_a[34];
  assign popcount35_2pl6_core_091 = input_a[20] ^ input_a[32];
  assign popcount35_2pl6_core_094 = ~input_a[12];
  assign popcount35_2pl6_core_097 = input_a[14] ^ input_a[3];
  assign popcount35_2pl6_core_100 = ~(input_a[7] & input_a[19]);
  assign popcount35_2pl6_core_101 = ~input_a[18];
  assign popcount35_2pl6_core_103 = input_a[16] | input_a[4];
  assign popcount35_2pl6_core_105 = ~input_a[6];
  assign popcount35_2pl6_core_107 = input_a[13] & input_a[20];
  assign popcount35_2pl6_core_108 = ~input_a[27];
  assign popcount35_2pl6_core_110 = ~input_a[29];
  assign popcount35_2pl6_core_111 = input_a[32] ^ input_a[34];
  assign popcount35_2pl6_core_112 = ~(input_a[17] | input_a[8]);
  assign popcount35_2pl6_core_113 = input_a[26] & input_a[7];
  assign popcount35_2pl6_core_114 = ~input_a[11];
  assign popcount35_2pl6_core_115 = ~(input_a[10] & input_a[24]);
  assign popcount35_2pl6_core_116 = input_a[11] & input_a[4];
  assign popcount35_2pl6_core_117 = ~(input_a[2] ^ input_a[26]);
  assign popcount35_2pl6_core_119 = ~input_a[22];
  assign popcount35_2pl6_core_123 = input_a[31] | input_a[23];
  assign popcount35_2pl6_core_126 = ~(input_a[4] | input_a[5]);
  assign popcount35_2pl6_core_127 = input_a[1] | input_a[29];
  assign popcount35_2pl6_core_128 = ~(input_a[21] & input_a[31]);
  assign popcount35_2pl6_core_129 = input_a[14] ^ input_a[23];
  assign popcount35_2pl6_core_130 = input_a[18] & input_a[23];
  assign popcount35_2pl6_core_131 = ~(input_a[7] & input_a[5]);
  assign popcount35_2pl6_core_134 = ~(input_a[14] & input_a[27]);
  assign popcount35_2pl6_core_135 = ~input_a[5];
  assign popcount35_2pl6_core_136 = ~(input_a[26] | input_a[1]);
  assign popcount35_2pl6_core_137 = ~(input_a[30] ^ input_a[26]);
  assign popcount35_2pl6_core_138 = input_a[21] & input_a[7];
  assign popcount35_2pl6_core_139 = ~(input_a[10] & input_a[31]);
  assign popcount35_2pl6_core_142 = ~(input_a[12] & input_a[32]);
  assign popcount35_2pl6_core_144 = input_a[21] | input_a[30];
  assign popcount35_2pl6_core_146 = ~(input_a[31] & input_a[17]);
  assign popcount35_2pl6_core_147 = ~(input_a[4] ^ input_a[0]);
  assign popcount35_2pl6_core_150 = ~(input_a[0] ^ input_a[28]);
  assign popcount35_2pl6_core_152 = ~(input_a[4] & input_a[14]);
  assign popcount35_2pl6_core_153 = input_a[11] ^ input_a[7];
  assign popcount35_2pl6_core_155_not = ~input_a[7];
  assign popcount35_2pl6_core_156 = input_a[8] | input_a[20];
  assign popcount35_2pl6_core_159 = ~input_a[32];
  assign popcount35_2pl6_core_160 = input_a[3] ^ input_a[4];
  assign popcount35_2pl6_core_161 = ~(input_a[0] | input_a[6]);
  assign popcount35_2pl6_core_162 = ~(input_a[11] & input_a[10]);
  assign popcount35_2pl6_core_165 = ~input_a[12];
  assign popcount35_2pl6_core_166 = input_a[28] ^ input_a[26];
  assign popcount35_2pl6_core_169 = ~(input_a[23] & input_a[13]);
  assign popcount35_2pl6_core_171 = input_a[26] | input_a[20];
  assign popcount35_2pl6_core_174 = ~(input_a[12] | input_a[20]);
  assign popcount35_2pl6_core_175 = ~(input_a[1] ^ input_a[28]);
  assign popcount35_2pl6_core_178 = ~(input_a[18] & input_a[28]);
  assign popcount35_2pl6_core_179 = ~(input_a[30] ^ input_a[27]);
  assign popcount35_2pl6_core_180 = input_a[25] | input_a[8];
  assign popcount35_2pl6_core_182 = input_a[27] ^ input_a[29];
  assign popcount35_2pl6_core_185 = ~input_a[11];
  assign popcount35_2pl6_core_187 = ~(input_a[28] & input_a[5]);
  assign popcount35_2pl6_core_188 = input_a[16] ^ input_a[23];
  assign popcount35_2pl6_core_190 = input_a[16] ^ input_a[12];
  assign popcount35_2pl6_core_191 = input_a[13] ^ input_a[8];
  assign popcount35_2pl6_core_192 = ~input_a[15];
  assign popcount35_2pl6_core_194 = ~input_a[5];
  assign popcount35_2pl6_core_195 = input_a[13] | input_a[33];
  assign popcount35_2pl6_core_196 = input_a[1] ^ input_a[6];
  assign popcount35_2pl6_core_197 = input_a[29] | input_a[5];
  assign popcount35_2pl6_core_198 = ~(input_a[14] ^ input_a[22]);
  assign popcount35_2pl6_core_199 = input_a[25] & input_a[17];
  assign popcount35_2pl6_core_201 = ~(input_a[11] | input_a[23]);
  assign popcount35_2pl6_core_202 = input_a[12] | input_a[16];
  assign popcount35_2pl6_core_203 = input_a[3] ^ input_a[16];
  assign popcount35_2pl6_core_204 = input_a[15] | input_a[22];
  assign popcount35_2pl6_core_207 = input_a[16] ^ input_a[12];
  assign popcount35_2pl6_core_208 = ~input_a[10];
  assign popcount35_2pl6_core_209 = input_a[25] | input_a[30];
  assign popcount35_2pl6_core_212 = ~(input_a[9] & input_a[2]);
  assign popcount35_2pl6_core_213 = input_a[17] | input_a[30];
  assign popcount35_2pl6_core_214 = input_a[20] | input_a[11];
  assign popcount35_2pl6_core_218 = input_a[18] | input_a[11];
  assign popcount35_2pl6_core_219 = input_a[31] & input_a[30];
  assign popcount35_2pl6_core_220 = ~(input_a[23] & input_a[13]);
  assign popcount35_2pl6_core_221 = input_a[8] | input_a[19];
  assign popcount35_2pl6_core_225 = input_a[11] & input_a[28];
  assign popcount35_2pl6_core_226 = ~(input_a[6] & input_a[27]);
  assign popcount35_2pl6_core_227 = input_a[6] | input_a[22];
  assign popcount35_2pl6_core_229 = input_a[33] | input_a[6];
  assign popcount35_2pl6_core_230 = ~input_a[34];
  assign popcount35_2pl6_core_231 = ~(input_a[4] | input_a[13]);
  assign popcount35_2pl6_core_233 = ~(input_a[34] | input_a[12]);
  assign popcount35_2pl6_core_234 = input_a[34] ^ input_a[10];
  assign popcount35_2pl6_core_235 = ~(input_a[26] | input_a[30]);
  assign popcount35_2pl6_core_238 = input_a[27] | input_a[17];
  assign popcount35_2pl6_core_244_not = ~input_a[30];
  assign popcount35_2pl6_core_248 = input_a[7] ^ input_a[11];
  assign popcount35_2pl6_core_249 = input_a[21] & input_a[7];
  assign popcount35_2pl6_core_250 = input_a[11] & input_a[29];
  assign popcount35_2pl6_core_251 = input_a[28] & input_a[0];
  assign popcount35_2pl6_core_252 = input_a[19] & input_a[9];
  assign popcount35_2pl6_core_253 = ~(input_a[3] ^ input_a[7]);
  assign popcount35_2pl6_core_254 = ~input_a[12];
  assign popcount35_2pl6_core_255 = input_a[2] ^ input_a[14];
  assign popcount35_2pl6_core_256 = ~(input_a[17] | input_a[2]);
  assign popcount35_2pl6_core_257_not = ~input_a[16];
  assign popcount35_2pl6_core_260 = input_a[8] & input_a[5];
  assign popcount35_2pl6_core_262 = ~(input_a[26] ^ input_a[31]);

  assign popcount35_2pl6_out[0] = 1'b1;
  assign popcount35_2pl6_out[1] = 1'b1;
  assign popcount35_2pl6_out[2] = 1'b1;
  assign popcount35_2pl6_out[3] = 1'b1;
  assign popcount35_2pl6_out[4] = 1'b0;
  assign popcount35_2pl6_out[5] = input_a[7];
endmodule