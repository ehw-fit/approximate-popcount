// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.52363
// WCE=27.0
// EP=0.990208%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_bt0q(input [37:0] input_a, output [5:0] popcount38_bt0q_out);
  wire popcount38_bt0q_core_040;
  wire popcount38_bt0q_core_041;
  wire popcount38_bt0q_core_042;
  wire popcount38_bt0q_core_044;
  wire popcount38_bt0q_core_046;
  wire popcount38_bt0q_core_047;
  wire popcount38_bt0q_core_048;
  wire popcount38_bt0q_core_051;
  wire popcount38_bt0q_core_052;
  wire popcount38_bt0q_core_054;
  wire popcount38_bt0q_core_055;
  wire popcount38_bt0q_core_056;
  wire popcount38_bt0q_core_058;
  wire popcount38_bt0q_core_060;
  wire popcount38_bt0q_core_062;
  wire popcount38_bt0q_core_063_not;
  wire popcount38_bt0q_core_064;
  wire popcount38_bt0q_core_065;
  wire popcount38_bt0q_core_067;
  wire popcount38_bt0q_core_068;
  wire popcount38_bt0q_core_069;
  wire popcount38_bt0q_core_070;
  wire popcount38_bt0q_core_071;
  wire popcount38_bt0q_core_072;
  wire popcount38_bt0q_core_073;
  wire popcount38_bt0q_core_075;
  wire popcount38_bt0q_core_076;
  wire popcount38_bt0q_core_077;
  wire popcount38_bt0q_core_080;
  wire popcount38_bt0q_core_081;
  wire popcount38_bt0q_core_084;
  wire popcount38_bt0q_core_087;
  wire popcount38_bt0q_core_088;
  wire popcount38_bt0q_core_090;
  wire popcount38_bt0q_core_091;
  wire popcount38_bt0q_core_092;
  wire popcount38_bt0q_core_095;
  wire popcount38_bt0q_core_097;
  wire popcount38_bt0q_core_099;
  wire popcount38_bt0q_core_102;
  wire popcount38_bt0q_core_103;
  wire popcount38_bt0q_core_104;
  wire popcount38_bt0q_core_108;
  wire popcount38_bt0q_core_109;
  wire popcount38_bt0q_core_110;
  wire popcount38_bt0q_core_111;
  wire popcount38_bt0q_core_112_not;
  wire popcount38_bt0q_core_113;
  wire popcount38_bt0q_core_114;
  wire popcount38_bt0q_core_115;
  wire popcount38_bt0q_core_118;
  wire popcount38_bt0q_core_119;
  wire popcount38_bt0q_core_120;
  wire popcount38_bt0q_core_121;
  wire popcount38_bt0q_core_122;
  wire popcount38_bt0q_core_123;
  wire popcount38_bt0q_core_125;
  wire popcount38_bt0q_core_126;
  wire popcount38_bt0q_core_128;
  wire popcount38_bt0q_core_129;
  wire popcount38_bt0q_core_130;
  wire popcount38_bt0q_core_131;
  wire popcount38_bt0q_core_133;
  wire popcount38_bt0q_core_134;
  wire popcount38_bt0q_core_136;
  wire popcount38_bt0q_core_142;
  wire popcount38_bt0q_core_143;
  wire popcount38_bt0q_core_145;
  wire popcount38_bt0q_core_146;
  wire popcount38_bt0q_core_147;
  wire popcount38_bt0q_core_148;
  wire popcount38_bt0q_core_150;
  wire popcount38_bt0q_core_151;
  wire popcount38_bt0q_core_152;
  wire popcount38_bt0q_core_153_not;
  wire popcount38_bt0q_core_154;
  wire popcount38_bt0q_core_156;
  wire popcount38_bt0q_core_160;
  wire popcount38_bt0q_core_161;
  wire popcount38_bt0q_core_163;
  wire popcount38_bt0q_core_165;
  wire popcount38_bt0q_core_166;
  wire popcount38_bt0q_core_167;
  wire popcount38_bt0q_core_168;
  wire popcount38_bt0q_core_169;
  wire popcount38_bt0q_core_171;
  wire popcount38_bt0q_core_172;
  wire popcount38_bt0q_core_174;
  wire popcount38_bt0q_core_176;
  wire popcount38_bt0q_core_177;
  wire popcount38_bt0q_core_179;
  wire popcount38_bt0q_core_181;
  wire popcount38_bt0q_core_183;
  wire popcount38_bt0q_core_184;
  wire popcount38_bt0q_core_185;
  wire popcount38_bt0q_core_186;
  wire popcount38_bt0q_core_188;
  wire popcount38_bt0q_core_189;
  wire popcount38_bt0q_core_190;
  wire popcount38_bt0q_core_193;
  wire popcount38_bt0q_core_195;
  wire popcount38_bt0q_core_196;
  wire popcount38_bt0q_core_198;
  wire popcount38_bt0q_core_199;
  wire popcount38_bt0q_core_200;
  wire popcount38_bt0q_core_201;
  wire popcount38_bt0q_core_202;
  wire popcount38_bt0q_core_203;
  wire popcount38_bt0q_core_204;
  wire popcount38_bt0q_core_205;
  wire popcount38_bt0q_core_206;
  wire popcount38_bt0q_core_208;
  wire popcount38_bt0q_core_210;
  wire popcount38_bt0q_core_213;
  wire popcount38_bt0q_core_214;
  wire popcount38_bt0q_core_216;
  wire popcount38_bt0q_core_218;
  wire popcount38_bt0q_core_219;
  wire popcount38_bt0q_core_221;
  wire popcount38_bt0q_core_222;
  wire popcount38_bt0q_core_225;
  wire popcount38_bt0q_core_226;
  wire popcount38_bt0q_core_227;
  wire popcount38_bt0q_core_228;
  wire popcount38_bt0q_core_229;
  wire popcount38_bt0q_core_230;
  wire popcount38_bt0q_core_231;
  wire popcount38_bt0q_core_233;
  wire popcount38_bt0q_core_234_not;
  wire popcount38_bt0q_core_237_not;
  wire popcount38_bt0q_core_239;
  wire popcount38_bt0q_core_244;
  wire popcount38_bt0q_core_246_not;
  wire popcount38_bt0q_core_247;
  wire popcount38_bt0q_core_250;
  wire popcount38_bt0q_core_251;
  wire popcount38_bt0q_core_252;
  wire popcount38_bt0q_core_253;
  wire popcount38_bt0q_core_254;
  wire popcount38_bt0q_core_256;
  wire popcount38_bt0q_core_257;
  wire popcount38_bt0q_core_258;
  wire popcount38_bt0q_core_259;
  wire popcount38_bt0q_core_260;
  wire popcount38_bt0q_core_262;
  wire popcount38_bt0q_core_264;
  wire popcount38_bt0q_core_267;
  wire popcount38_bt0q_core_268;
  wire popcount38_bt0q_core_270;
  wire popcount38_bt0q_core_272;
  wire popcount38_bt0q_core_273;
  wire popcount38_bt0q_core_274;
  wire popcount38_bt0q_core_275;
  wire popcount38_bt0q_core_276;
  wire popcount38_bt0q_core_277;
  wire popcount38_bt0q_core_279;
  wire popcount38_bt0q_core_280;
  wire popcount38_bt0q_core_282;
  wire popcount38_bt0q_core_284;
  wire popcount38_bt0q_core_285;
  wire popcount38_bt0q_core_287;
  wire popcount38_bt0q_core_288;
  wire popcount38_bt0q_core_291;
  wire popcount38_bt0q_core_292;
  wire popcount38_bt0q_core_293;
  wire popcount38_bt0q_core_296;

  assign popcount38_bt0q_core_040 = input_a[11] & input_a[10];
  assign popcount38_bt0q_core_041 = ~(input_a[3] ^ input_a[34]);
  assign popcount38_bt0q_core_042 = ~(input_a[27] ^ input_a[33]);
  assign popcount38_bt0q_core_044 = ~(input_a[9] & input_a[12]);
  assign popcount38_bt0q_core_046 = input_a[36] ^ input_a[16];
  assign popcount38_bt0q_core_047 = input_a[14] ^ input_a[19];
  assign popcount38_bt0q_core_048 = ~(input_a[35] & input_a[13]);
  assign popcount38_bt0q_core_051 = input_a[7] & input_a[11];
  assign popcount38_bt0q_core_052 = ~(input_a[11] ^ input_a[16]);
  assign popcount38_bt0q_core_054 = ~(input_a[31] ^ input_a[5]);
  assign popcount38_bt0q_core_055 = input_a[21] | input_a[22];
  assign popcount38_bt0q_core_056 = ~input_a[10];
  assign popcount38_bt0q_core_058 = input_a[8] | input_a[2];
  assign popcount38_bt0q_core_060 = input_a[5] & input_a[4];
  assign popcount38_bt0q_core_062 = input_a[34] & input_a[1];
  assign popcount38_bt0q_core_063_not = ~input_a[21];
  assign popcount38_bt0q_core_064 = input_a[2] & input_a[10];
  assign popcount38_bt0q_core_065 = ~(input_a[13] & input_a[24]);
  assign popcount38_bt0q_core_067 = ~(input_a[37] | input_a[30]);
  assign popcount38_bt0q_core_068 = input_a[33] ^ input_a[9];
  assign popcount38_bt0q_core_069 = ~input_a[0];
  assign popcount38_bt0q_core_070 = input_a[11] & input_a[27];
  assign popcount38_bt0q_core_071 = input_a[20] ^ input_a[28];
  assign popcount38_bt0q_core_072 = ~(input_a[0] ^ input_a[27]);
  assign popcount38_bt0q_core_073 = ~(input_a[28] ^ input_a[34]);
  assign popcount38_bt0q_core_075 = ~(input_a[37] & input_a[21]);
  assign popcount38_bt0q_core_076 = input_a[8] | input_a[29];
  assign popcount38_bt0q_core_077 = ~input_a[20];
  assign popcount38_bt0q_core_080 = ~input_a[12];
  assign popcount38_bt0q_core_081 = input_a[33] & input_a[31];
  assign popcount38_bt0q_core_084 = input_a[21] & input_a[1];
  assign popcount38_bt0q_core_087 = input_a[23] & input_a[34];
  assign popcount38_bt0q_core_088 = ~(input_a[22] & input_a[20]);
  assign popcount38_bt0q_core_090 = ~(input_a[17] & input_a[26]);
  assign popcount38_bt0q_core_091 = ~(input_a[35] & input_a[1]);
  assign popcount38_bt0q_core_092 = ~input_a[34];
  assign popcount38_bt0q_core_095 = ~(input_a[34] | input_a[21]);
  assign popcount38_bt0q_core_097 = ~input_a[9];
  assign popcount38_bt0q_core_099 = input_a[15] ^ input_a[34];
  assign popcount38_bt0q_core_102 = input_a[25] & input_a[10];
  assign popcount38_bt0q_core_103 = ~(input_a[9] ^ input_a[26]);
  assign popcount38_bt0q_core_104 = ~(input_a[22] | input_a[31]);
  assign popcount38_bt0q_core_108 = ~(input_a[7] ^ input_a[33]);
  assign popcount38_bt0q_core_109 = ~(input_a[26] ^ input_a[5]);
  assign popcount38_bt0q_core_110 = ~(input_a[15] ^ input_a[7]);
  assign popcount38_bt0q_core_111 = input_a[3] | input_a[13];
  assign popcount38_bt0q_core_112_not = ~input_a[7];
  assign popcount38_bt0q_core_113 = input_a[7] ^ input_a[8];
  assign popcount38_bt0q_core_114 = ~(input_a[27] | input_a[5]);
  assign popcount38_bt0q_core_115 = ~(input_a[9] | input_a[18]);
  assign popcount38_bt0q_core_118 = ~input_a[2];
  assign popcount38_bt0q_core_119 = input_a[29] & input_a[21];
  assign popcount38_bt0q_core_120 = ~(input_a[30] & input_a[35]);
  assign popcount38_bt0q_core_121 = input_a[33] ^ input_a[8];
  assign popcount38_bt0q_core_122 = ~(input_a[18] ^ input_a[34]);
  assign popcount38_bt0q_core_123 = input_a[2] | input_a[33];
  assign popcount38_bt0q_core_125 = ~(input_a[30] & input_a[23]);
  assign popcount38_bt0q_core_126 = ~(input_a[30] ^ input_a[23]);
  assign popcount38_bt0q_core_128 = ~input_a[19];
  assign popcount38_bt0q_core_129 = ~(input_a[27] & input_a[0]);
  assign popcount38_bt0q_core_130 = ~input_a[31];
  assign popcount38_bt0q_core_131 = input_a[5] ^ input_a[22];
  assign popcount38_bt0q_core_133 = ~(input_a[15] | input_a[31]);
  assign popcount38_bt0q_core_134 = input_a[2] | input_a[26];
  assign popcount38_bt0q_core_136 = input_a[7] ^ input_a[1];
  assign popcount38_bt0q_core_142 = ~(input_a[19] | input_a[31]);
  assign popcount38_bt0q_core_143 = input_a[9] ^ input_a[16];
  assign popcount38_bt0q_core_145 = ~(input_a[3] ^ input_a[11]);
  assign popcount38_bt0q_core_146 = input_a[24] | input_a[2];
  assign popcount38_bt0q_core_147 = input_a[29] & input_a[3];
  assign popcount38_bt0q_core_148 = ~(input_a[30] & input_a[30]);
  assign popcount38_bt0q_core_150 = input_a[37] & input_a[14];
  assign popcount38_bt0q_core_151 = ~(input_a[34] & input_a[7]);
  assign popcount38_bt0q_core_152 = ~(input_a[32] & input_a[25]);
  assign popcount38_bt0q_core_153_not = ~input_a[24];
  assign popcount38_bt0q_core_154 = input_a[32] ^ input_a[27];
  assign popcount38_bt0q_core_156 = input_a[34] & input_a[0];
  assign popcount38_bt0q_core_160 = input_a[35] & input_a[28];
  assign popcount38_bt0q_core_161 = input_a[22] & input_a[12];
  assign popcount38_bt0q_core_163 = ~input_a[23];
  assign popcount38_bt0q_core_165 = ~input_a[5];
  assign popcount38_bt0q_core_166 = input_a[34] & input_a[33];
  assign popcount38_bt0q_core_167 = ~(input_a[10] ^ input_a[21]);
  assign popcount38_bt0q_core_168 = input_a[12] ^ input_a[1];
  assign popcount38_bt0q_core_169 = ~input_a[14];
  assign popcount38_bt0q_core_171 = input_a[16] | input_a[1];
  assign popcount38_bt0q_core_172 = ~(input_a[5] ^ input_a[21]);
  assign popcount38_bt0q_core_174 = input_a[15] ^ input_a[3];
  assign popcount38_bt0q_core_176 = input_a[17] | input_a[15];
  assign popcount38_bt0q_core_177 = ~(input_a[29] & input_a[0]);
  assign popcount38_bt0q_core_179 = input_a[3] & input_a[2];
  assign popcount38_bt0q_core_181 = ~(input_a[20] ^ input_a[30]);
  assign popcount38_bt0q_core_183 = ~(input_a[32] & input_a[37]);
  assign popcount38_bt0q_core_184 = ~(input_a[8] ^ input_a[12]);
  assign popcount38_bt0q_core_185 = input_a[6] ^ input_a[33];
  assign popcount38_bt0q_core_186 = input_a[28] ^ input_a[18];
  assign popcount38_bt0q_core_188 = ~(input_a[15] & input_a[0]);
  assign popcount38_bt0q_core_189 = ~(input_a[31] & input_a[13]);
  assign popcount38_bt0q_core_190 = ~(input_a[24] ^ input_a[24]);
  assign popcount38_bt0q_core_193 = ~(input_a[24] ^ input_a[36]);
  assign popcount38_bt0q_core_195 = input_a[19] | input_a[26];
  assign popcount38_bt0q_core_196 = ~(input_a[6] | input_a[19]);
  assign popcount38_bt0q_core_198 = ~(input_a[9] & input_a[32]);
  assign popcount38_bt0q_core_199 = input_a[11] & input_a[30];
  assign popcount38_bt0q_core_200 = input_a[6] | input_a[23];
  assign popcount38_bt0q_core_201 = ~(input_a[11] ^ input_a[7]);
  assign popcount38_bt0q_core_202 = input_a[29] ^ input_a[36];
  assign popcount38_bt0q_core_203 = ~(input_a[26] ^ input_a[17]);
  assign popcount38_bt0q_core_204 = input_a[4] ^ input_a[15];
  assign popcount38_bt0q_core_205 = input_a[26] ^ input_a[33];
  assign popcount38_bt0q_core_206 = input_a[35] & input_a[30];
  assign popcount38_bt0q_core_208 = input_a[3] | input_a[2];
  assign popcount38_bt0q_core_210 = ~(input_a[34] & input_a[19]);
  assign popcount38_bt0q_core_213 = input_a[32] | input_a[9];
  assign popcount38_bt0q_core_214 = input_a[13] ^ input_a[6];
  assign popcount38_bt0q_core_216 = ~(input_a[29] | input_a[28]);
  assign popcount38_bt0q_core_218 = ~(input_a[21] ^ input_a[25]);
  assign popcount38_bt0q_core_219 = ~input_a[14];
  assign popcount38_bt0q_core_221 = ~input_a[28];
  assign popcount38_bt0q_core_222 = ~(input_a[9] | input_a[0]);
  assign popcount38_bt0q_core_225 = ~(input_a[37] | input_a[7]);
  assign popcount38_bt0q_core_226 = input_a[13] ^ input_a[27];
  assign popcount38_bt0q_core_227 = input_a[24] ^ input_a[26];
  assign popcount38_bt0q_core_228 = ~input_a[37];
  assign popcount38_bt0q_core_229 = ~(input_a[11] ^ input_a[37]);
  assign popcount38_bt0q_core_230 = ~(input_a[27] | input_a[18]);
  assign popcount38_bt0q_core_231 = ~input_a[1];
  assign popcount38_bt0q_core_233 = input_a[2] & input_a[3];
  assign popcount38_bt0q_core_234_not = ~input_a[32];
  assign popcount38_bt0q_core_237_not = ~input_a[4];
  assign popcount38_bt0q_core_239 = input_a[17] | input_a[12];
  assign popcount38_bt0q_core_244 = ~(input_a[25] & input_a[20]);
  assign popcount38_bt0q_core_246_not = ~input_a[14];
  assign popcount38_bt0q_core_247 = input_a[18] | input_a[13];
  assign popcount38_bt0q_core_250 = ~input_a[0];
  assign popcount38_bt0q_core_251 = input_a[21] ^ input_a[4];
  assign popcount38_bt0q_core_252 = ~(input_a[5] ^ input_a[13]);
  assign popcount38_bt0q_core_253 = ~input_a[24];
  assign popcount38_bt0q_core_254 = input_a[31] ^ input_a[8];
  assign popcount38_bt0q_core_256 = input_a[17] ^ input_a[14];
  assign popcount38_bt0q_core_257 = input_a[2] | input_a[9];
  assign popcount38_bt0q_core_258 = ~(input_a[10] | input_a[27]);
  assign popcount38_bt0q_core_259 = input_a[31] | input_a[9];
  assign popcount38_bt0q_core_260 = input_a[18] & input_a[17];
  assign popcount38_bt0q_core_262 = input_a[4] & input_a[32];
  assign popcount38_bt0q_core_264 = ~(input_a[21] | input_a[20]);
  assign popcount38_bt0q_core_267 = input_a[18] | input_a[23];
  assign popcount38_bt0q_core_268 = ~(input_a[14] ^ input_a[18]);
  assign popcount38_bt0q_core_270 = ~input_a[11];
  assign popcount38_bt0q_core_272 = ~input_a[15];
  assign popcount38_bt0q_core_273 = input_a[23] | input_a[19];
  assign popcount38_bt0q_core_274 = input_a[12] ^ input_a[21];
  assign popcount38_bt0q_core_275 = ~(input_a[16] | input_a[23]);
  assign popcount38_bt0q_core_276 = ~input_a[0];
  assign popcount38_bt0q_core_277 = ~input_a[18];
  assign popcount38_bt0q_core_279 = ~(input_a[35] & input_a[17]);
  assign popcount38_bt0q_core_280 = ~(input_a[27] | input_a[4]);
  assign popcount38_bt0q_core_282 = input_a[8] ^ input_a[11];
  assign popcount38_bt0q_core_284 = ~(input_a[22] ^ input_a[1]);
  assign popcount38_bt0q_core_285 = input_a[13] & input_a[4];
  assign popcount38_bt0q_core_287 = input_a[9] ^ input_a[37];
  assign popcount38_bt0q_core_288 = input_a[31] ^ input_a[7];
  assign popcount38_bt0q_core_291 = input_a[17] ^ input_a[25];
  assign popcount38_bt0q_core_292 = ~(input_a[6] & input_a[17]);
  assign popcount38_bt0q_core_293 = ~(input_a[21] ^ input_a[13]);
  assign popcount38_bt0q_core_296 = ~(input_a[34] | input_a[21]);

  assign popcount38_bt0q_out[0] = 1'b1;
  assign popcount38_bt0q_out[1] = 1'b0;
  assign popcount38_bt0q_out[2] = input_a[22];
  assign popcount38_bt0q_out[3] = 1'b1;
  assign popcount38_bt0q_out[4] = input_a[36];
  assign popcount38_bt0q_out[5] = 1'b0;
endmodule