// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.69417
// WCE=21.0
// EP=0.953061%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_37rn(input [29:0] input_a, output [4:0] popcount30_37rn_out);
  wire popcount30_37rn_core_032;
  wire popcount30_37rn_core_033;
  wire popcount30_37rn_core_034;
  wire popcount30_37rn_core_035;
  wire popcount30_37rn_core_038;
  wire popcount30_37rn_core_039;
  wire popcount30_37rn_core_040;
  wire popcount30_37rn_core_043;
  wire popcount30_37rn_core_044;
  wire popcount30_37rn_core_046;
  wire popcount30_37rn_core_047;
  wire popcount30_37rn_core_049;
  wire popcount30_37rn_core_051;
  wire popcount30_37rn_core_054;
  wire popcount30_37rn_core_056;
  wire popcount30_37rn_core_057_not;
  wire popcount30_37rn_core_059;
  wire popcount30_37rn_core_062;
  wire popcount30_37rn_core_065;
  wire popcount30_37rn_core_066;
  wire popcount30_37rn_core_067;
  wire popcount30_37rn_core_069;
  wire popcount30_37rn_core_072;
  wire popcount30_37rn_core_074;
  wire popcount30_37rn_core_076;
  wire popcount30_37rn_core_080;
  wire popcount30_37rn_core_082;
  wire popcount30_37rn_core_083;
  wire popcount30_37rn_core_085;
  wire popcount30_37rn_core_086;
  wire popcount30_37rn_core_087;
  wire popcount30_37rn_core_089;
  wire popcount30_37rn_core_092_not;
  wire popcount30_37rn_core_093;
  wire popcount30_37rn_core_094;
  wire popcount30_37rn_core_095;
  wire popcount30_37rn_core_098;
  wire popcount30_37rn_core_099;
  wire popcount30_37rn_core_101;
  wire popcount30_37rn_core_102;
  wire popcount30_37rn_core_107;
  wire popcount30_37rn_core_108;
  wire popcount30_37rn_core_109;
  wire popcount30_37rn_core_111;
  wire popcount30_37rn_core_113;
  wire popcount30_37rn_core_115;
  wire popcount30_37rn_core_116;
  wire popcount30_37rn_core_117;
  wire popcount30_37rn_core_120;
  wire popcount30_37rn_core_121;
  wire popcount30_37rn_core_122;
  wire popcount30_37rn_core_123_not;
  wire popcount30_37rn_core_125;
  wire popcount30_37rn_core_126;
  wire popcount30_37rn_core_127;
  wire popcount30_37rn_core_128;
  wire popcount30_37rn_core_130;
  wire popcount30_37rn_core_131;
  wire popcount30_37rn_core_132;
  wire popcount30_37rn_core_135;
  wire popcount30_37rn_core_137;
  wire popcount30_37rn_core_138;
  wire popcount30_37rn_core_139;
  wire popcount30_37rn_core_141;
  wire popcount30_37rn_core_142;
  wire popcount30_37rn_core_143;
  wire popcount30_37rn_core_144;
  wire popcount30_37rn_core_146;
  wire popcount30_37rn_core_147;
  wire popcount30_37rn_core_149;
  wire popcount30_37rn_core_150_not;
  wire popcount30_37rn_core_152;
  wire popcount30_37rn_core_153;
  wire popcount30_37rn_core_156;
  wire popcount30_37rn_core_157;
  wire popcount30_37rn_core_158;
  wire popcount30_37rn_core_159;
  wire popcount30_37rn_core_160;
  wire popcount30_37rn_core_162;
  wire popcount30_37rn_core_163;
  wire popcount30_37rn_core_164;
  wire popcount30_37rn_core_165;
  wire popcount30_37rn_core_167;
  wire popcount30_37rn_core_168_not;
  wire popcount30_37rn_core_170;
  wire popcount30_37rn_core_171;
  wire popcount30_37rn_core_172;
  wire popcount30_37rn_core_173;
  wire popcount30_37rn_core_175;
  wire popcount30_37rn_core_177;
  wire popcount30_37rn_core_178;
  wire popcount30_37rn_core_179;
  wire popcount30_37rn_core_180;
  wire popcount30_37rn_core_181;
  wire popcount30_37rn_core_182_not;
  wire popcount30_37rn_core_184;
  wire popcount30_37rn_core_185;
  wire popcount30_37rn_core_187;
  wire popcount30_37rn_core_188;
  wire popcount30_37rn_core_189;
  wire popcount30_37rn_core_190;
  wire popcount30_37rn_core_191;
  wire popcount30_37rn_core_193;
  wire popcount30_37rn_core_194;
  wire popcount30_37rn_core_195;
  wire popcount30_37rn_core_197;
  wire popcount30_37rn_core_198;
  wire popcount30_37rn_core_199;
  wire popcount30_37rn_core_201;
  wire popcount30_37rn_core_203;
  wire popcount30_37rn_core_204;
  wire popcount30_37rn_core_205;
  wire popcount30_37rn_core_206;
  wire popcount30_37rn_core_208;
  wire popcount30_37rn_core_209;
  wire popcount30_37rn_core_210;
  wire popcount30_37rn_core_212;

  assign popcount30_37rn_core_032 = input_a[6] & input_a[8];
  assign popcount30_37rn_core_033 = ~input_a[24];
  assign popcount30_37rn_core_034 = ~input_a[23];
  assign popcount30_37rn_core_035 = ~(input_a[1] | input_a[20]);
  assign popcount30_37rn_core_038 = input_a[10] ^ input_a[18];
  assign popcount30_37rn_core_039 = input_a[11] ^ input_a[3];
  assign popcount30_37rn_core_040 = ~(input_a[21] | input_a[9]);
  assign popcount30_37rn_core_043 = ~(input_a[15] | input_a[25]);
  assign popcount30_37rn_core_044 = ~(input_a[4] ^ input_a[23]);
  assign popcount30_37rn_core_046 = ~input_a[22];
  assign popcount30_37rn_core_047 = ~(input_a[12] ^ input_a[10]);
  assign popcount30_37rn_core_049 = ~input_a[13];
  assign popcount30_37rn_core_051 = input_a[24] | input_a[5];
  assign popcount30_37rn_core_054 = input_a[10] | input_a[18];
  assign popcount30_37rn_core_056 = ~(input_a[29] | input_a[22]);
  assign popcount30_37rn_core_057_not = ~input_a[15];
  assign popcount30_37rn_core_059 = ~input_a[5];
  assign popcount30_37rn_core_062 = input_a[25] ^ input_a[6];
  assign popcount30_37rn_core_065 = input_a[18] & input_a[26];
  assign popcount30_37rn_core_066 = input_a[24] | input_a[7];
  assign popcount30_37rn_core_067 = ~(input_a[24] | input_a[17]);
  assign popcount30_37rn_core_069 = ~(input_a[19] | input_a[13]);
  assign popcount30_37rn_core_072 = ~(input_a[22] | input_a[2]);
  assign popcount30_37rn_core_074 = ~input_a[26];
  assign popcount30_37rn_core_076 = input_a[29] ^ input_a[2];
  assign popcount30_37rn_core_080 = ~(input_a[26] | input_a[22]);
  assign popcount30_37rn_core_082 = ~(input_a[1] & input_a[13]);
  assign popcount30_37rn_core_083 = ~(input_a[20] | input_a[25]);
  assign popcount30_37rn_core_085 = ~(input_a[0] ^ input_a[6]);
  assign popcount30_37rn_core_086 = ~input_a[25];
  assign popcount30_37rn_core_087 = input_a[11] ^ input_a[25];
  assign popcount30_37rn_core_089 = input_a[23] & input_a[22];
  assign popcount30_37rn_core_092_not = ~input_a[22];
  assign popcount30_37rn_core_093 = ~(input_a[23] & input_a[20]);
  assign popcount30_37rn_core_094 = ~(input_a[5] ^ input_a[25]);
  assign popcount30_37rn_core_095 = ~(input_a[25] & input_a[1]);
  assign popcount30_37rn_core_098 = ~input_a[21];
  assign popcount30_37rn_core_099 = ~(input_a[5] | input_a[6]);
  assign popcount30_37rn_core_101 = input_a[0] ^ input_a[9];
  assign popcount30_37rn_core_102 = input_a[12] ^ input_a[20];
  assign popcount30_37rn_core_107 = ~(input_a[28] ^ input_a[22]);
  assign popcount30_37rn_core_108 = ~(input_a[26] ^ input_a[6]);
  assign popcount30_37rn_core_109 = input_a[15] ^ input_a[28];
  assign popcount30_37rn_core_111 = ~(input_a[0] ^ input_a[12]);
  assign popcount30_37rn_core_113 = input_a[3] | input_a[15];
  assign popcount30_37rn_core_115 = ~(input_a[18] | input_a[0]);
  assign popcount30_37rn_core_116 = ~input_a[7];
  assign popcount30_37rn_core_117 = ~(input_a[4] ^ input_a[23]);
  assign popcount30_37rn_core_120 = ~(input_a[6] ^ input_a[23]);
  assign popcount30_37rn_core_121 = ~(input_a[13] & input_a[20]);
  assign popcount30_37rn_core_122 = ~(input_a[28] ^ input_a[21]);
  assign popcount30_37rn_core_123_not = ~input_a[24];
  assign popcount30_37rn_core_125 = input_a[24] | input_a[0];
  assign popcount30_37rn_core_126 = input_a[19] ^ input_a[3];
  assign popcount30_37rn_core_127 = input_a[22] | input_a[27];
  assign popcount30_37rn_core_128 = ~(input_a[6] | input_a[10]);
  assign popcount30_37rn_core_130 = ~input_a[12];
  assign popcount30_37rn_core_131 = ~(input_a[24] & input_a[20]);
  assign popcount30_37rn_core_132 = input_a[12] ^ input_a[3];
  assign popcount30_37rn_core_135 = ~(input_a[17] & input_a[24]);
  assign popcount30_37rn_core_137 = ~(input_a[12] ^ input_a[6]);
  assign popcount30_37rn_core_138 = input_a[16] & input_a[26];
  assign popcount30_37rn_core_139 = ~(input_a[14] & input_a[15]);
  assign popcount30_37rn_core_141 = ~(input_a[22] | input_a[3]);
  assign popcount30_37rn_core_142 = ~(input_a[11] | input_a[29]);
  assign popcount30_37rn_core_143 = ~input_a[17];
  assign popcount30_37rn_core_144 = ~input_a[5];
  assign popcount30_37rn_core_146 = ~(input_a[17] ^ input_a[28]);
  assign popcount30_37rn_core_147 = ~(input_a[8] ^ input_a[15]);
  assign popcount30_37rn_core_149 = input_a[18] & input_a[15];
  assign popcount30_37rn_core_150_not = ~input_a[10];
  assign popcount30_37rn_core_152 = ~(input_a[27] & input_a[13]);
  assign popcount30_37rn_core_153 = ~(input_a[23] & input_a[29]);
  assign popcount30_37rn_core_156 = ~(input_a[22] & input_a[10]);
  assign popcount30_37rn_core_157 = ~(input_a[25] & input_a[5]);
  assign popcount30_37rn_core_158 = ~input_a[4];
  assign popcount30_37rn_core_159 = input_a[1] | input_a[6];
  assign popcount30_37rn_core_160 = ~(input_a[13] & input_a[28]);
  assign popcount30_37rn_core_162 = ~input_a[13];
  assign popcount30_37rn_core_163 = input_a[28] ^ input_a[12];
  assign popcount30_37rn_core_164 = input_a[15] ^ input_a[2];
  assign popcount30_37rn_core_165 = input_a[15] | input_a[18];
  assign popcount30_37rn_core_167 = ~input_a[6];
  assign popcount30_37rn_core_168_not = ~input_a[10];
  assign popcount30_37rn_core_170 = ~(input_a[26] & input_a[17]);
  assign popcount30_37rn_core_171 = input_a[18] | input_a[2];
  assign popcount30_37rn_core_172 = ~(input_a[28] & input_a[28]);
  assign popcount30_37rn_core_173 = input_a[3] | input_a[13];
  assign popcount30_37rn_core_175 = ~(input_a[7] & input_a[28]);
  assign popcount30_37rn_core_177 = input_a[17] ^ input_a[13];
  assign popcount30_37rn_core_178 = input_a[2] | input_a[16];
  assign popcount30_37rn_core_179 = input_a[20] | input_a[13];
  assign popcount30_37rn_core_180 = ~(input_a[16] ^ input_a[21]);
  assign popcount30_37rn_core_181 = input_a[25] ^ input_a[8];
  assign popcount30_37rn_core_182_not = ~input_a[3];
  assign popcount30_37rn_core_184 = input_a[8] & input_a[21];
  assign popcount30_37rn_core_185 = ~(input_a[26] ^ input_a[8]);
  assign popcount30_37rn_core_187 = ~(input_a[17] | input_a[12]);
  assign popcount30_37rn_core_188 = input_a[2] ^ input_a[16];
  assign popcount30_37rn_core_189 = ~(input_a[23] ^ input_a[28]);
  assign popcount30_37rn_core_190 = input_a[7] ^ input_a[5];
  assign popcount30_37rn_core_191 = ~(input_a[9] | input_a[27]);
  assign popcount30_37rn_core_193 = input_a[14] & input_a[1];
  assign popcount30_37rn_core_194 = input_a[3] & input_a[17];
  assign popcount30_37rn_core_195 = ~(input_a[12] ^ input_a[22]);
  assign popcount30_37rn_core_197 = ~(input_a[2] | input_a[1]);
  assign popcount30_37rn_core_198 = input_a[26] | input_a[17];
  assign popcount30_37rn_core_199 = ~(input_a[15] & input_a[4]);
  assign popcount30_37rn_core_201 = ~(input_a[20] ^ input_a[25]);
  assign popcount30_37rn_core_203 = ~input_a[25];
  assign popcount30_37rn_core_204 = input_a[12] & input_a[2];
  assign popcount30_37rn_core_205 = ~(input_a[10] & input_a[9]);
  assign popcount30_37rn_core_206 = input_a[28] & input_a[12];
  assign popcount30_37rn_core_208 = ~(input_a[24] & input_a[22]);
  assign popcount30_37rn_core_209 = ~(input_a[13] | input_a[25]);
  assign popcount30_37rn_core_210 = ~(input_a[24] | input_a[23]);
  assign popcount30_37rn_core_212 = input_a[5] ^ input_a[29];

  assign popcount30_37rn_out[0] = 1'b1;
  assign popcount30_37rn_out[1] = input_a[28];
  assign popcount30_37rn_out[2] = input_a[10];
  assign popcount30_37rn_out[3] = 1'b0;
  assign popcount30_37rn_out[4] = 1'b1;
endmodule