// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.244
// WCE=6.0
// EP=0.753931%
// Printed PDK parameters:
//  Area=35697113.0
//  Delay=48375384.0
//  Power=1881900.0

module popcount25_qjqh(input [24:0] input_a, output [4:0] popcount25_qjqh_out);
  wire popcount25_qjqh_core_028;
  wire popcount25_qjqh_core_032;
  wire popcount25_qjqh_core_033;
  wire popcount25_qjqh_core_034;
  wire popcount25_qjqh_core_035;
  wire popcount25_qjqh_core_036;
  wire popcount25_qjqh_core_037;
  wire popcount25_qjqh_core_038;
  wire popcount25_qjqh_core_039;
  wire popcount25_qjqh_core_041;
  wire popcount25_qjqh_core_042;
  wire popcount25_qjqh_core_043;
  wire popcount25_qjqh_core_044;
  wire popcount25_qjqh_core_045;
  wire popcount25_qjqh_core_047_not;
  wire popcount25_qjqh_core_050;
  wire popcount25_qjqh_core_051;
  wire popcount25_qjqh_core_052;
  wire popcount25_qjqh_core_053_not;
  wire popcount25_qjqh_core_054;
  wire popcount25_qjqh_core_055;
  wire popcount25_qjqh_core_056;
  wire popcount25_qjqh_core_057;
  wire popcount25_qjqh_core_058;
  wire popcount25_qjqh_core_059;
  wire popcount25_qjqh_core_060;
  wire popcount25_qjqh_core_061;
  wire popcount25_qjqh_core_063;
  wire popcount25_qjqh_core_064;
  wire popcount25_qjqh_core_065;
  wire popcount25_qjqh_core_067;
  wire popcount25_qjqh_core_069;
  wire popcount25_qjqh_core_071;
  wire popcount25_qjqh_core_074;
  wire popcount25_qjqh_core_075;
  wire popcount25_qjqh_core_077;
  wire popcount25_qjqh_core_078;
  wire popcount25_qjqh_core_080;
  wire popcount25_qjqh_core_082;
  wire popcount25_qjqh_core_083;
  wire popcount25_qjqh_core_084;
  wire popcount25_qjqh_core_085;
  wire popcount25_qjqh_core_086;
  wire popcount25_qjqh_core_090;
  wire popcount25_qjqh_core_092;
  wire popcount25_qjqh_core_093;
  wire popcount25_qjqh_core_095;
  wire popcount25_qjqh_core_096;
  wire popcount25_qjqh_core_097;
  wire popcount25_qjqh_core_098;
  wire popcount25_qjqh_core_099;
  wire popcount25_qjqh_core_100;
  wire popcount25_qjqh_core_101;
  wire popcount25_qjqh_core_102;
  wire popcount25_qjqh_core_104;
  wire popcount25_qjqh_core_105;
  wire popcount25_qjqh_core_106;
  wire popcount25_qjqh_core_107;
  wire popcount25_qjqh_core_109_not;
  wire popcount25_qjqh_core_112;
  wire popcount25_qjqh_core_114;
  wire popcount25_qjqh_core_116;
  wire popcount25_qjqh_core_117;
  wire popcount25_qjqh_core_119;
  wire popcount25_qjqh_core_120;
  wire popcount25_qjqh_core_121;
  wire popcount25_qjqh_core_122;
  wire popcount25_qjqh_core_123;
  wire popcount25_qjqh_core_124;
  wire popcount25_qjqh_core_125;
  wire popcount25_qjqh_core_126;
  wire popcount25_qjqh_core_128;
  wire popcount25_qjqh_core_131_not;
  wire popcount25_qjqh_core_132;
  wire popcount25_qjqh_core_133;
  wire popcount25_qjqh_core_134;
  wire popcount25_qjqh_core_135;
  wire popcount25_qjqh_core_136;
  wire popcount25_qjqh_core_143;
  wire popcount25_qjqh_core_144;
  wire popcount25_qjqh_core_145;
  wire popcount25_qjqh_core_146;
  wire popcount25_qjqh_core_147;
  wire popcount25_qjqh_core_149;
  wire popcount25_qjqh_core_151;
  wire popcount25_qjqh_core_152;
  wire popcount25_qjqh_core_153;
  wire popcount25_qjqh_core_154;
  wire popcount25_qjqh_core_155;
  wire popcount25_qjqh_core_156;
  wire popcount25_qjqh_core_160;
  wire popcount25_qjqh_core_162;
  wire popcount25_qjqh_core_163;
  wire popcount25_qjqh_core_164;
  wire popcount25_qjqh_core_165;
  wire popcount25_qjqh_core_166;
  wire popcount25_qjqh_core_169;
  wire popcount25_qjqh_core_170;
  wire popcount25_qjqh_core_171;
  wire popcount25_qjqh_core_172;
  wire popcount25_qjqh_core_173;
  wire popcount25_qjqh_core_174;
  wire popcount25_qjqh_core_175;
  wire popcount25_qjqh_core_176;
  wire popcount25_qjqh_core_177;
  wire popcount25_qjqh_core_178;
  wire popcount25_qjqh_core_179;
  wire popcount25_qjqh_core_180;
  wire popcount25_qjqh_core_182;

  assign popcount25_qjqh_core_028 = input_a[12] & input_a[2];
  assign popcount25_qjqh_core_032 = input_a[16] & input_a[14];
  assign popcount25_qjqh_core_033 = input_a[4] ^ input_a[5];
  assign popcount25_qjqh_core_034 = input_a[4] & input_a[5];
  assign popcount25_qjqh_core_035 = input_a[3] ^ popcount25_qjqh_core_033;
  assign popcount25_qjqh_core_036 = input_a[3] & popcount25_qjqh_core_033;
  assign popcount25_qjqh_core_037 = popcount25_qjqh_core_034 | popcount25_qjqh_core_036;
  assign popcount25_qjqh_core_038 = input_a[9] & input_a[20];
  assign popcount25_qjqh_core_039 = ~input_a[15];
  assign popcount25_qjqh_core_041 = popcount25_qjqh_core_028 ^ popcount25_qjqh_core_037;
  assign popcount25_qjqh_core_042 = popcount25_qjqh_core_028 & popcount25_qjqh_core_037;
  assign popcount25_qjqh_core_043 = popcount25_qjqh_core_041 ^ popcount25_qjqh_core_035;
  assign popcount25_qjqh_core_044 = popcount25_qjqh_core_041 & popcount25_qjqh_core_035;
  assign popcount25_qjqh_core_045 = popcount25_qjqh_core_042 | popcount25_qjqh_core_044;
  assign popcount25_qjqh_core_047_not = ~input_a[18];
  assign popcount25_qjqh_core_050 = ~(input_a[16] ^ input_a[14]);
  assign popcount25_qjqh_core_051 = input_a[7] | input_a[8];
  assign popcount25_qjqh_core_052 = input_a[7] & input_a[8];
  assign popcount25_qjqh_core_053_not = ~input_a[20];
  assign popcount25_qjqh_core_054 = input_a[6] & popcount25_qjqh_core_051;
  assign popcount25_qjqh_core_055 = popcount25_qjqh_core_052 | popcount25_qjqh_core_054;
  assign popcount25_qjqh_core_056 = input_a[21] ^ input_a[2];
  assign popcount25_qjqh_core_057 = input_a[10] | input_a[11];
  assign popcount25_qjqh_core_058 = input_a[10] & input_a[11];
  assign popcount25_qjqh_core_059 = input_a[5] | input_a[10];
  assign popcount25_qjqh_core_060 = input_a[9] & popcount25_qjqh_core_057;
  assign popcount25_qjqh_core_061 = popcount25_qjqh_core_058 | popcount25_qjqh_core_060;
  assign popcount25_qjqh_core_063 = input_a[16] | input_a[13];
  assign popcount25_qjqh_core_064 = ~(input_a[20] & input_a[9]);
  assign popcount25_qjqh_core_065 = popcount25_qjqh_core_055 ^ popcount25_qjqh_core_061;
  assign popcount25_qjqh_core_067 = ~popcount25_qjqh_core_065;
  assign popcount25_qjqh_core_069 = popcount25_qjqh_core_055 | popcount25_qjqh_core_065;
  assign popcount25_qjqh_core_071 = ~input_a[1];
  assign popcount25_qjqh_core_074 = input_a[19] ^ input_a[6];
  assign popcount25_qjqh_core_075 = input_a[5] | input_a[16];
  assign popcount25_qjqh_core_077 = popcount25_qjqh_core_043 ^ popcount25_qjqh_core_067;
  assign popcount25_qjqh_core_078 = popcount25_qjqh_core_043 & popcount25_qjqh_core_067;
  assign popcount25_qjqh_core_080 = ~(input_a[0] ^ input_a[16]);
  assign popcount25_qjqh_core_082 = popcount25_qjqh_core_045 ^ popcount25_qjqh_core_069;
  assign popcount25_qjqh_core_083 = popcount25_qjqh_core_045 & popcount25_qjqh_core_069;
  assign popcount25_qjqh_core_084 = popcount25_qjqh_core_082 ^ popcount25_qjqh_core_078;
  assign popcount25_qjqh_core_085 = popcount25_qjqh_core_082 & popcount25_qjqh_core_078;
  assign popcount25_qjqh_core_086 = popcount25_qjqh_core_083 | popcount25_qjqh_core_085;
  assign popcount25_qjqh_core_090 = input_a[2] | input_a[22];
  assign popcount25_qjqh_core_092 = input_a[13] | input_a[14];
  assign popcount25_qjqh_core_093 = input_a[13] & input_a[14];
  assign popcount25_qjqh_core_095 = input_a[0] & popcount25_qjqh_core_092;
  assign popcount25_qjqh_core_096 = popcount25_qjqh_core_093 | popcount25_qjqh_core_095;
  assign popcount25_qjqh_core_097 = ~(input_a[2] | input_a[9]);
  assign popcount25_qjqh_core_098 = input_a[3] | input_a[7];
  assign popcount25_qjqh_core_099 = input_a[17] & input_a[16];
  assign popcount25_qjqh_core_100 = input_a[3] | input_a[21];
  assign popcount25_qjqh_core_101 = input_a[17] & input_a[15];
  assign popcount25_qjqh_core_102 = popcount25_qjqh_core_099 | popcount25_qjqh_core_101;
  assign popcount25_qjqh_core_104 = ~(input_a[15] ^ input_a[16]);
  assign popcount25_qjqh_core_105 = ~(input_a[23] | input_a[4]);
  assign popcount25_qjqh_core_106 = popcount25_qjqh_core_096 ^ popcount25_qjqh_core_102;
  assign popcount25_qjqh_core_107 = popcount25_qjqh_core_096 & popcount25_qjqh_core_102;
  assign popcount25_qjqh_core_109_not = ~input_a[3];
  assign popcount25_qjqh_core_112 = input_a[11] & input_a[14];
  assign popcount25_qjqh_core_114 = input_a[14] & input_a[19];
  assign popcount25_qjqh_core_116 = input_a[22] & input_a[17];
  assign popcount25_qjqh_core_117 = input_a[19] & input_a[20];
  assign popcount25_qjqh_core_119 = input_a[18] & input_a[1];
  assign popcount25_qjqh_core_120 = popcount25_qjqh_core_117 | popcount25_qjqh_core_119;
  assign popcount25_qjqh_core_121 = input_a[14] & input_a[24];
  assign popcount25_qjqh_core_122 = ~(input_a[17] ^ input_a[0]);
  assign popcount25_qjqh_core_123 = input_a[21] & input_a[22];
  assign popcount25_qjqh_core_124 = ~(input_a[17] | input_a[10]);
  assign popcount25_qjqh_core_125 = input_a[23] & input_a[24];
  assign popcount25_qjqh_core_126 = input_a[21] | input_a[3];
  assign popcount25_qjqh_core_128 = popcount25_qjqh_core_123 | popcount25_qjqh_core_125;
  assign popcount25_qjqh_core_131_not = ~input_a[1];
  assign popcount25_qjqh_core_132 = ~input_a[24];
  assign popcount25_qjqh_core_133 = input_a[6] | input_a[12];
  assign popcount25_qjqh_core_134 = ~(input_a[22] ^ input_a[21]);
  assign popcount25_qjqh_core_135 = popcount25_qjqh_core_120 ^ popcount25_qjqh_core_128;
  assign popcount25_qjqh_core_136 = popcount25_qjqh_core_120 & popcount25_qjqh_core_128;
  assign popcount25_qjqh_core_143 = ~input_a[8];
  assign popcount25_qjqh_core_144 = ~input_a[2];
  assign popcount25_qjqh_core_145 = input_a[8] | input_a[13];
  assign popcount25_qjqh_core_146 = input_a[22] ^ input_a[9];
  assign popcount25_qjqh_core_147 = popcount25_qjqh_core_106 ^ popcount25_qjqh_core_135;
  assign popcount25_qjqh_core_149 = ~popcount25_qjqh_core_147;
  assign popcount25_qjqh_core_151 = popcount25_qjqh_core_106 | popcount25_qjqh_core_147;
  assign popcount25_qjqh_core_152 = popcount25_qjqh_core_107 ^ popcount25_qjqh_core_136;
  assign popcount25_qjqh_core_153 = popcount25_qjqh_core_107 & popcount25_qjqh_core_136;
  assign popcount25_qjqh_core_154 = popcount25_qjqh_core_152 ^ popcount25_qjqh_core_151;
  assign popcount25_qjqh_core_155 = popcount25_qjqh_core_152 & popcount25_qjqh_core_151;
  assign popcount25_qjqh_core_156 = popcount25_qjqh_core_153 | popcount25_qjqh_core_155;
  assign popcount25_qjqh_core_160 = input_a[13] | input_a[8];
  assign popcount25_qjqh_core_162 = input_a[17] ^ input_a[15];
  assign popcount25_qjqh_core_163 = ~(input_a[22] | input_a[15]);
  assign popcount25_qjqh_core_164 = popcount25_qjqh_core_077 ^ popcount25_qjqh_core_149;
  assign popcount25_qjqh_core_165 = popcount25_qjqh_core_077 & popcount25_qjqh_core_149;
  assign popcount25_qjqh_core_166 = ~(input_a[16] & input_a[12]);
  assign popcount25_qjqh_core_169 = popcount25_qjqh_core_084 ^ popcount25_qjqh_core_154;
  assign popcount25_qjqh_core_170 = popcount25_qjqh_core_084 & popcount25_qjqh_core_154;
  assign popcount25_qjqh_core_171 = popcount25_qjqh_core_169 ^ popcount25_qjqh_core_165;
  assign popcount25_qjqh_core_172 = popcount25_qjqh_core_169 & popcount25_qjqh_core_165;
  assign popcount25_qjqh_core_173 = popcount25_qjqh_core_170 | popcount25_qjqh_core_172;
  assign popcount25_qjqh_core_174 = popcount25_qjqh_core_086 ^ popcount25_qjqh_core_156;
  assign popcount25_qjqh_core_175 = popcount25_qjqh_core_086 & popcount25_qjqh_core_156;
  assign popcount25_qjqh_core_176 = popcount25_qjqh_core_174 ^ popcount25_qjqh_core_173;
  assign popcount25_qjqh_core_177 = popcount25_qjqh_core_174 & popcount25_qjqh_core_173;
  assign popcount25_qjqh_core_178 = popcount25_qjqh_core_175 | popcount25_qjqh_core_177;
  assign popcount25_qjqh_core_179 = ~(input_a[17] ^ input_a[16]);
  assign popcount25_qjqh_core_180 = input_a[5] | input_a[22];
  assign popcount25_qjqh_core_182 = ~input_a[2];

  assign popcount25_qjqh_out[0] = popcount25_qjqh_core_173;
  assign popcount25_qjqh_out[1] = popcount25_qjqh_core_164;
  assign popcount25_qjqh_out[2] = popcount25_qjqh_core_171;
  assign popcount25_qjqh_out[3] = popcount25_qjqh_core_176;
  assign popcount25_qjqh_out[4] = popcount25_qjqh_core_178;
endmodule