// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.89676
// WCE=17.0
// EP=0.893849%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_22bo(input [28:0] input_a, output [4:0] popcount29_22bo_out);
  wire popcount29_22bo_core_034;
  wire popcount29_22bo_core_035;
  wire popcount29_22bo_core_036;
  wire popcount29_22bo_core_039;
  wire popcount29_22bo_core_040;
  wire popcount29_22bo_core_041;
  wire popcount29_22bo_core_042;
  wire popcount29_22bo_core_043_not;
  wire popcount29_22bo_core_044;
  wire popcount29_22bo_core_045;
  wire popcount29_22bo_core_046;
  wire popcount29_22bo_core_047;
  wire popcount29_22bo_core_048;
  wire popcount29_22bo_core_053;
  wire popcount29_22bo_core_054;
  wire popcount29_22bo_core_055;
  wire popcount29_22bo_core_057;
  wire popcount29_22bo_core_061;
  wire popcount29_22bo_core_062;
  wire popcount29_22bo_core_063;
  wire popcount29_22bo_core_064;
  wire popcount29_22bo_core_065;
  wire popcount29_22bo_core_066;
  wire popcount29_22bo_core_067;
  wire popcount29_22bo_core_068;
  wire popcount29_22bo_core_069;
  wire popcount29_22bo_core_070_not;
  wire popcount29_22bo_core_072;
  wire popcount29_22bo_core_074;
  wire popcount29_22bo_core_075;
  wire popcount29_22bo_core_076;
  wire popcount29_22bo_core_079;
  wire popcount29_22bo_core_080;
  wire popcount29_22bo_core_081;
  wire popcount29_22bo_core_082;
  wire popcount29_22bo_core_084;
  wire popcount29_22bo_core_086;
  wire popcount29_22bo_core_090;
  wire popcount29_22bo_core_091;
  wire popcount29_22bo_core_092;
  wire popcount29_22bo_core_094;
  wire popcount29_22bo_core_096;
  wire popcount29_22bo_core_097;
  wire popcount29_22bo_core_099;
  wire popcount29_22bo_core_100_not;
  wire popcount29_22bo_core_102;
  wire popcount29_22bo_core_103;
  wire popcount29_22bo_core_104;
  wire popcount29_22bo_core_105;
  wire popcount29_22bo_core_107;
  wire popcount29_22bo_core_108;
  wire popcount29_22bo_core_109;
  wire popcount29_22bo_core_110;
  wire popcount29_22bo_core_111;
  wire popcount29_22bo_core_113;
  wire popcount29_22bo_core_117;
  wire popcount29_22bo_core_122;
  wire popcount29_22bo_core_123;
  wire popcount29_22bo_core_124;
  wire popcount29_22bo_core_125;
  wire popcount29_22bo_core_126;
  wire popcount29_22bo_core_128;
  wire popcount29_22bo_core_129;
  wire popcount29_22bo_core_132;
  wire popcount29_22bo_core_136;
  wire popcount29_22bo_core_137;
  wire popcount29_22bo_core_138;
  wire popcount29_22bo_core_139;
  wire popcount29_22bo_core_141;
  wire popcount29_22bo_core_142;
  wire popcount29_22bo_core_143;
  wire popcount29_22bo_core_146;
  wire popcount29_22bo_core_148;
  wire popcount29_22bo_core_152;
  wire popcount29_22bo_core_153;
  wire popcount29_22bo_core_154;
  wire popcount29_22bo_core_156;
  wire popcount29_22bo_core_157;
  wire popcount29_22bo_core_160;
  wire popcount29_22bo_core_161;
  wire popcount29_22bo_core_163;
  wire popcount29_22bo_core_164;
  wire popcount29_22bo_core_165;
  wire popcount29_22bo_core_166;
  wire popcount29_22bo_core_170;
  wire popcount29_22bo_core_172;
  wire popcount29_22bo_core_173;
  wire popcount29_22bo_core_174;
  wire popcount29_22bo_core_176;
  wire popcount29_22bo_core_178;
  wire popcount29_22bo_core_179;
  wire popcount29_22bo_core_181;
  wire popcount29_22bo_core_183;
  wire popcount29_22bo_core_184;
  wire popcount29_22bo_core_185;
  wire popcount29_22bo_core_186;
  wire popcount29_22bo_core_187;
  wire popcount29_22bo_core_190_not;
  wire popcount29_22bo_core_192;
  wire popcount29_22bo_core_195;
  wire popcount29_22bo_core_196;
  wire popcount29_22bo_core_199;
  wire popcount29_22bo_core_200;
  wire popcount29_22bo_core_201;
  wire popcount29_22bo_core_204;
  wire popcount29_22bo_core_205;
  wire popcount29_22bo_core_206;
  wire popcount29_22bo_core_207;

  assign popcount29_22bo_core_034 = input_a[24] & input_a[26];
  assign popcount29_22bo_core_035 = ~(input_a[0] & input_a[8]);
  assign popcount29_22bo_core_036 = ~input_a[16];
  assign popcount29_22bo_core_039 = input_a[6] & input_a[2];
  assign popcount29_22bo_core_040 = ~(input_a[22] | input_a[6]);
  assign popcount29_22bo_core_041 = input_a[27] | input_a[17];
  assign popcount29_22bo_core_042 = ~input_a[0];
  assign popcount29_22bo_core_043_not = ~input_a[25];
  assign popcount29_22bo_core_044 = input_a[21] | input_a[5];
  assign popcount29_22bo_core_045 = ~(input_a[5] & input_a[26]);
  assign popcount29_22bo_core_046 = input_a[9] ^ input_a[3];
  assign popcount29_22bo_core_047 = ~(input_a[12] & input_a[21]);
  assign popcount29_22bo_core_048 = ~input_a[9];
  assign popcount29_22bo_core_053 = input_a[9] | input_a[21];
  assign popcount29_22bo_core_054 = input_a[28] & input_a[23];
  assign popcount29_22bo_core_055 = input_a[2] & input_a[17];
  assign popcount29_22bo_core_057 = input_a[2] & input_a[4];
  assign popcount29_22bo_core_061 = ~(input_a[19] & input_a[6]);
  assign popcount29_22bo_core_062 = ~(input_a[26] & input_a[23]);
  assign popcount29_22bo_core_063 = input_a[15] ^ input_a[24];
  assign popcount29_22bo_core_064 = input_a[18] | input_a[5];
  assign popcount29_22bo_core_065 = ~input_a[6];
  assign popcount29_22bo_core_066 = ~(input_a[22] & input_a[11]);
  assign popcount29_22bo_core_067 = input_a[21] & input_a[22];
  assign popcount29_22bo_core_068 = ~(input_a[27] & input_a[17]);
  assign popcount29_22bo_core_069 = ~input_a[8];
  assign popcount29_22bo_core_070_not = ~input_a[24];
  assign popcount29_22bo_core_072 = input_a[1] | input_a[12];
  assign popcount29_22bo_core_074 = ~input_a[24];
  assign popcount29_22bo_core_075 = ~input_a[3];
  assign popcount29_22bo_core_076 = ~input_a[20];
  assign popcount29_22bo_core_079 = input_a[8] ^ input_a[28];
  assign popcount29_22bo_core_080 = ~input_a[20];
  assign popcount29_22bo_core_081 = ~(input_a[16] | input_a[4]);
  assign popcount29_22bo_core_082 = ~(input_a[11] & input_a[26]);
  assign popcount29_22bo_core_084 = input_a[19] | input_a[28];
  assign popcount29_22bo_core_086 = ~(input_a[4] & input_a[0]);
  assign popcount29_22bo_core_090 = input_a[1] | input_a[17];
  assign popcount29_22bo_core_091 = ~(input_a[5] & input_a[20]);
  assign popcount29_22bo_core_092 = input_a[3] | input_a[28];
  assign popcount29_22bo_core_094 = ~(input_a[6] & input_a[24]);
  assign popcount29_22bo_core_096 = ~(input_a[8] | input_a[26]);
  assign popcount29_22bo_core_097 = ~(input_a[4] | input_a[21]);
  assign popcount29_22bo_core_099 = input_a[15] | input_a[22];
  assign popcount29_22bo_core_100_not = ~input_a[15];
  assign popcount29_22bo_core_102 = ~(input_a[4] & input_a[8]);
  assign popcount29_22bo_core_103 = input_a[14] ^ input_a[20];
  assign popcount29_22bo_core_104 = input_a[7] | input_a[19];
  assign popcount29_22bo_core_105 = ~(input_a[12] ^ input_a[21]);
  assign popcount29_22bo_core_107 = ~(input_a[14] & input_a[12]);
  assign popcount29_22bo_core_108 = input_a[15] ^ input_a[11];
  assign popcount29_22bo_core_109 = ~(input_a[17] ^ input_a[5]);
  assign popcount29_22bo_core_110 = input_a[21] | input_a[11];
  assign popcount29_22bo_core_111 = ~(input_a[16] ^ input_a[10]);
  assign popcount29_22bo_core_113 = input_a[6] ^ input_a[12];
  assign popcount29_22bo_core_117 = ~(input_a[25] & input_a[18]);
  assign popcount29_22bo_core_122 = ~(input_a[2] ^ input_a[25]);
  assign popcount29_22bo_core_123 = ~(input_a[7] | input_a[27]);
  assign popcount29_22bo_core_124 = ~(input_a[24] & input_a[23]);
  assign popcount29_22bo_core_125 = input_a[28] ^ input_a[14];
  assign popcount29_22bo_core_126 = ~(input_a[16] ^ input_a[19]);
  assign popcount29_22bo_core_128 = ~(input_a[1] | input_a[1]);
  assign popcount29_22bo_core_129 = input_a[22] ^ input_a[4];
  assign popcount29_22bo_core_132 = ~input_a[26];
  assign popcount29_22bo_core_136 = ~input_a[21];
  assign popcount29_22bo_core_137 = input_a[14] ^ input_a[24];
  assign popcount29_22bo_core_138 = input_a[10] ^ input_a[15];
  assign popcount29_22bo_core_139 = input_a[0] ^ input_a[6];
  assign popcount29_22bo_core_141 = ~(input_a[0] ^ input_a[26]);
  assign popcount29_22bo_core_142 = input_a[24] & input_a[27];
  assign popcount29_22bo_core_143 = ~(input_a[16] | input_a[9]);
  assign popcount29_22bo_core_146 = input_a[7] | input_a[22];
  assign popcount29_22bo_core_148 = ~input_a[26];
  assign popcount29_22bo_core_152 = ~(input_a[25] | input_a[3]);
  assign popcount29_22bo_core_153 = input_a[8] ^ input_a[17];
  assign popcount29_22bo_core_154 = input_a[8] | input_a[13];
  assign popcount29_22bo_core_156 = ~(input_a[25] & input_a[6]);
  assign popcount29_22bo_core_157 = ~(input_a[10] & input_a[27]);
  assign popcount29_22bo_core_160 = input_a[16] ^ input_a[24];
  assign popcount29_22bo_core_161 = ~(input_a[28] | input_a[10]);
  assign popcount29_22bo_core_163 = ~(input_a[9] & input_a[27]);
  assign popcount29_22bo_core_164 = ~(input_a[5] ^ input_a[26]);
  assign popcount29_22bo_core_165 = input_a[10] | input_a[24];
  assign popcount29_22bo_core_166 = input_a[2] ^ input_a[24];
  assign popcount29_22bo_core_170 = input_a[15] & input_a[12];
  assign popcount29_22bo_core_172 = ~input_a[9];
  assign popcount29_22bo_core_173 = ~(input_a[16] | input_a[7]);
  assign popcount29_22bo_core_174 = input_a[8] & input_a[23];
  assign popcount29_22bo_core_176 = ~(input_a[20] ^ input_a[22]);
  assign popcount29_22bo_core_178 = input_a[12] | input_a[9];
  assign popcount29_22bo_core_179 = ~(input_a[21] | input_a[22]);
  assign popcount29_22bo_core_181 = input_a[9] | input_a[2];
  assign popcount29_22bo_core_183 = ~(input_a[10] & input_a[28]);
  assign popcount29_22bo_core_184 = ~(input_a[25] | input_a[26]);
  assign popcount29_22bo_core_185 = input_a[4] | input_a[16];
  assign popcount29_22bo_core_186 = ~(input_a[10] & input_a[18]);
  assign popcount29_22bo_core_187 = ~(input_a[14] | input_a[26]);
  assign popcount29_22bo_core_190_not = ~input_a[17];
  assign popcount29_22bo_core_192 = input_a[3] & input_a[6];
  assign popcount29_22bo_core_195 = ~(input_a[6] | input_a[26]);
  assign popcount29_22bo_core_196 = input_a[13] ^ input_a[7];
  assign popcount29_22bo_core_199 = ~(input_a[14] | input_a[16]);
  assign popcount29_22bo_core_200 = ~(input_a[21] ^ input_a[3]);
  assign popcount29_22bo_core_201 = ~(input_a[25] ^ input_a[5]);
  assign popcount29_22bo_core_204 = ~(input_a[5] & input_a[25]);
  assign popcount29_22bo_core_205 = ~(input_a[21] ^ input_a[6]);
  assign popcount29_22bo_core_206 = input_a[18] & input_a[2];
  assign popcount29_22bo_core_207 = input_a[1] & input_a[12];

  assign popcount29_22bo_out[0] = input_a[13];
  assign popcount29_22bo_out[1] = 1'b1;
  assign popcount29_22bo_out[2] = input_a[26];
  assign popcount29_22bo_out[3] = 1'b1;
  assign popcount29_22bo_out[4] = 1'b0;
endmodule