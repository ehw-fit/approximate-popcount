// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.32472
// WCE=14.0
// EP=0.867159%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_gm8j(input [24:0] input_a, output [4:0] popcount25_gm8j_out);
  wire popcount25_gm8j_core_028;
  wire popcount25_gm8j_core_029;
  wire popcount25_gm8j_core_030;
  wire popcount25_gm8j_core_032;
  wire popcount25_gm8j_core_035;
  wire popcount25_gm8j_core_036;
  wire popcount25_gm8j_core_037;
  wire popcount25_gm8j_core_038;
  wire popcount25_gm8j_core_039;
  wire popcount25_gm8j_core_043;
  wire popcount25_gm8j_core_045;
  wire popcount25_gm8j_core_047;
  wire popcount25_gm8j_core_048;
  wire popcount25_gm8j_core_049;
  wire popcount25_gm8j_core_051;
  wire popcount25_gm8j_core_052;
  wire popcount25_gm8j_core_055;
  wire popcount25_gm8j_core_056;
  wire popcount25_gm8j_core_057;
  wire popcount25_gm8j_core_059;
  wire popcount25_gm8j_core_060;
  wire popcount25_gm8j_core_061;
  wire popcount25_gm8j_core_062;
  wire popcount25_gm8j_core_064;
  wire popcount25_gm8j_core_066;
  wire popcount25_gm8j_core_067;
  wire popcount25_gm8j_core_068;
  wire popcount25_gm8j_core_069;
  wire popcount25_gm8j_core_070;
  wire popcount25_gm8j_core_073;
  wire popcount25_gm8j_core_075;
  wire popcount25_gm8j_core_076;
  wire popcount25_gm8j_core_077;
  wire popcount25_gm8j_core_078;
  wire popcount25_gm8j_core_079;
  wire popcount25_gm8j_core_080;
  wire popcount25_gm8j_core_081;
  wire popcount25_gm8j_core_082;
  wire popcount25_gm8j_core_083;
  wire popcount25_gm8j_core_084;
  wire popcount25_gm8j_core_085;
  wire popcount25_gm8j_core_087;
  wire popcount25_gm8j_core_090;
  wire popcount25_gm8j_core_094;
  wire popcount25_gm8j_core_095;
  wire popcount25_gm8j_core_099;
  wire popcount25_gm8j_core_100;
  wire popcount25_gm8j_core_101;
  wire popcount25_gm8j_core_102;
  wire popcount25_gm8j_core_103;
  wire popcount25_gm8j_core_104;
  wire popcount25_gm8j_core_105;
  wire popcount25_gm8j_core_106;
  wire popcount25_gm8j_core_107;
  wire popcount25_gm8j_core_108;
  wire popcount25_gm8j_core_109;
  wire popcount25_gm8j_core_110;
  wire popcount25_gm8j_core_111;
  wire popcount25_gm8j_core_113;
  wire popcount25_gm8j_core_114;
  wire popcount25_gm8j_core_115;
  wire popcount25_gm8j_core_116;
  wire popcount25_gm8j_core_117;
  wire popcount25_gm8j_core_118;
  wire popcount25_gm8j_core_120;
  wire popcount25_gm8j_core_121;
  wire popcount25_gm8j_core_122;
  wire popcount25_gm8j_core_124;
  wire popcount25_gm8j_core_128;
  wire popcount25_gm8j_core_129;
  wire popcount25_gm8j_core_130;
  wire popcount25_gm8j_core_131;
  wire popcount25_gm8j_core_132;
  wire popcount25_gm8j_core_134;
  wire popcount25_gm8j_core_135;
  wire popcount25_gm8j_core_136;
  wire popcount25_gm8j_core_137;
  wire popcount25_gm8j_core_138;
  wire popcount25_gm8j_core_141;
  wire popcount25_gm8j_core_143;
  wire popcount25_gm8j_core_144;
  wire popcount25_gm8j_core_145_not;
  wire popcount25_gm8j_core_147;
  wire popcount25_gm8j_core_148;
  wire popcount25_gm8j_core_149;
  wire popcount25_gm8j_core_150;
  wire popcount25_gm8j_core_152;
  wire popcount25_gm8j_core_153;
  wire popcount25_gm8j_core_154;
  wire popcount25_gm8j_core_155;
  wire popcount25_gm8j_core_156;
  wire popcount25_gm8j_core_158;
  wire popcount25_gm8j_core_159;
  wire popcount25_gm8j_core_160;
  wire popcount25_gm8j_core_161;
  wire popcount25_gm8j_core_166;
  wire popcount25_gm8j_core_167;
  wire popcount25_gm8j_core_168;
  wire popcount25_gm8j_core_169;
  wire popcount25_gm8j_core_170;
  wire popcount25_gm8j_core_173;
  wire popcount25_gm8j_core_174;
  wire popcount25_gm8j_core_175;
  wire popcount25_gm8j_core_176;
  wire popcount25_gm8j_core_177;
  wire popcount25_gm8j_core_179;
  wire popcount25_gm8j_core_180;
  wire popcount25_gm8j_core_181;
  wire popcount25_gm8j_core_182;

  assign popcount25_gm8j_core_028 = input_a[1] | input_a[17];
  assign popcount25_gm8j_core_029 = ~(input_a[10] & input_a[20]);
  assign popcount25_gm8j_core_030 = ~input_a[8];
  assign popcount25_gm8j_core_032 = ~(input_a[7] & input_a[21]);
  assign popcount25_gm8j_core_035 = input_a[8] | input_a[11];
  assign popcount25_gm8j_core_036 = ~(input_a[22] & input_a[0]);
  assign popcount25_gm8j_core_037 = input_a[23] & input_a[8];
  assign popcount25_gm8j_core_038 = input_a[21] ^ input_a[17];
  assign popcount25_gm8j_core_039 = ~input_a[24];
  assign popcount25_gm8j_core_043 = ~(input_a[18] & input_a[9]);
  assign popcount25_gm8j_core_045 = ~input_a[0];
  assign popcount25_gm8j_core_047 = ~(input_a[4] ^ input_a[8]);
  assign popcount25_gm8j_core_048 = ~input_a[9];
  assign popcount25_gm8j_core_049 = ~(input_a[12] & input_a[15]);
  assign popcount25_gm8j_core_051 = input_a[19] & input_a[6];
  assign popcount25_gm8j_core_052 = input_a[23] & input_a[3];
  assign popcount25_gm8j_core_055 = input_a[22] | input_a[18];
  assign popcount25_gm8j_core_056 = ~(input_a[7] | input_a[3]);
  assign popcount25_gm8j_core_057 = input_a[5] ^ input_a[4];
  assign popcount25_gm8j_core_059 = input_a[10] | input_a[15];
  assign popcount25_gm8j_core_060 = input_a[20] | input_a[14];
  assign popcount25_gm8j_core_061 = ~input_a[11];
  assign popcount25_gm8j_core_062 = input_a[8] | input_a[1];
  assign popcount25_gm8j_core_064 = input_a[2] & input_a[18];
  assign popcount25_gm8j_core_066 = input_a[13] ^ input_a[11];
  assign popcount25_gm8j_core_067 = input_a[8] & input_a[4];
  assign popcount25_gm8j_core_068 = ~input_a[19];
  assign popcount25_gm8j_core_069 = ~(input_a[3] & input_a[2]);
  assign popcount25_gm8j_core_070 = input_a[13] | input_a[0];
  assign popcount25_gm8j_core_073 = ~(input_a[7] & input_a[10]);
  assign popcount25_gm8j_core_075 = ~(input_a[11] | input_a[21]);
  assign popcount25_gm8j_core_076 = input_a[16] & input_a[1];
  assign popcount25_gm8j_core_077 = ~(input_a[0] ^ input_a[5]);
  assign popcount25_gm8j_core_078 = input_a[24] | input_a[12];
  assign popcount25_gm8j_core_079 = ~input_a[10];
  assign popcount25_gm8j_core_080 = input_a[4] & input_a[13];
  assign popcount25_gm8j_core_081 = input_a[18] & input_a[1];
  assign popcount25_gm8j_core_082 = ~(input_a[4] & input_a[10]);
  assign popcount25_gm8j_core_083 = ~(input_a[20] & input_a[3]);
  assign popcount25_gm8j_core_084 = input_a[1] ^ input_a[0];
  assign popcount25_gm8j_core_085 = ~input_a[22];
  assign popcount25_gm8j_core_087 = ~input_a[23];
  assign popcount25_gm8j_core_090 = input_a[9] ^ input_a[21];
  assign popcount25_gm8j_core_094 = ~(input_a[0] | input_a[14]);
  assign popcount25_gm8j_core_095 = ~(input_a[22] | input_a[18]);
  assign popcount25_gm8j_core_099 = ~(input_a[6] ^ input_a[0]);
  assign popcount25_gm8j_core_100 = ~(input_a[7] | input_a[10]);
  assign popcount25_gm8j_core_101 = input_a[0] | input_a[10];
  assign popcount25_gm8j_core_102 = ~input_a[20];
  assign popcount25_gm8j_core_103 = ~(input_a[10] & input_a[17]);
  assign popcount25_gm8j_core_104 = ~input_a[11];
  assign popcount25_gm8j_core_105 = ~(input_a[2] ^ input_a[10]);
  assign popcount25_gm8j_core_106 = ~(input_a[18] ^ input_a[21]);
  assign popcount25_gm8j_core_107 = input_a[14] & input_a[4];
  assign popcount25_gm8j_core_108 = ~(input_a[4] ^ input_a[22]);
  assign popcount25_gm8j_core_109 = ~(input_a[19] ^ input_a[8]);
  assign popcount25_gm8j_core_110 = ~input_a[17];
  assign popcount25_gm8j_core_111 = input_a[9] & input_a[13];
  assign popcount25_gm8j_core_113 = input_a[2] | input_a[23];
  assign popcount25_gm8j_core_114 = ~(input_a[4] | input_a[17]);
  assign popcount25_gm8j_core_115 = ~(input_a[20] | input_a[7]);
  assign popcount25_gm8j_core_116 = input_a[8] & input_a[10];
  assign popcount25_gm8j_core_117 = ~(input_a[16] & input_a[10]);
  assign popcount25_gm8j_core_118 = input_a[19] | input_a[5];
  assign popcount25_gm8j_core_120 = ~(input_a[0] & input_a[2]);
  assign popcount25_gm8j_core_121 = ~(input_a[15] | input_a[21]);
  assign popcount25_gm8j_core_122 = input_a[19] & input_a[24];
  assign popcount25_gm8j_core_124 = input_a[24] | input_a[16];
  assign popcount25_gm8j_core_128 = ~input_a[4];
  assign popcount25_gm8j_core_129 = input_a[15] ^ input_a[20];
  assign popcount25_gm8j_core_130 = ~(input_a[7] ^ input_a[23]);
  assign popcount25_gm8j_core_131 = ~(input_a[24] | input_a[0]);
  assign popcount25_gm8j_core_132 = ~(input_a[22] | input_a[8]);
  assign popcount25_gm8j_core_134 = input_a[22] | input_a[3];
  assign popcount25_gm8j_core_135 = ~(input_a[21] & input_a[6]);
  assign popcount25_gm8j_core_136 = ~(input_a[0] & input_a[8]);
  assign popcount25_gm8j_core_137 = ~input_a[5];
  assign popcount25_gm8j_core_138 = input_a[4] & input_a[12];
  assign popcount25_gm8j_core_141 = ~(input_a[17] & input_a[9]);
  assign popcount25_gm8j_core_143 = input_a[20] | input_a[0];
  assign popcount25_gm8j_core_144 = ~(input_a[12] & input_a[8]);
  assign popcount25_gm8j_core_145_not = ~input_a[17];
  assign popcount25_gm8j_core_147 = ~(input_a[24] | input_a[7]);
  assign popcount25_gm8j_core_148 = ~(input_a[0] ^ input_a[20]);
  assign popcount25_gm8j_core_149 = ~(input_a[2] | input_a[22]);
  assign popcount25_gm8j_core_150 = input_a[17] & input_a[11];
  assign popcount25_gm8j_core_152 = input_a[14] ^ input_a[12];
  assign popcount25_gm8j_core_153 = ~input_a[12];
  assign popcount25_gm8j_core_154 = ~(input_a[9] & input_a[7]);
  assign popcount25_gm8j_core_155 = ~input_a[5];
  assign popcount25_gm8j_core_156 = input_a[10] & input_a[13];
  assign popcount25_gm8j_core_158 = ~(input_a[15] ^ input_a[9]);
  assign popcount25_gm8j_core_159 = input_a[3] ^ input_a[8];
  assign popcount25_gm8j_core_160 = input_a[21] & input_a[23];
  assign popcount25_gm8j_core_161 = ~(input_a[18] & input_a[23]);
  assign popcount25_gm8j_core_166 = ~(input_a[0] | input_a[5]);
  assign popcount25_gm8j_core_167 = input_a[4] | input_a[18];
  assign popcount25_gm8j_core_168 = input_a[1] ^ input_a[12];
  assign popcount25_gm8j_core_169 = input_a[22] ^ input_a[21];
  assign popcount25_gm8j_core_170 = input_a[0] & input_a[20];
  assign popcount25_gm8j_core_173 = input_a[15] & input_a[24];
  assign popcount25_gm8j_core_174 = input_a[9] ^ input_a[9];
  assign popcount25_gm8j_core_175 = ~(input_a[0] & input_a[3]);
  assign popcount25_gm8j_core_176 = ~input_a[10];
  assign popcount25_gm8j_core_177 = input_a[23] & input_a[2];
  assign popcount25_gm8j_core_179 = input_a[20] & input_a[9];
  assign popcount25_gm8j_core_180 = ~(input_a[14] | input_a[11]);
  assign popcount25_gm8j_core_181 = ~(input_a[18] & input_a[0]);
  assign popcount25_gm8j_core_182 = input_a[20] | input_a[24];

  assign popcount25_gm8j_out[0] = 1'b1;
  assign popcount25_gm8j_out[1] = input_a[10];
  assign popcount25_gm8j_out[2] = input_a[24];
  assign popcount25_gm8j_out[3] = 1'b1;
  assign popcount25_gm8j_out[4] = 1'b0;
endmodule