// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.73271
// WCE=18.0
// EP=0.935558%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_uob2(input [28:0] input_a, output [4:0] popcount29_uob2_out);
  wire popcount29_uob2_core_031;
  wire popcount29_uob2_core_032;
  wire popcount29_uob2_core_033;
  wire popcount29_uob2_core_038;
  wire popcount29_uob2_core_040;
  wire popcount29_uob2_core_041;
  wire popcount29_uob2_core_042;
  wire popcount29_uob2_core_048;
  wire popcount29_uob2_core_052;
  wire popcount29_uob2_core_053;
  wire popcount29_uob2_core_056;
  wire popcount29_uob2_core_057;
  wire popcount29_uob2_core_058;
  wire popcount29_uob2_core_059;
  wire popcount29_uob2_core_060;
  wire popcount29_uob2_core_061;
  wire popcount29_uob2_core_062;
  wire popcount29_uob2_core_064;
  wire popcount29_uob2_core_065;
  wire popcount29_uob2_core_066;
  wire popcount29_uob2_core_067;
  wire popcount29_uob2_core_068;
  wire popcount29_uob2_core_069;
  wire popcount29_uob2_core_071;
  wire popcount29_uob2_core_072;
  wire popcount29_uob2_core_073;
  wire popcount29_uob2_core_075;
  wire popcount29_uob2_core_076;
  wire popcount29_uob2_core_077;
  wire popcount29_uob2_core_079;
  wire popcount29_uob2_core_080;
  wire popcount29_uob2_core_081;
  wire popcount29_uob2_core_083;
  wire popcount29_uob2_core_084;
  wire popcount29_uob2_core_085;
  wire popcount29_uob2_core_086;
  wire popcount29_uob2_core_087;
  wire popcount29_uob2_core_092;
  wire popcount29_uob2_core_095;
  wire popcount29_uob2_core_096;
  wire popcount29_uob2_core_097;
  wire popcount29_uob2_core_098;
  wire popcount29_uob2_core_099;
  wire popcount29_uob2_core_100;
  wire popcount29_uob2_core_101;
  wire popcount29_uob2_core_102;
  wire popcount29_uob2_core_104;
  wire popcount29_uob2_core_105;
  wire popcount29_uob2_core_106;
  wire popcount29_uob2_core_107;
  wire popcount29_uob2_core_110;
  wire popcount29_uob2_core_111;
  wire popcount29_uob2_core_112;
  wire popcount29_uob2_core_113;
  wire popcount29_uob2_core_117;
  wire popcount29_uob2_core_118;
  wire popcount29_uob2_core_120;
  wire popcount29_uob2_core_123;
  wire popcount29_uob2_core_126;
  wire popcount29_uob2_core_127;
  wire popcount29_uob2_core_129;
  wire popcount29_uob2_core_130;
  wire popcount29_uob2_core_131;
  wire popcount29_uob2_core_132;
  wire popcount29_uob2_core_134;
  wire popcount29_uob2_core_138;
  wire popcount29_uob2_core_139;
  wire popcount29_uob2_core_143;
  wire popcount29_uob2_core_147;
  wire popcount29_uob2_core_148;
  wire popcount29_uob2_core_149;
  wire popcount29_uob2_core_151;
  wire popcount29_uob2_core_152;
  wire popcount29_uob2_core_153;
  wire popcount29_uob2_core_154;
  wire popcount29_uob2_core_156;
  wire popcount29_uob2_core_157;
  wire popcount29_uob2_core_158;
  wire popcount29_uob2_core_159;
  wire popcount29_uob2_core_160;
  wire popcount29_uob2_core_161;
  wire popcount29_uob2_core_162_not;
  wire popcount29_uob2_core_163;
  wire popcount29_uob2_core_164;
  wire popcount29_uob2_core_165;
  wire popcount29_uob2_core_166;
  wire popcount29_uob2_core_167;
  wire popcount29_uob2_core_168;
  wire popcount29_uob2_core_169;
  wire popcount29_uob2_core_171;
  wire popcount29_uob2_core_173;
  wire popcount29_uob2_core_174;
  wire popcount29_uob2_core_175;
  wire popcount29_uob2_core_176;
  wire popcount29_uob2_core_181;
  wire popcount29_uob2_core_183;
  wire popcount29_uob2_core_189;
  wire popcount29_uob2_core_191;
  wire popcount29_uob2_core_192;
  wire popcount29_uob2_core_194;
  wire popcount29_uob2_core_198;
  wire popcount29_uob2_core_201;
  wire popcount29_uob2_core_203;
  wire popcount29_uob2_core_205;
  wire popcount29_uob2_core_206;
  wire popcount29_uob2_core_207;

  assign popcount29_uob2_core_031 = input_a[24] | input_a[17];
  assign popcount29_uob2_core_032 = ~(input_a[24] & input_a[6]);
  assign popcount29_uob2_core_033 = ~(input_a[13] & input_a[13]);
  assign popcount29_uob2_core_038 = ~(input_a[4] ^ input_a[11]);
  assign popcount29_uob2_core_040 = ~input_a[9];
  assign popcount29_uob2_core_041 = ~input_a[15];
  assign popcount29_uob2_core_042 = input_a[8] & input_a[5];
  assign popcount29_uob2_core_048 = ~(input_a[20] & input_a[7]);
  assign popcount29_uob2_core_052 = input_a[15] ^ input_a[7];
  assign popcount29_uob2_core_053 = ~(input_a[13] | input_a[5]);
  assign popcount29_uob2_core_056 = input_a[27] & input_a[9];
  assign popcount29_uob2_core_057 = ~(input_a[24] ^ input_a[27]);
  assign popcount29_uob2_core_058 = ~(input_a[10] & input_a[28]);
  assign popcount29_uob2_core_059 = input_a[27] | input_a[2];
  assign popcount29_uob2_core_060 = ~input_a[22];
  assign popcount29_uob2_core_061 = ~(input_a[16] | input_a[1]);
  assign popcount29_uob2_core_062 = ~input_a[18];
  assign popcount29_uob2_core_064 = ~(input_a[26] | input_a[8]);
  assign popcount29_uob2_core_065 = input_a[7] | input_a[11];
  assign popcount29_uob2_core_066 = input_a[11] ^ input_a[0];
  assign popcount29_uob2_core_067 = ~input_a[2];
  assign popcount29_uob2_core_068 = ~(input_a[18] ^ input_a[14]);
  assign popcount29_uob2_core_069 = ~(input_a[10] | input_a[20]);
  assign popcount29_uob2_core_071 = ~(input_a[15] | input_a[21]);
  assign popcount29_uob2_core_072 = input_a[27] | input_a[21];
  assign popcount29_uob2_core_073 = ~(input_a[12] & input_a[26]);
  assign popcount29_uob2_core_075 = ~(input_a[1] ^ input_a[16]);
  assign popcount29_uob2_core_076 = ~(input_a[17] & input_a[11]);
  assign popcount29_uob2_core_077 = input_a[16] ^ input_a[10];
  assign popcount29_uob2_core_079 = ~input_a[16];
  assign popcount29_uob2_core_080 = input_a[10] & input_a[28];
  assign popcount29_uob2_core_081 = input_a[25] & input_a[12];
  assign popcount29_uob2_core_083 = ~(input_a[0] & input_a[12]);
  assign popcount29_uob2_core_084 = ~(input_a[28] | input_a[22]);
  assign popcount29_uob2_core_085 = input_a[3] ^ input_a[8];
  assign popcount29_uob2_core_086 = ~(input_a[7] & input_a[5]);
  assign popcount29_uob2_core_087 = input_a[7] & input_a[1];
  assign popcount29_uob2_core_092 = input_a[8] & input_a[4];
  assign popcount29_uob2_core_095 = ~(input_a[2] & input_a[4]);
  assign popcount29_uob2_core_096 = ~input_a[24];
  assign popcount29_uob2_core_097 = ~(input_a[9] & input_a[15]);
  assign popcount29_uob2_core_098 = ~input_a[20];
  assign popcount29_uob2_core_099 = input_a[27] | input_a[19];
  assign popcount29_uob2_core_100 = input_a[24] | input_a[21];
  assign popcount29_uob2_core_101 = ~(input_a[23] | input_a[4]);
  assign popcount29_uob2_core_102 = ~(input_a[14] & input_a[12]);
  assign popcount29_uob2_core_104 = input_a[12] ^ input_a[2];
  assign popcount29_uob2_core_105 = ~(input_a[21] & input_a[9]);
  assign popcount29_uob2_core_106 = ~(input_a[17] ^ input_a[19]);
  assign popcount29_uob2_core_107 = input_a[19] ^ input_a[4];
  assign popcount29_uob2_core_110 = ~(input_a[21] | input_a[7]);
  assign popcount29_uob2_core_111 = input_a[7] | input_a[6];
  assign popcount29_uob2_core_112 = ~input_a[26];
  assign popcount29_uob2_core_113 = input_a[17] | input_a[17];
  assign popcount29_uob2_core_117 = ~(input_a[18] & input_a[19]);
  assign popcount29_uob2_core_118 = ~(input_a[15] | input_a[16]);
  assign popcount29_uob2_core_120 = ~(input_a[26] | input_a[23]);
  assign popcount29_uob2_core_123 = ~input_a[9];
  assign popcount29_uob2_core_126 = ~(input_a[18] ^ input_a[1]);
  assign popcount29_uob2_core_127 = input_a[11] & input_a[14];
  assign popcount29_uob2_core_129 = input_a[3] & input_a[18];
  assign popcount29_uob2_core_130 = ~(input_a[21] ^ input_a[26]);
  assign popcount29_uob2_core_131 = ~(input_a[10] & input_a[15]);
  assign popcount29_uob2_core_132 = input_a[5] ^ input_a[21];
  assign popcount29_uob2_core_134 = input_a[21] & input_a[9];
  assign popcount29_uob2_core_138 = ~(input_a[7] | input_a[0]);
  assign popcount29_uob2_core_139 = input_a[18] | input_a[9];
  assign popcount29_uob2_core_143 = input_a[9] | input_a[4];
  assign popcount29_uob2_core_147 = ~(input_a[20] & input_a[8]);
  assign popcount29_uob2_core_148 = ~input_a[22];
  assign popcount29_uob2_core_149 = input_a[10] | input_a[15];
  assign popcount29_uob2_core_151 = ~(input_a[15] ^ input_a[27]);
  assign popcount29_uob2_core_152 = ~input_a[9];
  assign popcount29_uob2_core_153 = ~(input_a[11] ^ input_a[4]);
  assign popcount29_uob2_core_154 = input_a[1] | input_a[14];
  assign popcount29_uob2_core_156 = input_a[27] | input_a[4];
  assign popcount29_uob2_core_157 = input_a[7] | input_a[6];
  assign popcount29_uob2_core_158 = ~input_a[10];
  assign popcount29_uob2_core_159 = ~(input_a[7] | input_a[22]);
  assign popcount29_uob2_core_160 = input_a[26] ^ input_a[9];
  assign popcount29_uob2_core_161 = ~input_a[7];
  assign popcount29_uob2_core_162_not = ~input_a[9];
  assign popcount29_uob2_core_163 = input_a[21] ^ input_a[1];
  assign popcount29_uob2_core_164 = ~input_a[16];
  assign popcount29_uob2_core_165 = input_a[26] & input_a[22];
  assign popcount29_uob2_core_166 = input_a[6] ^ input_a[6];
  assign popcount29_uob2_core_167 = ~(input_a[27] | input_a[4]);
  assign popcount29_uob2_core_168 = ~(input_a[10] | input_a[13]);
  assign popcount29_uob2_core_169 = ~(input_a[14] ^ input_a[1]);
  assign popcount29_uob2_core_171 = ~input_a[23];
  assign popcount29_uob2_core_173 = input_a[17] ^ input_a[28];
  assign popcount29_uob2_core_174 = ~(input_a[22] | input_a[8]);
  assign popcount29_uob2_core_175 = ~(input_a[0] ^ input_a[11]);
  assign popcount29_uob2_core_176 = input_a[12] ^ input_a[8];
  assign popcount29_uob2_core_181 = input_a[20] ^ input_a[25];
  assign popcount29_uob2_core_183 = input_a[6] & input_a[21];
  assign popcount29_uob2_core_189 = ~(input_a[22] | input_a[15]);
  assign popcount29_uob2_core_191 = input_a[14] & input_a[27];
  assign popcount29_uob2_core_192 = input_a[8] & input_a[18];
  assign popcount29_uob2_core_194 = ~(input_a[6] ^ input_a[22]);
  assign popcount29_uob2_core_198 = input_a[7] | input_a[7];
  assign popcount29_uob2_core_201 = ~(input_a[21] ^ input_a[15]);
  assign popcount29_uob2_core_203 = input_a[11] | input_a[9];
  assign popcount29_uob2_core_205 = ~(input_a[18] & input_a[20]);
  assign popcount29_uob2_core_206 = ~(input_a[19] & input_a[6]);
  assign popcount29_uob2_core_207 = ~(input_a[4] ^ input_a[4]);

  assign popcount29_uob2_out[0] = 1'b1;
  assign popcount29_uob2_out[1] = input_a[5];
  assign popcount29_uob2_out[2] = 1'b0;
  assign popcount29_uob2_out[3] = 1'b0;
  assign popcount29_uob2_out[4] = 1'b1;
endmodule