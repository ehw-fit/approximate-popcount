
module cmp_pos(input [44:0] input_a, output [5:0] cgp_out);
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_054;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_081;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_114;
  wire cgp_core_117;
  wire cgp_core_118;
  wire cgp_core_121;
  wire cgp_core_122;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_130;
  wire cgp_core_131;
  wire cgp_core_132;
  wire cgp_core_133;
  wire cgp_core_134;
  wire cgp_core_136;
  wire cgp_core_137;
  wire cgp_core_139;
  wire cgp_core_140;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_145;
  wire cgp_core_147;
  wire cgp_core_149;
  wire cgp_core_150;
  wire cgp_core_151;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_159;
  wire cgp_core_167;
  wire cgp_core_168;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_181;
  wire cgp_core_185;
  wire cgp_core_191;
  wire cgp_core_194;
  wire cgp_core_195;
  wire cgp_core_196;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_206;
  wire cgp_core_207;
  wire cgp_core_208;
  wire cgp_core_209;
  wire cgp_core_210;
  wire cgp_core_211;
  wire cgp_core_213;
  wire cgp_core_216;
  wire cgp_core_220;
  wire cgp_core_221;
  wire cgp_core_224;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_231;
  wire cgp_core_234;
  wire cgp_core_240;
  wire cgp_core_241;
  wire cgp_core_249;
  wire cgp_core_250;
  wire cgp_core_252;
  wire cgp_core_253;
  wire cgp_core_254;
  wire cgp_core_255;
  wire cgp_core_257;
  wire cgp_core_258;
  wire cgp_core_259;
  wire cgp_core_260;
  wire cgp_core_263;
  wire cgp_core_265;
  wire cgp_core_266;
  wire cgp_core_267;
  wire cgp_core_268;
  wire cgp_core_269;
  wire cgp_core_271;
  wire cgp_core_275;
  wire cgp_core_277;
  wire cgp_core_278;
  wire cgp_core_281;
  wire cgp_core_282;
  wire cgp_core_283;
  wire cgp_core_284;
  wire cgp_core_286;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_290;
  wire cgp_core_291;
  wire cgp_core_292;
  wire cgp_core_293;
  wire cgp_core_294;
  wire cgp_core_295;
  wire cgp_core_298;
  wire cgp_core_299;
  wire cgp_core_300;
  wire cgp_core_301;
  wire cgp_core_302;
  wire cgp_core_303;
  wire cgp_core_305;
  wire cgp_core_306;
  wire cgp_core_309;
  wire cgp_core_310;
  wire cgp_core_312;
  wire cgp_core_316;
  wire cgp_core_318;
  wire cgp_core_319;
  wire cgp_core_320;
  wire cgp_core_321;
  wire cgp_core_323;
  wire cgp_core_324;
  wire cgp_core_326;
  wire cgp_core_327;
  wire cgp_core_328;
  wire cgp_core_329;
  wire cgp_core_330;
  wire cgp_core_332;
  wire cgp_core_333;
  wire cgp_core_336;
  wire cgp_core_337;
  wire cgp_core_338;
  wire cgp_core_342;
  wire cgp_core_344;
  wire cgp_core_345;
  wire cgp_core_346;
  wire cgp_core_347;
  wire cgp_core_348;
  wire cgp_core_349;
  wire cgp_core_350;
  wire cgp_core_351;
  wire cgp_core_352;
  wire cgp_core_353;
  wire cgp_core_354;
  wire cgp_core_355;
  wire cgp_core_356;

  assign cgp_core_047 = input_a[13] | input_a[31];
  assign cgp_core_048 = ~(input_a[11] ^ input_a[34]);
  assign cgp_core_049 = input_a[8] ^ input_a[41];
  assign cgp_core_050 = ~input_a[22];
  assign cgp_core_051 = input_a[1] ^ input_a[16];
  assign cgp_core_052 = input_a[25] | input_a[10];
  assign cgp_core_054 = input_a[37] | input_a[18];
  assign cgp_core_056 = input_a[1] | input_a[31];
  assign cgp_core_057 = input_a[12] ^ input_a[18];
  assign cgp_core_058 = input_a[22] ^ input_a[32];
  assign cgp_core_059 = input_a[36] ^ input_a[44];
  assign cgp_core_060 = ~(input_a[42] | input_a[13]);
  assign cgp_core_061 = input_a[11] ^ input_a[37];
  assign cgp_core_062 = ~(input_a[41] ^ input_a[31]);
  assign cgp_core_063 = ~(input_a[35] ^ input_a[14]);
  assign cgp_core_068 = ~(input_a[29] & input_a[22]);
  assign cgp_core_069 = input_a[27] ^ input_a[25];
  assign cgp_core_070 = input_a[35] & input_a[26];
  assign cgp_core_072 = input_a[33] ^ input_a[40];
  assign cgp_core_073 = input_a[36] ^ input_a[44];
  assign cgp_core_074 = ~(input_a[32] ^ input_a[31]);
  assign cgp_core_075 = ~input_a[25];
  assign cgp_core_076 = input_a[21] & input_a[11];
  assign cgp_core_077 = input_a[20] & input_a[26];
  assign cgp_core_079 = ~(input_a[36] & input_a[6]);
  assign cgp_core_081 = ~(input_a[12] & input_a[20]);
  assign cgp_core_084 = ~(input_a[17] | input_a[3]);
  assign cgp_core_086 = input_a[19] ^ input_a[3];
  assign cgp_core_087 = ~(input_a[11] ^ input_a[12]);
  assign cgp_core_089 = ~(input_a[39] | input_a[24]);
  assign cgp_core_090 = ~(input_a[2] & input_a[4]);
  assign cgp_core_093 = input_a[37] & input_a[40];
  assign cgp_core_094 = ~input_a[22];
  assign cgp_core_095 = ~(input_a[38] | input_a[20]);
  assign cgp_core_099 = ~(input_a[14] | input_a[33]);
  assign cgp_core_100 = ~(input_a[15] & input_a[39]);
  assign cgp_core_101 = input_a[31] & input_a[19];
  assign cgp_core_104 = ~input_a[28];
  assign cgp_core_105 = ~(input_a[27] ^ input_a[35]);
  assign cgp_core_106 = input_a[5] & input_a[41];
  assign cgp_core_107 = ~(input_a[3] | input_a[4]);
  assign cgp_core_109 = ~(input_a[21] & input_a[43]);
  assign cgp_core_110 = ~(input_a[32] | input_a[24]);
  assign cgp_core_114 = input_a[20] & input_a[8];
  assign cgp_core_117 = ~(input_a[43] | input_a[24]);
  assign cgp_core_118 = cgp_core_106 & cgp_core_114;
  assign cgp_core_121 = input_a[0] | input_a[36];
  assign cgp_core_122 = ~input_a[4];
  assign cgp_core_123 = ~(input_a[14] ^ input_a[13]);
  assign cgp_core_124 = input_a[34] | input_a[19];
  assign cgp_core_125 = ~(input_a[32] & input_a[16]);
  assign cgp_core_126 = ~(input_a[12] & input_a[28]);
  assign cgp_core_127 = input_a[43] & input_a[34];
  assign cgp_core_128 = ~(input_a[42] ^ input_a[20]);
  assign cgp_core_130 = ~(input_a[10] & input_a[35]);
  assign cgp_core_131 = ~(input_a[14] | input_a[19]);
  assign cgp_core_132 = input_a[16] & input_a[42];
  assign cgp_core_133 = input_a[26] ^ input_a[21];
  assign cgp_core_134 = input_a[40] | input_a[13];
  assign cgp_core_136 = ~input_a[44];
  assign cgp_core_137 = ~input_a[11];
  assign cgp_core_139 = ~(input_a[22] & input_a[37]);
  assign cgp_core_140 = input_a[12] ^ input_a[10];
  assign cgp_core_141 = ~(input_a[1] ^ input_a[19]);
  assign cgp_core_142 = ~(input_a[38] | input_a[44]);
  assign cgp_core_143 = input_a[11] | input_a[26];
  assign cgp_core_145 = input_a[36] | input_a[34];
  assign cgp_core_147 = input_a[38] & input_a[41];
  assign cgp_core_149 = input_a[15] & cgp_core_136;
  assign cgp_core_150 = ~(input_a[10] ^ input_a[12]);
  assign cgp_core_151 = input_a[18] ^ input_a[21];
  assign cgp_core_153 = cgp_core_118 ^ cgp_core_143;
  assign cgp_core_154 = cgp_core_118 & cgp_core_143;
  assign cgp_core_155 = cgp_core_153 ^ cgp_core_149;
  assign cgp_core_156 = cgp_core_153 & cgp_core_149;
  assign cgp_core_157 = cgp_core_154 | cgp_core_156;
  assign cgp_core_159 = ~(input_a[35] & input_a[26]);
  assign cgp_core_167 = input_a[0] | input_a[7];
  assign cgp_core_168 = input_a[10] & input_a[1];
  assign cgp_core_170 = input_a[44] ^ cgp_core_155;
  assign cgp_core_171 = input_a[44] & cgp_core_155;
  assign cgp_core_172 = cgp_core_170 ^ cgp_core_168;
  assign cgp_core_173 = cgp_core_170 & cgp_core_168;
  assign cgp_core_174 = cgp_core_171 | cgp_core_173;
  assign cgp_core_177 = cgp_core_157 ^ cgp_core_174;
  assign cgp_core_178 = cgp_core_157 & cgp_core_174;
  assign cgp_core_181 = ~(input_a[44] | input_a[0]);
  assign cgp_core_185 = ~(input_a[12] ^ input_a[42]);
  assign cgp_core_191 = ~input_a[5];
  assign cgp_core_194 = ~(input_a[6] | input_a[0]);
  assign cgp_core_195 = ~(input_a[12] | input_a[35]);
  assign cgp_core_196 = input_a[12] ^ input_a[41];
  assign cgp_core_200 = input_a[39] & input_a[3];
  assign cgp_core_201 = ~(input_a[14] & input_a[1]);
  assign cgp_core_202 = ~(input_a[20] ^ input_a[9]);
  assign cgp_core_206 = ~input_a[37];
  assign cgp_core_207 = ~(input_a[26] | input_a[13]);
  assign cgp_core_208 = ~(input_a[37] | input_a[17]);
  assign cgp_core_209 = input_a[14] | input_a[44];
  assign cgp_core_210 = input_a[12] & input_a[7];
  assign cgp_core_211 = ~(input_a[34] & input_a[24]);
  assign cgp_core_213 = input_a[22] | input_a[41];
  assign cgp_core_216 = ~(input_a[10] & input_a[19]);
  assign cgp_core_220 = ~(input_a[7] & input_a[18]);
  assign cgp_core_221 = ~(input_a[23] & input_a[39]);
  assign cgp_core_224 = ~(input_a[35] & input_a[15]);
  assign cgp_core_228 = input_a[6] & input_a[5];
  assign cgp_core_229 = ~(input_a[8] & input_a[31]);
  assign cgp_core_231 = ~(input_a[30] | input_a[43]);
  assign cgp_core_234 = ~input_a[14];
  assign cgp_core_240 = ~(input_a[20] & input_a[12]);
  assign cgp_core_241 = ~(input_a[13] ^ input_a[25]);
  assign cgp_core_249 = ~input_a[23];
  assign cgp_core_250 = ~(input_a[10] ^ input_a[30]);
  assign cgp_core_252 = ~(input_a[34] | input_a[9]);
  assign cgp_core_253 = ~(input_a[43] | input_a[3]);
  assign cgp_core_254 = ~(input_a[21] & input_a[43]);
  assign cgp_core_255 = ~(input_a[32] & input_a[33]);
  assign cgp_core_257 = ~(input_a[34] | input_a[27]);
  assign cgp_core_258 = ~(input_a[20] & input_a[15]);
  assign cgp_core_259 = ~(input_a[35] | input_a[41]);
  assign cgp_core_260 = input_a[15] | input_a[42];
  assign cgp_core_263 = ~(input_a[27] & input_a[2]);
  assign cgp_core_265 = ~input_a[24];
  assign cgp_core_266 = input_a[2] & input_a[41];
  assign cgp_core_267 = ~input_a[13];
  assign cgp_core_268 = input_a[24] | input_a[43];
  assign cgp_core_269 = ~input_a[43];
  assign cgp_core_271 = input_a[33] & input_a[6];
  assign cgp_core_275 = input_a[11] ^ input_a[21];
  assign cgp_core_277 = ~(input_a[20] | input_a[17]);
  assign cgp_core_278 = ~(input_a[35] | input_a[17]);
  assign cgp_core_281 = ~input_a[14];
  assign cgp_core_282 = input_a[27] ^ input_a[23];
  assign cgp_core_283 = ~input_a[2];
  assign cgp_core_284 = ~input_a[30];
  assign cgp_core_286 = ~input_a[21];
  assign cgp_core_287 = ~input_a[17];
  assign cgp_core_288 = ~input_a[8];
  assign cgp_core_289 = ~(input_a[2] ^ input_a[23]);
  assign cgp_core_290 = ~(input_a[15] & input_a[25]);
  assign cgp_core_291 = ~input_a[15];
  assign cgp_core_292 = ~(input_a[2] & input_a[1]);
  assign cgp_core_293 = ~(input_a[35] ^ input_a[1]);
  assign cgp_core_294 = ~(input_a[40] ^ input_a[30]);
  assign cgp_core_295 = input_a[11] | input_a[13];
  assign cgp_core_298 = ~input_a[39];
  assign cgp_core_299 = ~(input_a[1] | input_a[30]);
  assign cgp_core_300 = ~input_a[35];
  assign cgp_core_301 = ~(input_a[0] ^ input_a[24]);
  assign cgp_core_302 = ~(input_a[11] | input_a[10]);
  assign cgp_core_303 = ~(input_a[32] & input_a[37]);
  assign cgp_core_305 = input_a[1] | input_a[20];
  assign cgp_core_306 = ~input_a[26];
  assign cgp_core_309 = input_a[35] ^ input_a[17];
  assign cgp_core_310 = input_a[27] ^ input_a[7];
  assign cgp_core_312 = input_a[33] & input_a[30];
  assign cgp_core_316 = ~input_a[29];
  assign cgp_core_318 = input_a[5] & input_a[2];
  assign cgp_core_319 = ~(input_a[28] & input_a[43]);
  assign cgp_core_320 = ~input_a[35];
  assign cgp_core_321 = input_a[31] & input_a[0];
  assign cgp_core_323 = ~input_a[40];
  assign cgp_core_324 = ~(input_a[23] & input_a[33]);
  assign cgp_core_326 = input_a[1] ^ input_a[6];
  assign cgp_core_327 = ~input_a[4];
  assign cgp_core_328 = input_a[33] & input_a[40];
  assign cgp_core_329 = input_a[41] | input_a[27];
  assign cgp_core_330 = ~(input_a[3] | input_a[37]);
  assign cgp_core_332 = input_a[38] ^ input_a[39];
  assign cgp_core_333 = input_a[13] | input_a[26];
  assign cgp_core_336 = input_a[4] & input_a[12];
  assign cgp_core_337 = cgp_core_172 ^ cgp_core_300;
  assign cgp_core_338 = cgp_core_172 & cgp_core_300;
  assign cgp_core_342 = cgp_core_177 ^ cgp_core_320;
  assign cgp_core_344 = cgp_core_342 ^ cgp_core_338;
  assign cgp_core_345 = cgp_core_342 & cgp_core_338;
  assign cgp_core_346 = cgp_core_177 | cgp_core_345;
  assign cgp_core_347 = cgp_core_178 ^ input_a[35];
  assign cgp_core_348 = cgp_core_178 & input_a[35];
  assign cgp_core_349 = cgp_core_347 | cgp_core_346;
  assign cgp_core_350 = input_a[27] | input_a[14];
  assign cgp_core_351 = ~input_a[26];
  assign cgp_core_352 = ~(input_a[37] & input_a[20]);
  assign cgp_core_353 = ~(input_a[5] & input_a[12]);
  assign cgp_core_354 = ~(input_a[42] | input_a[35]);
  assign cgp_core_355 = ~(input_a[8] ^ input_a[15]);
  assign cgp_core_356 = ~(input_a[13] | input_a[13]);

  assign cgp_out[0] = input_a[23];
  assign cgp_out[1] = cgp_core_300;
  assign cgp_out[2] = cgp_core_337;
  assign cgp_out[3] = cgp_core_344;
  assign cgp_out[4] = cgp_core_349;
  assign cgp_out[5] = cgp_core_348;
endmodule

module cmp_neg(input [38:0] input_a, output [5:0] cgp_out);
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_111;
  wire cgp_core_113;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_119;
  wire cgp_core_121;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_133;
  wire cgp_core_134;
  wire cgp_core_136;
  wire cgp_core_138;
  wire cgp_core_140;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_158;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_162;
  wire cgp_core_164;
  wire cgp_core_166;
  wire cgp_core_167;
  wire cgp_core_168;
  wire cgp_core_169;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_189;
  wire cgp_core_190;
  wire cgp_core_193;
  wire cgp_core_197;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_203;
  wire cgp_core_210;
  wire cgp_core_212;
  wire cgp_core_213;
  wire cgp_core_216;
  wire cgp_core_217;
  wire cgp_core_222;
  wire cgp_core_225;
  wire cgp_core_226;
  wire cgp_core_227;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_230;
  wire cgp_core_232;
  wire cgp_core_233;
  wire cgp_core_235;
  wire cgp_core_237;
  wire cgp_core_238;
  wire cgp_core_239;
  wire cgp_core_240;
  wire cgp_core_243;
  wire cgp_core_244;
  wire cgp_core_246;
  wire cgp_core_247;
  wire cgp_core_252;
  wire cgp_core_255;
  wire cgp_core_256;
  wire cgp_core_258;
  wire cgp_core_259;
  wire cgp_core_262;
  wire cgp_core_265;
  wire cgp_core_267;
  wire cgp_core_268;
  wire cgp_core_271;
  wire cgp_core_272;
  wire cgp_core_276;
  wire cgp_core_278;
  wire cgp_core_279;
  wire cgp_core_280;
  wire cgp_core_282;
  wire cgp_core_283;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_290;
  wire cgp_core_291;
  wire cgp_core_292;
  wire cgp_core_293;
  wire cgp_core_294;
  wire cgp_core_295;
  wire cgp_core_296;
  wire cgp_core_298;
  wire cgp_core_299;
  wire cgp_core_302;
  wire cgp_core_303;
  wire cgp_core_305;
  wire cgp_core_306;

  assign cgp_core_041 = input_a[0] ^ input_a[1];
  assign cgp_core_042 = input_a[0] & input_a[1];
  assign cgp_core_043 = ~(input_a[2] & input_a[3]);
  assign cgp_core_044 = input_a[2] & input_a[3];
  assign cgp_core_045 = ~(input_a[23] ^ input_a[1]);
  assign cgp_core_046 = input_a[37] & cgp_core_043;
  assign cgp_core_047 = cgp_core_042 ^ cgp_core_044;
  assign cgp_core_048 = cgp_core_042 & cgp_core_044;
  assign cgp_core_049 = cgp_core_047 | cgp_core_046;
  assign cgp_core_052 = ~(input_a[22] | input_a[35]);
  assign cgp_core_053 = ~(input_a[19] ^ input_a[3]);
  assign cgp_core_055 = ~(input_a[16] & input_a[7]);
  assign cgp_core_057 = input_a[7] ^ input_a[16];
  assign cgp_core_060 = ~input_a[30];
  assign cgp_core_062 = input_a[16] | input_a[30];
  assign cgp_core_066 = ~input_a[2];
  assign cgp_core_068 = input_a[26] ^ input_a[31];
  assign cgp_core_069 = ~(input_a[22] ^ input_a[3]);
  assign cgp_core_071 = cgp_core_049 ^ cgp_core_062;
  assign cgp_core_072 = cgp_core_049 & cgp_core_062;
  assign cgp_core_074 = input_a[21] & input_a[10];
  assign cgp_core_077 = ~(input_a[15] | input_a[20]);
  assign cgp_core_078 = cgp_core_048 | cgp_core_072;
  assign cgp_core_079 = ~input_a[8];
  assign cgp_core_080 = ~(input_a[28] & input_a[32]);
  assign cgp_core_082 = input_a[20] ^ input_a[38];
  assign cgp_core_084 = input_a[5] & input_a[4];
  assign cgp_core_085 = input_a[12] ^ input_a[13];
  assign cgp_core_086 = input_a[12] & input_a[13];
  assign cgp_core_087 = ~(input_a[38] | input_a[36]);
  assign cgp_core_088 = input_a[11] & cgp_core_085;
  assign cgp_core_089 = cgp_core_086 | cgp_core_088;
  assign cgp_core_092 = input_a[32] & input_a[23];
  assign cgp_core_093 = cgp_core_084 ^ cgp_core_089;
  assign cgp_core_094 = cgp_core_084 & cgp_core_089;
  assign cgp_core_095 = cgp_core_093 ^ cgp_core_092;
  assign cgp_core_096 = cgp_core_093 & cgp_core_092;
  assign cgp_core_097 = cgp_core_094 | cgp_core_096;
  assign cgp_core_099 = ~input_a[35];
  assign cgp_core_101 = input_a[20] & input_a[15];
  assign cgp_core_102 = input_a[17] ^ input_a[18];
  assign cgp_core_103 = input_a[17] & input_a[18];
  assign cgp_core_104 = ~(input_a[31] | input_a[15]);
  assign cgp_core_105 = input_a[33] & cgp_core_102;
  assign cgp_core_106 = cgp_core_103 | cgp_core_105;
  assign cgp_core_109 = input_a[4] ^ input_a[34];
  assign cgp_core_110 = cgp_core_101 ^ cgp_core_106;
  assign cgp_core_111 = cgp_core_101 & cgp_core_106;
  assign cgp_core_113 = ~(input_a[4] & input_a[12]);
  assign cgp_core_116 = input_a[19] & input_a[8];
  assign cgp_core_117 = ~input_a[4];
  assign cgp_core_119 = cgp_core_095 ^ cgp_core_110;
  assign cgp_core_121 = ~cgp_core_119;
  assign cgp_core_123 = cgp_core_095 | cgp_core_119;
  assign cgp_core_124 = cgp_core_097 ^ cgp_core_111;
  assign cgp_core_125 = cgp_core_097 & cgp_core_111;
  assign cgp_core_126 = cgp_core_124 ^ cgp_core_123;
  assign cgp_core_127 = cgp_core_124 & cgp_core_123;
  assign cgp_core_128 = cgp_core_125 | cgp_core_127;
  assign cgp_core_133 = ~input_a[5];
  assign cgp_core_134 = ~input_a[5];
  assign cgp_core_136 = cgp_core_071 ^ cgp_core_121;
  assign cgp_core_138 = ~cgp_core_136;
  assign cgp_core_140 = cgp_core_071 | cgp_core_136;
  assign cgp_core_141 = cgp_core_078 ^ cgp_core_126;
  assign cgp_core_142 = cgp_core_078 & cgp_core_126;
  assign cgp_core_143 = cgp_core_141 ^ cgp_core_140;
  assign cgp_core_144 = cgp_core_141 & cgp_core_140;
  assign cgp_core_145 = cgp_core_142 | cgp_core_144;
  assign cgp_core_148 = cgp_core_128 ^ cgp_core_145;
  assign cgp_core_149 = cgp_core_128 & cgp_core_145;
  assign cgp_core_154 = ~(input_a[9] | input_a[25]);
  assign cgp_core_155 = input_a[5] ^ input_a[10];
  assign cgp_core_156 = input_a[19] ^ input_a[36];
  assign cgp_core_157 = input_a[19] & input_a[8];
  assign cgp_core_158 = input_a[17] ^ input_a[10];
  assign cgp_core_159 = input_a[31] & input_a[9];
  assign cgp_core_160 = ~(input_a[2] | input_a[38]);
  assign cgp_core_162 = cgp_core_159 | input_a[35];
  assign cgp_core_164 = ~input_a[7];
  assign cgp_core_166 = cgp_core_157 ^ cgp_core_162;
  assign cgp_core_167 = cgp_core_157 & input_a[35];
  assign cgp_core_168 = cgp_core_166 ^ input_a[14];
  assign cgp_core_169 = cgp_core_166 & input_a[14];
  assign cgp_core_170 = cgp_core_167 | cgp_core_169;
  assign cgp_core_171 = cgp_core_159 | cgp_core_170;
  assign cgp_core_172 = input_a[30] ^ input_a[34];
  assign cgp_core_173 = input_a[24] ^ input_a[25];
  assign cgp_core_174 = input_a[24] & input_a[25];
  assign cgp_core_175 = input_a[27] ^ input_a[28];
  assign cgp_core_176 = input_a[27] & input_a[28];
  assign cgp_core_177 = input_a[26] ^ cgp_core_175;
  assign cgp_core_178 = input_a[26] & cgp_core_175;
  assign cgp_core_179 = cgp_core_176 | cgp_core_178;
  assign cgp_core_182 = cgp_core_173 & cgp_core_177;
  assign cgp_core_183 = cgp_core_174 ^ cgp_core_179;
  assign cgp_core_184 = cgp_core_174 & cgp_core_179;
  assign cgp_core_185 = cgp_core_183 ^ cgp_core_182;
  assign cgp_core_186 = cgp_core_183 & cgp_core_182;
  assign cgp_core_187 = cgp_core_184 | cgp_core_186;
  assign cgp_core_189 = input_a[10] | input_a[1];
  assign cgp_core_190 = input_a[13] ^ input_a[3];
  assign cgp_core_193 = cgp_core_168 & cgp_core_185;
  assign cgp_core_197 = cgp_core_171 ^ cgp_core_187;
  assign cgp_core_199 = cgp_core_197 | cgp_core_193;
  assign cgp_core_200 = input_a[34] & cgp_core_193;
  assign cgp_core_201 = cgp_core_171 | cgp_core_200;
  assign cgp_core_203 = ~input_a[34];
  assign cgp_core_210 = ~(input_a[4] ^ input_a[35]);
  assign cgp_core_212 = input_a[36] | input_a[20];
  assign cgp_core_213 = input_a[38] ^ input_a[37];
  assign cgp_core_216 = ~(input_a[2] ^ input_a[0]);
  assign cgp_core_217 = input_a[18] ^ input_a[18];
  assign cgp_core_222 = input_a[3] | input_a[6];
  assign cgp_core_225 = input_a[38] & input_a[22];
  assign cgp_core_226 = ~(input_a[1] & input_a[36]);
  assign cgp_core_227 = ~(input_a[33] ^ input_a[4]);
  assign cgp_core_228 = input_a[34] ^ input_a[14];
  assign cgp_core_229 = input_a[37] | input_a[13];
  assign cgp_core_230 = ~(input_a[16] | input_a[31]);
  assign cgp_core_232 = ~(input_a[33] | input_a[12]);
  assign cgp_core_233 = input_a[4] | input_a[21];
  assign cgp_core_235 = ~input_a[15];
  assign cgp_core_237 = ~(input_a[19] & input_a[19]);
  assign cgp_core_238 = input_a[33] ^ input_a[38];
  assign cgp_core_239 = ~input_a[38];
  assign cgp_core_240 = ~(input_a[12] ^ input_a[3]);
  assign cgp_core_243 = ~cgp_core_225;
  assign cgp_core_244 = input_a[4] & cgp_core_225;
  assign cgp_core_246 = ~cgp_core_243;
  assign cgp_core_247 = cgp_core_244 | cgp_core_246;
  assign cgp_core_252 = input_a[37] ^ input_a[21];
  assign cgp_core_255 = ~(input_a[30] & input_a[7]);
  assign cgp_core_256 = ~(input_a[5] ^ input_a[7]);
  assign cgp_core_258 = input_a[20] & input_a[22];
  assign cgp_core_259 = input_a[8] & input_a[10];
  assign cgp_core_262 = ~cgp_core_243;
  assign cgp_core_265 = cgp_core_199 ^ cgp_core_247;
  assign cgp_core_267 = cgp_core_265 ^ cgp_core_243;
  assign cgp_core_268 = input_a[20] & input_a[14];
  assign cgp_core_271 = ~(input_a[0] | input_a[37]);
  assign cgp_core_272 = cgp_core_201 | cgp_core_199;
  assign cgp_core_276 = input_a[15] & input_a[6];
  assign cgp_core_278 = ~(input_a[22] ^ input_a[17]);
  assign cgp_core_279 = ~input_a[0];
  assign cgp_core_280 = input_a[27] & input_a[18];
  assign cgp_core_282 = cgp_core_138 ^ cgp_core_262;
  assign cgp_core_283 = cgp_core_138 & cgp_core_262;
  assign cgp_core_287 = cgp_core_143 ^ cgp_core_267;
  assign cgp_core_288 = cgp_core_143 & cgp_core_267;
  assign cgp_core_289 = cgp_core_287 ^ cgp_core_283;
  assign cgp_core_290 = cgp_core_287 & cgp_core_283;
  assign cgp_core_291 = cgp_core_288 | cgp_core_290;
  assign cgp_core_292 = cgp_core_148 ^ cgp_core_272;
  assign cgp_core_293 = cgp_core_148 & cgp_core_272;
  assign cgp_core_294 = cgp_core_292 ^ cgp_core_291;
  assign cgp_core_295 = cgp_core_292 & cgp_core_291;
  assign cgp_core_296 = cgp_core_293 | cgp_core_295;
  assign cgp_core_298 = input_a[10] & input_a[27];
  assign cgp_core_299 = cgp_core_149 ^ cgp_core_296;
  assign cgp_core_302 = ~(input_a[35] ^ input_a[1]);
  assign cgp_core_303 = ~(input_a[30] ^ input_a[35]);
  assign cgp_core_305 = input_a[30] & input_a[15];
  assign cgp_core_306 = input_a[23] ^ input_a[17];

  assign cgp_out[0] = input_a[34];
  assign cgp_out[1] = cgp_core_282;
  assign cgp_out[2] = cgp_core_289;
  assign cgp_out[3] = cgp_core_294;
  assign cgp_out[4] = cgp_core_299;
  assign cgp_out[5] = 1'b0;
endmodule
module pcc(input [44:0] pos, input [38:0] neg, output outval);
    wire [5:0] cnt_pos;
    wire [5:0] cnt_neg;

    cmp_pos ipos(pos, cnt_pos);
    cmp_neg ineg(neg, cnt_neg);

    assign outval = (cnt_pos >= cnt_neg);
endmodule
