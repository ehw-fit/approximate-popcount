// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.31641
// WCE=15.0
// EP=0.865499%
// Printed PDK parameters:
//  Area=476280.0
//  Delay=2551099.0
//  Power=3460.8

module popcount30_uea4(input [29:0] input_a, output [4:0] popcount30_uea4_out);
  wire popcount30_uea4_core_032;
  wire popcount30_uea4_core_033;
  wire popcount30_uea4_core_038;
  wire popcount30_uea4_core_041;
  wire popcount30_uea4_core_043;
  wire popcount30_uea4_core_044;
  wire popcount30_uea4_core_045;
  wire popcount30_uea4_core_046;
  wire popcount30_uea4_core_048;
  wire popcount30_uea4_core_049;
  wire popcount30_uea4_core_050;
  wire popcount30_uea4_core_053;
  wire popcount30_uea4_core_054;
  wire popcount30_uea4_core_055;
  wire popcount30_uea4_core_056;
  wire popcount30_uea4_core_057;
  wire popcount30_uea4_core_060;
  wire popcount30_uea4_core_061;
  wire popcount30_uea4_core_062;
  wire popcount30_uea4_core_063;
  wire popcount30_uea4_core_066;
  wire popcount30_uea4_core_067;
  wire popcount30_uea4_core_068;
  wire popcount30_uea4_core_069;
  wire popcount30_uea4_core_070;
  wire popcount30_uea4_core_071;
  wire popcount30_uea4_core_072;
  wire popcount30_uea4_core_073;
  wire popcount30_uea4_core_074;
  wire popcount30_uea4_core_075;
  wire popcount30_uea4_core_078;
  wire popcount30_uea4_core_079;
  wire popcount30_uea4_core_081;
  wire popcount30_uea4_core_083;
  wire popcount30_uea4_core_084;
  wire popcount30_uea4_core_085;
  wire popcount30_uea4_core_086;
  wire popcount30_uea4_core_087;
  wire popcount30_uea4_core_091;
  wire popcount30_uea4_core_092;
  wire popcount30_uea4_core_093_not;
  wire popcount30_uea4_core_094;
  wire popcount30_uea4_core_096;
  wire popcount30_uea4_core_097;
  wire popcount30_uea4_core_098;
  wire popcount30_uea4_core_101;
  wire popcount30_uea4_core_102;
  wire popcount30_uea4_core_103;
  wire popcount30_uea4_core_105;
  wire popcount30_uea4_core_106;
  wire popcount30_uea4_core_107;
  wire popcount30_uea4_core_108;
  wire popcount30_uea4_core_109;
  wire popcount30_uea4_core_110;
  wire popcount30_uea4_core_112;
  wire popcount30_uea4_core_113;
  wire popcount30_uea4_core_114;
  wire popcount30_uea4_core_116;
  wire popcount30_uea4_core_117;
  wire popcount30_uea4_core_118;
  wire popcount30_uea4_core_119;
  wire popcount30_uea4_core_120;
  wire popcount30_uea4_core_121;
  wire popcount30_uea4_core_123;
  wire popcount30_uea4_core_126;
  wire popcount30_uea4_core_127;
  wire popcount30_uea4_core_128;
  wire popcount30_uea4_core_129;
  wire popcount30_uea4_core_131;
  wire popcount30_uea4_core_132;
  wire popcount30_uea4_core_133;
  wire popcount30_uea4_core_135;
  wire popcount30_uea4_core_137;
  wire popcount30_uea4_core_138;
  wire popcount30_uea4_core_140;
  wire popcount30_uea4_core_143;
  wire popcount30_uea4_core_145;
  wire popcount30_uea4_core_146;
  wire popcount30_uea4_core_147;
  wire popcount30_uea4_core_148;
  wire popcount30_uea4_core_149;
  wire popcount30_uea4_core_151;
  wire popcount30_uea4_core_155;
  wire popcount30_uea4_core_157;
  wire popcount30_uea4_core_158;
  wire popcount30_uea4_core_159;
  wire popcount30_uea4_core_160;
  wire popcount30_uea4_core_161;
  wire popcount30_uea4_core_162;
  wire popcount30_uea4_core_163;
  wire popcount30_uea4_core_164;
  wire popcount30_uea4_core_165;
  wire popcount30_uea4_core_166;
  wire popcount30_uea4_core_167;
  wire popcount30_uea4_core_168;
  wire popcount30_uea4_core_169;
  wire popcount30_uea4_core_171;
  wire popcount30_uea4_core_173;
  wire popcount30_uea4_core_174;
  wire popcount30_uea4_core_175;
  wire popcount30_uea4_core_177;
  wire popcount30_uea4_core_178;
  wire popcount30_uea4_core_179;
  wire popcount30_uea4_core_180;
  wire popcount30_uea4_core_181;
  wire popcount30_uea4_core_182;
  wire popcount30_uea4_core_183;
  wire popcount30_uea4_core_186;
  wire popcount30_uea4_core_187;
  wire popcount30_uea4_core_194;
  wire popcount30_uea4_core_196;
  wire popcount30_uea4_core_197;
  wire popcount30_uea4_core_198;
  wire popcount30_uea4_core_199;
  wire popcount30_uea4_core_200;
  wire popcount30_uea4_core_201;
  wire popcount30_uea4_core_202;
  wire popcount30_uea4_core_203;
  wire popcount30_uea4_core_204;
  wire popcount30_uea4_core_205;
  wire popcount30_uea4_core_206;
  wire popcount30_uea4_core_208;
  wire popcount30_uea4_core_209;
  wire popcount30_uea4_core_210;
  wire popcount30_uea4_core_212;
  wire popcount30_uea4_core_213;

  assign popcount30_uea4_core_032 = ~input_a[1];
  assign popcount30_uea4_core_033 = input_a[28] & input_a[25];
  assign popcount30_uea4_core_038 = input_a[19] & input_a[24];
  assign popcount30_uea4_core_041 = input_a[7] ^ input_a[20];
  assign popcount30_uea4_core_043 = ~(input_a[1] & input_a[3]);
  assign popcount30_uea4_core_044 = ~(input_a[8] & input_a[10]);
  assign popcount30_uea4_core_045 = input_a[24] & input_a[6];
  assign popcount30_uea4_core_046 = ~(input_a[28] & input_a[0]);
  assign popcount30_uea4_core_048 = input_a[14] | input_a[12];
  assign popcount30_uea4_core_049 = input_a[25] | input_a[18];
  assign popcount30_uea4_core_050 = ~(input_a[29] & input_a[7]);
  assign popcount30_uea4_core_053 = ~(input_a[18] & input_a[0]);
  assign popcount30_uea4_core_054 = ~(input_a[12] & input_a[6]);
  assign popcount30_uea4_core_055 = ~input_a[18];
  assign popcount30_uea4_core_056 = input_a[8] ^ input_a[8];
  assign popcount30_uea4_core_057 = ~(input_a[15] | input_a[2]);
  assign popcount30_uea4_core_060 = ~input_a[11];
  assign popcount30_uea4_core_061 = ~(input_a[8] & input_a[5]);
  assign popcount30_uea4_core_062 = input_a[9] & input_a[24];
  assign popcount30_uea4_core_063 = input_a[8] ^ input_a[21];
  assign popcount30_uea4_core_066 = ~(input_a[1] | input_a[14]);
  assign popcount30_uea4_core_067 = ~(input_a[27] ^ input_a[0]);
  assign popcount30_uea4_core_068 = ~(input_a[6] & input_a[8]);
  assign popcount30_uea4_core_069 = ~(input_a[13] & input_a[14]);
  assign popcount30_uea4_core_070 = input_a[20] ^ input_a[2];
  assign popcount30_uea4_core_071 = input_a[1] & input_a[7];
  assign popcount30_uea4_core_072 = ~(input_a[16] ^ input_a[23]);
  assign popcount30_uea4_core_073 = ~(input_a[18] ^ input_a[21]);
  assign popcount30_uea4_core_074 = input_a[25] & input_a[4];
  assign popcount30_uea4_core_075 = ~(input_a[23] ^ input_a[12]);
  assign popcount30_uea4_core_078 = input_a[3] ^ input_a[3];
  assign popcount30_uea4_core_079 = ~(input_a[26] ^ input_a[16]);
  assign popcount30_uea4_core_081 = ~(input_a[14] ^ input_a[15]);
  assign popcount30_uea4_core_083 = ~(input_a[20] ^ input_a[22]);
  assign popcount30_uea4_core_084 = input_a[6] | input_a[16];
  assign popcount30_uea4_core_085 = ~input_a[11];
  assign popcount30_uea4_core_086 = ~(input_a[24] | input_a[19]);
  assign popcount30_uea4_core_087 = ~input_a[4];
  assign popcount30_uea4_core_091 = ~(input_a[9] ^ input_a[1]);
  assign popcount30_uea4_core_092 = ~input_a[11];
  assign popcount30_uea4_core_093_not = ~input_a[0];
  assign popcount30_uea4_core_094 = input_a[9] | input_a[6];
  assign popcount30_uea4_core_096 = input_a[16] ^ input_a[13];
  assign popcount30_uea4_core_097 = ~(input_a[0] ^ input_a[0]);
  assign popcount30_uea4_core_098 = ~(input_a[14] & input_a[5]);
  assign popcount30_uea4_core_101 = ~(input_a[15] ^ input_a[24]);
  assign popcount30_uea4_core_102 = ~(input_a[24] | input_a[28]);
  assign popcount30_uea4_core_103 = ~(input_a[21] | input_a[4]);
  assign popcount30_uea4_core_105 = ~input_a[29];
  assign popcount30_uea4_core_106 = input_a[29] ^ input_a[3];
  assign popcount30_uea4_core_107 = input_a[12] & input_a[11];
  assign popcount30_uea4_core_108 = ~(input_a[11] | input_a[26]);
  assign popcount30_uea4_core_109 = input_a[20] & input_a[25];
  assign popcount30_uea4_core_110 = ~(input_a[11] | input_a[9]);
  assign popcount30_uea4_core_112 = ~(input_a[4] ^ input_a[0]);
  assign popcount30_uea4_core_113 = input_a[0] & input_a[27];
  assign popcount30_uea4_core_114 = input_a[8] ^ input_a[6];
  assign popcount30_uea4_core_116 = input_a[3] | input_a[5];
  assign popcount30_uea4_core_117 = input_a[17] & input_a[8];
  assign popcount30_uea4_core_118 = ~(input_a[16] & input_a[18]);
  assign popcount30_uea4_core_119 = input_a[24] & input_a[2];
  assign popcount30_uea4_core_120 = input_a[29] & input_a[22];
  assign popcount30_uea4_core_121 = input_a[17] | input_a[9];
  assign popcount30_uea4_core_123 = input_a[8] ^ input_a[2];
  assign popcount30_uea4_core_126 = ~(input_a[1] | input_a[14]);
  assign popcount30_uea4_core_127 = input_a[15] & input_a[28];
  assign popcount30_uea4_core_128 = input_a[15] | input_a[24];
  assign popcount30_uea4_core_129 = ~input_a[23];
  assign popcount30_uea4_core_131 = input_a[5] | input_a[13];
  assign popcount30_uea4_core_132 = input_a[26] & input_a[0];
  assign popcount30_uea4_core_133 = input_a[0] ^ input_a[23];
  assign popcount30_uea4_core_135 = ~input_a[16];
  assign popcount30_uea4_core_137 = ~input_a[22];
  assign popcount30_uea4_core_138 = ~(input_a[0] | input_a[28]);
  assign popcount30_uea4_core_140 = input_a[2] & input_a[10];
  assign popcount30_uea4_core_143 = ~(input_a[10] ^ input_a[11]);
  assign popcount30_uea4_core_145 = input_a[18] | input_a[6];
  assign popcount30_uea4_core_146 = input_a[18] & input_a[1];
  assign popcount30_uea4_core_147 = ~(input_a[23] | input_a[10]);
  assign popcount30_uea4_core_148 = input_a[26] | input_a[11];
  assign popcount30_uea4_core_149 = input_a[11] & input_a[3];
  assign popcount30_uea4_core_151 = ~input_a[16];
  assign popcount30_uea4_core_155 = ~(input_a[3] | input_a[1]);
  assign popcount30_uea4_core_157 = ~(input_a[0] ^ input_a[11]);
  assign popcount30_uea4_core_158 = ~(input_a[3] & input_a[14]);
  assign popcount30_uea4_core_159 = input_a[23] ^ input_a[26];
  assign popcount30_uea4_core_160 = input_a[23] & input_a[28];
  assign popcount30_uea4_core_161 = input_a[8] & input_a[18];
  assign popcount30_uea4_core_162 = input_a[16] & input_a[3];
  assign popcount30_uea4_core_163 = input_a[18] & input_a[7];
  assign popcount30_uea4_core_164 = ~(input_a[13] | input_a[22]);
  assign popcount30_uea4_core_165 = input_a[26] | input_a[16];
  assign popcount30_uea4_core_166 = ~(input_a[26] ^ input_a[14]);
  assign popcount30_uea4_core_167 = ~(input_a[27] | input_a[4]);
  assign popcount30_uea4_core_168 = input_a[29] & input_a[17];
  assign popcount30_uea4_core_169 = ~input_a[21];
  assign popcount30_uea4_core_171 = ~(input_a[29] & input_a[17]);
  assign popcount30_uea4_core_173 = ~input_a[2];
  assign popcount30_uea4_core_174 = ~(input_a[9] | input_a[9]);
  assign popcount30_uea4_core_175 = input_a[17] | input_a[14];
  assign popcount30_uea4_core_177 = ~(input_a[15] ^ input_a[10]);
  assign popcount30_uea4_core_178 = input_a[27] & input_a[9];
  assign popcount30_uea4_core_179 = input_a[27] & input_a[12];
  assign popcount30_uea4_core_180 = ~(input_a[0] | input_a[12]);
  assign popcount30_uea4_core_181 = input_a[10] & input_a[12];
  assign popcount30_uea4_core_182 = ~(input_a[8] | input_a[18]);
  assign popcount30_uea4_core_183 = ~(input_a[25] ^ input_a[27]);
  assign popcount30_uea4_core_186 = ~(input_a[9] | input_a[24]);
  assign popcount30_uea4_core_187 = ~(input_a[8] ^ input_a[3]);
  assign popcount30_uea4_core_194 = input_a[11] & input_a[4];
  assign popcount30_uea4_core_196 = ~(input_a[24] & input_a[24]);
  assign popcount30_uea4_core_197 = ~(input_a[24] | input_a[3]);
  assign popcount30_uea4_core_198 = input_a[19] & input_a[2];
  assign popcount30_uea4_core_199 = ~(input_a[15] & input_a[11]);
  assign popcount30_uea4_core_200 = input_a[15] & input_a[14];
  assign popcount30_uea4_core_201 = ~(input_a[6] & input_a[24]);
  assign popcount30_uea4_core_202 = ~(input_a[10] | input_a[27]);
  assign popcount30_uea4_core_203 = input_a[15] | input_a[23];
  assign popcount30_uea4_core_204 = input_a[15] | input_a[24];
  assign popcount30_uea4_core_205 = input_a[0] & input_a[2];
  assign popcount30_uea4_core_206 = input_a[12] & input_a[9];
  assign popcount30_uea4_core_208 = input_a[3] & input_a[0];
  assign popcount30_uea4_core_209 = input_a[12] ^ input_a[11];
  assign popcount30_uea4_core_210 = ~(input_a[20] | input_a[12]);
  assign popcount30_uea4_core_212 = ~(input_a[19] ^ input_a[15]);
  assign popcount30_uea4_core_213 = input_a[5] & input_a[4];

  assign popcount30_uea4_out[0] = input_a[20];
  assign popcount30_uea4_out[1] = input_a[29];
  assign popcount30_uea4_out[2] = popcount30_uea4_core_201;
  assign popcount30_uea4_out[3] = popcount30_uea4_core_201;
  assign popcount30_uea4_out[4] = popcount30_uea4_core_045;
endmodule