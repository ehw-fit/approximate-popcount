// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.93621
// WCE=28.0
// EP=0.939096%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount40_5o2k(input [39:0] input_a, output [5:0] popcount40_5o2k_out);
  wire popcount40_5o2k_core_042;
  wire popcount40_5o2k_core_047;
  wire popcount40_5o2k_core_048;
  wire popcount40_5o2k_core_050;
  wire popcount40_5o2k_core_052;
  wire popcount40_5o2k_core_054;
  wire popcount40_5o2k_core_055;
  wire popcount40_5o2k_core_056;
  wire popcount40_5o2k_core_059;
  wire popcount40_5o2k_core_060;
  wire popcount40_5o2k_core_062;
  wire popcount40_5o2k_core_063;
  wire popcount40_5o2k_core_064;
  wire popcount40_5o2k_core_065;
  wire popcount40_5o2k_core_066;
  wire popcount40_5o2k_core_067;
  wire popcount40_5o2k_core_069;
  wire popcount40_5o2k_core_070;
  wire popcount40_5o2k_core_071;
  wire popcount40_5o2k_core_072;
  wire popcount40_5o2k_core_073;
  wire popcount40_5o2k_core_074;
  wire popcount40_5o2k_core_075;
  wire popcount40_5o2k_core_076;
  wire popcount40_5o2k_core_077;
  wire popcount40_5o2k_core_078;
  wire popcount40_5o2k_core_079_not;
  wire popcount40_5o2k_core_080;
  wire popcount40_5o2k_core_081;
  wire popcount40_5o2k_core_083;
  wire popcount40_5o2k_core_084;
  wire popcount40_5o2k_core_085;
  wire popcount40_5o2k_core_086;
  wire popcount40_5o2k_core_087;
  wire popcount40_5o2k_core_088;
  wire popcount40_5o2k_core_089;
  wire popcount40_5o2k_core_090;
  wire popcount40_5o2k_core_091;
  wire popcount40_5o2k_core_092;
  wire popcount40_5o2k_core_093;
  wire popcount40_5o2k_core_094;
  wire popcount40_5o2k_core_096;
  wire popcount40_5o2k_core_102;
  wire popcount40_5o2k_core_104;
  wire popcount40_5o2k_core_105;
  wire popcount40_5o2k_core_106;
  wire popcount40_5o2k_core_109_not;
  wire popcount40_5o2k_core_111;
  wire popcount40_5o2k_core_113;
  wire popcount40_5o2k_core_114;
  wire popcount40_5o2k_core_115;
  wire popcount40_5o2k_core_116;
  wire popcount40_5o2k_core_117;
  wire popcount40_5o2k_core_120;
  wire popcount40_5o2k_core_121;
  wire popcount40_5o2k_core_123;
  wire popcount40_5o2k_core_128;
  wire popcount40_5o2k_core_129;
  wire popcount40_5o2k_core_130;
  wire popcount40_5o2k_core_131;
  wire popcount40_5o2k_core_132;
  wire popcount40_5o2k_core_133;
  wire popcount40_5o2k_core_134;
  wire popcount40_5o2k_core_135;
  wire popcount40_5o2k_core_136;
  wire popcount40_5o2k_core_137;
  wire popcount40_5o2k_core_140;
  wire popcount40_5o2k_core_141;
  wire popcount40_5o2k_core_142;
  wire popcount40_5o2k_core_144_not;
  wire popcount40_5o2k_core_148_not;
  wire popcount40_5o2k_core_149;
  wire popcount40_5o2k_core_150;
  wire popcount40_5o2k_core_151;
  wire popcount40_5o2k_core_152;
  wire popcount40_5o2k_core_153;
  wire popcount40_5o2k_core_154;
  wire popcount40_5o2k_core_157;
  wire popcount40_5o2k_core_158;
  wire popcount40_5o2k_core_159;
  wire popcount40_5o2k_core_161;
  wire popcount40_5o2k_core_163;
  wire popcount40_5o2k_core_165;
  wire popcount40_5o2k_core_166;
  wire popcount40_5o2k_core_168;
  wire popcount40_5o2k_core_169;
  wire popcount40_5o2k_core_173;
  wire popcount40_5o2k_core_174;
  wire popcount40_5o2k_core_175;
  wire popcount40_5o2k_core_176;
  wire popcount40_5o2k_core_177;
  wire popcount40_5o2k_core_178;
  wire popcount40_5o2k_core_179;
  wire popcount40_5o2k_core_180;
  wire popcount40_5o2k_core_182;
  wire popcount40_5o2k_core_183;
  wire popcount40_5o2k_core_184;
  wire popcount40_5o2k_core_187_not;
  wire popcount40_5o2k_core_189;
  wire popcount40_5o2k_core_190;
  wire popcount40_5o2k_core_191;
  wire popcount40_5o2k_core_193;
  wire popcount40_5o2k_core_195;
  wire popcount40_5o2k_core_196;
  wire popcount40_5o2k_core_198;
  wire popcount40_5o2k_core_199;
  wire popcount40_5o2k_core_200;
  wire popcount40_5o2k_core_201;
  wire popcount40_5o2k_core_203;
  wire popcount40_5o2k_core_205;
  wire popcount40_5o2k_core_207;
  wire popcount40_5o2k_core_208;
  wire popcount40_5o2k_core_209;
  wire popcount40_5o2k_core_210;
  wire popcount40_5o2k_core_211;
  wire popcount40_5o2k_core_214;
  wire popcount40_5o2k_core_215;
  wire popcount40_5o2k_core_216;
  wire popcount40_5o2k_core_217;
  wire popcount40_5o2k_core_219;
  wire popcount40_5o2k_core_220;
  wire popcount40_5o2k_core_221;
  wire popcount40_5o2k_core_222;
  wire popcount40_5o2k_core_223_not;
  wire popcount40_5o2k_core_225;
  wire popcount40_5o2k_core_226;
  wire popcount40_5o2k_core_227;
  wire popcount40_5o2k_core_228;
  wire popcount40_5o2k_core_229;
  wire popcount40_5o2k_core_230;
  wire popcount40_5o2k_core_231;
  wire popcount40_5o2k_core_232;
  wire popcount40_5o2k_core_233;
  wire popcount40_5o2k_core_235;
  wire popcount40_5o2k_core_236;
  wire popcount40_5o2k_core_237;
  wire popcount40_5o2k_core_238;
  wire popcount40_5o2k_core_239;
  wire popcount40_5o2k_core_241;
  wire popcount40_5o2k_core_242_not;
  wire popcount40_5o2k_core_243;
  wire popcount40_5o2k_core_244;
  wire popcount40_5o2k_core_247_not;
  wire popcount40_5o2k_core_248;
  wire popcount40_5o2k_core_251;
  wire popcount40_5o2k_core_253;
  wire popcount40_5o2k_core_256;
  wire popcount40_5o2k_core_258;
  wire popcount40_5o2k_core_260;
  wire popcount40_5o2k_core_261;
  wire popcount40_5o2k_core_263;
  wire popcount40_5o2k_core_265;
  wire popcount40_5o2k_core_266;
  wire popcount40_5o2k_core_267;
  wire popcount40_5o2k_core_270;
  wire popcount40_5o2k_core_273;
  wire popcount40_5o2k_core_274;
  wire popcount40_5o2k_core_276;
  wire popcount40_5o2k_core_277;
  wire popcount40_5o2k_core_278;
  wire popcount40_5o2k_core_282;
  wire popcount40_5o2k_core_284;
  wire popcount40_5o2k_core_288;
  wire popcount40_5o2k_core_290;
  wire popcount40_5o2k_core_291;
  wire popcount40_5o2k_core_293;
  wire popcount40_5o2k_core_295;
  wire popcount40_5o2k_core_296;
  wire popcount40_5o2k_core_299;
  wire popcount40_5o2k_core_300;
  wire popcount40_5o2k_core_302;
  wire popcount40_5o2k_core_304;
  wire popcount40_5o2k_core_305;
  wire popcount40_5o2k_core_306;
  wire popcount40_5o2k_core_307;
  wire popcount40_5o2k_core_308;
  wire popcount40_5o2k_core_309_not;
  wire popcount40_5o2k_core_310;
  wire popcount40_5o2k_core_312;

  assign popcount40_5o2k_core_042 = input_a[8] | input_a[0];
  assign popcount40_5o2k_core_047 = ~(input_a[2] & input_a[15]);
  assign popcount40_5o2k_core_048 = ~(input_a[3] | input_a[15]);
  assign popcount40_5o2k_core_050 = ~(input_a[11] ^ input_a[29]);
  assign popcount40_5o2k_core_052 = input_a[22] & input_a[17];
  assign popcount40_5o2k_core_054 = input_a[15] ^ input_a[33];
  assign popcount40_5o2k_core_055 = ~input_a[11];
  assign popcount40_5o2k_core_056 = input_a[9] ^ input_a[11];
  assign popcount40_5o2k_core_059 = input_a[36] ^ input_a[34];
  assign popcount40_5o2k_core_060 = ~(input_a[8] | input_a[35]);
  assign popcount40_5o2k_core_062 = input_a[25] & input_a[17];
  assign popcount40_5o2k_core_063 = input_a[3] & input_a[26];
  assign popcount40_5o2k_core_064 = ~(input_a[5] & input_a[21]);
  assign popcount40_5o2k_core_065 = ~(input_a[4] | input_a[38]);
  assign popcount40_5o2k_core_066 = ~(input_a[29] | input_a[20]);
  assign popcount40_5o2k_core_067 = input_a[26] ^ input_a[12];
  assign popcount40_5o2k_core_069 = input_a[35] & input_a[13];
  assign popcount40_5o2k_core_070 = ~(input_a[0] | input_a[6]);
  assign popcount40_5o2k_core_071 = input_a[7] & input_a[29];
  assign popcount40_5o2k_core_072 = input_a[25] ^ input_a[2];
  assign popcount40_5o2k_core_073 = input_a[3] & input_a[28];
  assign popcount40_5o2k_core_074 = ~(input_a[4] ^ input_a[36]);
  assign popcount40_5o2k_core_075 = input_a[3] & input_a[1];
  assign popcount40_5o2k_core_076 = ~input_a[2];
  assign popcount40_5o2k_core_077 = ~(input_a[3] | input_a[0]);
  assign popcount40_5o2k_core_078 = ~(input_a[16] ^ input_a[38]);
  assign popcount40_5o2k_core_079_not = ~input_a[18];
  assign popcount40_5o2k_core_080 = ~(input_a[2] ^ input_a[24]);
  assign popcount40_5o2k_core_081 = ~(input_a[31] ^ input_a[36]);
  assign popcount40_5o2k_core_083 = input_a[24] & input_a[19];
  assign popcount40_5o2k_core_084 = input_a[5] ^ input_a[6];
  assign popcount40_5o2k_core_085 = ~(input_a[16] | input_a[33]);
  assign popcount40_5o2k_core_086 = ~(input_a[17] & input_a[31]);
  assign popcount40_5o2k_core_087 = ~(input_a[7] ^ input_a[7]);
  assign popcount40_5o2k_core_088 = ~input_a[10];
  assign popcount40_5o2k_core_089 = ~(input_a[0] | input_a[19]);
  assign popcount40_5o2k_core_090 = input_a[28] & input_a[9];
  assign popcount40_5o2k_core_091 = input_a[30] ^ input_a[29];
  assign popcount40_5o2k_core_092 = ~input_a[3];
  assign popcount40_5o2k_core_093 = input_a[24] ^ input_a[19];
  assign popcount40_5o2k_core_094 = ~input_a[1];
  assign popcount40_5o2k_core_096 = ~input_a[2];
  assign popcount40_5o2k_core_102 = ~(input_a[0] & input_a[22]);
  assign popcount40_5o2k_core_104 = input_a[7] | input_a[31];
  assign popcount40_5o2k_core_105 = input_a[29] | input_a[27];
  assign popcount40_5o2k_core_106 = input_a[37] & input_a[20];
  assign popcount40_5o2k_core_109_not = ~input_a[37];
  assign popcount40_5o2k_core_111 = input_a[38] | input_a[6];
  assign popcount40_5o2k_core_113 = input_a[6] ^ input_a[32];
  assign popcount40_5o2k_core_114 = input_a[37] ^ input_a[21];
  assign popcount40_5o2k_core_115 = ~(input_a[27] & input_a[27]);
  assign popcount40_5o2k_core_116 = input_a[23] | input_a[25];
  assign popcount40_5o2k_core_117 = ~(input_a[28] | input_a[6]);
  assign popcount40_5o2k_core_120 = input_a[35] ^ input_a[8];
  assign popcount40_5o2k_core_121 = ~(input_a[7] & input_a[38]);
  assign popcount40_5o2k_core_123 = ~(input_a[10] & input_a[5]);
  assign popcount40_5o2k_core_128 = input_a[3] & input_a[5];
  assign popcount40_5o2k_core_129 = ~(input_a[37] | input_a[6]);
  assign popcount40_5o2k_core_130 = input_a[14] | input_a[6];
  assign popcount40_5o2k_core_131 = ~input_a[16];
  assign popcount40_5o2k_core_132 = ~input_a[36];
  assign popcount40_5o2k_core_133 = ~(input_a[33] & input_a[34]);
  assign popcount40_5o2k_core_134 = ~(input_a[4] ^ input_a[29]);
  assign popcount40_5o2k_core_135 = ~(input_a[7] & input_a[19]);
  assign popcount40_5o2k_core_136 = input_a[2] & input_a[39];
  assign popcount40_5o2k_core_137 = input_a[7] & input_a[33];
  assign popcount40_5o2k_core_140 = ~input_a[2];
  assign popcount40_5o2k_core_141 = ~(input_a[5] & input_a[9]);
  assign popcount40_5o2k_core_142 = input_a[2] ^ input_a[36];
  assign popcount40_5o2k_core_144_not = ~input_a[2];
  assign popcount40_5o2k_core_148_not = ~input_a[25];
  assign popcount40_5o2k_core_149 = ~(input_a[0] ^ input_a[36]);
  assign popcount40_5o2k_core_150 = input_a[14] ^ input_a[34];
  assign popcount40_5o2k_core_151 = ~(input_a[28] | input_a[19]);
  assign popcount40_5o2k_core_152 = input_a[30] ^ input_a[32];
  assign popcount40_5o2k_core_153 = ~(input_a[36] ^ input_a[29]);
  assign popcount40_5o2k_core_154 = input_a[18] | input_a[31];
  assign popcount40_5o2k_core_157 = ~(input_a[4] & input_a[19]);
  assign popcount40_5o2k_core_158 = ~input_a[23];
  assign popcount40_5o2k_core_159 = ~(input_a[38] | input_a[24]);
  assign popcount40_5o2k_core_161 = ~(input_a[19] & input_a[21]);
  assign popcount40_5o2k_core_163 = ~(input_a[25] ^ input_a[21]);
  assign popcount40_5o2k_core_165 = input_a[2] ^ input_a[18];
  assign popcount40_5o2k_core_166 = input_a[10] & input_a[0];
  assign popcount40_5o2k_core_168 = ~input_a[26];
  assign popcount40_5o2k_core_169 = input_a[1] & input_a[34];
  assign popcount40_5o2k_core_173 = ~(input_a[21] | input_a[35]);
  assign popcount40_5o2k_core_174 = input_a[22] | input_a[28];
  assign popcount40_5o2k_core_175 = input_a[27] & input_a[29];
  assign popcount40_5o2k_core_176 = ~(input_a[9] | input_a[33]);
  assign popcount40_5o2k_core_177 = ~(input_a[26] ^ input_a[11]);
  assign popcount40_5o2k_core_178 = input_a[13] & input_a[23];
  assign popcount40_5o2k_core_179 = ~input_a[38];
  assign popcount40_5o2k_core_180 = input_a[17] & input_a[29];
  assign popcount40_5o2k_core_182 = input_a[34] & input_a[34];
  assign popcount40_5o2k_core_183 = ~(input_a[33] | input_a[31]);
  assign popcount40_5o2k_core_184 = ~(input_a[29] & input_a[7]);
  assign popcount40_5o2k_core_187_not = ~input_a[37];
  assign popcount40_5o2k_core_189 = ~(input_a[10] | input_a[6]);
  assign popcount40_5o2k_core_190 = input_a[39] & input_a[33];
  assign popcount40_5o2k_core_191 = input_a[22] & input_a[28];
  assign popcount40_5o2k_core_193 = input_a[23] ^ input_a[32];
  assign popcount40_5o2k_core_195 = ~(input_a[9] & input_a[9]);
  assign popcount40_5o2k_core_196 = ~(input_a[12] ^ input_a[27]);
  assign popcount40_5o2k_core_198 = input_a[36] | input_a[7];
  assign popcount40_5o2k_core_199 = input_a[18] & input_a[29];
  assign popcount40_5o2k_core_200 = ~(input_a[15] & input_a[31]);
  assign popcount40_5o2k_core_201 = input_a[32] | input_a[37];
  assign popcount40_5o2k_core_203 = input_a[2] ^ input_a[26];
  assign popcount40_5o2k_core_205 = ~(input_a[34] & input_a[30]);
  assign popcount40_5o2k_core_207 = ~(input_a[6] & input_a[1]);
  assign popcount40_5o2k_core_208 = ~(input_a[7] & input_a[13]);
  assign popcount40_5o2k_core_209 = input_a[28] ^ input_a[17];
  assign popcount40_5o2k_core_210 = ~(input_a[2] & input_a[35]);
  assign popcount40_5o2k_core_211 = ~(input_a[18] & input_a[24]);
  assign popcount40_5o2k_core_214 = ~input_a[29];
  assign popcount40_5o2k_core_215 = input_a[22] & input_a[37];
  assign popcount40_5o2k_core_216 = ~input_a[32];
  assign popcount40_5o2k_core_217 = ~(input_a[35] ^ input_a[39]);
  assign popcount40_5o2k_core_219 = input_a[15] & input_a[20];
  assign popcount40_5o2k_core_220 = ~input_a[35];
  assign popcount40_5o2k_core_221 = ~input_a[22];
  assign popcount40_5o2k_core_222 = input_a[32] & input_a[27];
  assign popcount40_5o2k_core_223_not = ~input_a[23];
  assign popcount40_5o2k_core_225 = input_a[29] | input_a[5];
  assign popcount40_5o2k_core_226 = input_a[7] & input_a[19];
  assign popcount40_5o2k_core_227 = input_a[36] & input_a[10];
  assign popcount40_5o2k_core_228 = ~(input_a[32] & input_a[21]);
  assign popcount40_5o2k_core_229 = input_a[9] ^ input_a[35];
  assign popcount40_5o2k_core_230 = ~(input_a[2] & input_a[4]);
  assign popcount40_5o2k_core_231 = ~(input_a[37] | input_a[29]);
  assign popcount40_5o2k_core_232 = ~input_a[9];
  assign popcount40_5o2k_core_233 = input_a[7] & input_a[35];
  assign popcount40_5o2k_core_235 = ~input_a[9];
  assign popcount40_5o2k_core_236 = ~input_a[10];
  assign popcount40_5o2k_core_237 = ~input_a[1];
  assign popcount40_5o2k_core_238 = ~(input_a[31] | input_a[17]);
  assign popcount40_5o2k_core_239 = input_a[11] & input_a[28];
  assign popcount40_5o2k_core_241 = ~(input_a[11] & input_a[18]);
  assign popcount40_5o2k_core_242_not = ~input_a[24];
  assign popcount40_5o2k_core_243 = input_a[32] | input_a[39];
  assign popcount40_5o2k_core_244 = ~(input_a[33] ^ input_a[13]);
  assign popcount40_5o2k_core_247_not = ~input_a[34];
  assign popcount40_5o2k_core_248 = ~(input_a[4] & input_a[29]);
  assign popcount40_5o2k_core_251 = input_a[22] | input_a[30];
  assign popcount40_5o2k_core_253 = ~input_a[18];
  assign popcount40_5o2k_core_256 = ~(input_a[19] ^ input_a[28]);
  assign popcount40_5o2k_core_258 = ~(input_a[0] | input_a[32]);
  assign popcount40_5o2k_core_260 = input_a[14] ^ input_a[13];
  assign popcount40_5o2k_core_261 = ~(input_a[19] ^ input_a[34]);
  assign popcount40_5o2k_core_263 = ~(input_a[16] & input_a[29]);
  assign popcount40_5o2k_core_265 = input_a[6] ^ input_a[6];
  assign popcount40_5o2k_core_266 = ~(input_a[16] | input_a[19]);
  assign popcount40_5o2k_core_267 = ~input_a[11];
  assign popcount40_5o2k_core_270 = ~(input_a[25] | input_a[23]);
  assign popcount40_5o2k_core_273 = ~(input_a[35] & input_a[0]);
  assign popcount40_5o2k_core_274 = input_a[32] ^ input_a[32];
  assign popcount40_5o2k_core_276 = ~(input_a[32] ^ input_a[1]);
  assign popcount40_5o2k_core_277 = ~(input_a[13] | input_a[23]);
  assign popcount40_5o2k_core_278 = input_a[19] & input_a[11];
  assign popcount40_5o2k_core_282 = input_a[23] ^ input_a[3];
  assign popcount40_5o2k_core_284 = input_a[19] ^ input_a[5];
  assign popcount40_5o2k_core_288 = input_a[19] & input_a[28];
  assign popcount40_5o2k_core_290 = input_a[9] ^ input_a[24];
  assign popcount40_5o2k_core_291 = input_a[33] ^ input_a[31];
  assign popcount40_5o2k_core_293 = input_a[28] ^ input_a[8];
  assign popcount40_5o2k_core_295 = input_a[3] | input_a[17];
  assign popcount40_5o2k_core_296 = ~(input_a[5] ^ input_a[8]);
  assign popcount40_5o2k_core_299 = input_a[2] ^ input_a[6];
  assign popcount40_5o2k_core_300 = ~(input_a[25] | input_a[15]);
  assign popcount40_5o2k_core_302 = input_a[17] & input_a[15];
  assign popcount40_5o2k_core_304 = ~(input_a[34] | input_a[27]);
  assign popcount40_5o2k_core_305 = ~(input_a[3] & input_a[7]);
  assign popcount40_5o2k_core_306 = ~(input_a[15] ^ input_a[25]);
  assign popcount40_5o2k_core_307 = input_a[17] & input_a[37];
  assign popcount40_5o2k_core_308 = input_a[8] | input_a[29];
  assign popcount40_5o2k_core_309_not = ~input_a[12];
  assign popcount40_5o2k_core_310 = input_a[10] & input_a[30];
  assign popcount40_5o2k_core_312 = ~(input_a[11] & input_a[5]);

  assign popcount40_5o2k_out[0] = 1'b0;
  assign popcount40_5o2k_out[1] = input_a[19];
  assign popcount40_5o2k_out[2] = input_a[19];
  assign popcount40_5o2k_out[3] = input_a[14];
  assign popcount40_5o2k_out[4] = 1'b1;
  assign popcount40_5o2k_out[5] = 1'b0;
endmodule