// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.55848
// WCE=24.0
// EP=0.976718%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_6cry(input [26:0] input_a, output [4:0] popcount27_6cry_out);
  wire popcount27_6cry_core_029;
  wire popcount27_6cry_core_032;
  wire popcount27_6cry_core_033;
  wire popcount27_6cry_core_034;
  wire popcount27_6cry_core_035;
  wire popcount27_6cry_core_036;
  wire popcount27_6cry_core_038_not;
  wire popcount27_6cry_core_039;
  wire popcount27_6cry_core_040;
  wire popcount27_6cry_core_041;
  wire popcount27_6cry_core_043;
  wire popcount27_6cry_core_045;
  wire popcount27_6cry_core_046;
  wire popcount27_6cry_core_048;
  wire popcount27_6cry_core_049;
  wire popcount27_6cry_core_050;
  wire popcount27_6cry_core_052;
  wire popcount27_6cry_core_053;
  wire popcount27_6cry_core_054;
  wire popcount27_6cry_core_055;
  wire popcount27_6cry_core_057;
  wire popcount27_6cry_core_058;
  wire popcount27_6cry_core_059;
  wire popcount27_6cry_core_060;
  wire popcount27_6cry_core_061;
  wire popcount27_6cry_core_064;
  wire popcount27_6cry_core_065;
  wire popcount27_6cry_core_066;
  wire popcount27_6cry_core_067;
  wire popcount27_6cry_core_068;
  wire popcount27_6cry_core_069;
  wire popcount27_6cry_core_070;
  wire popcount27_6cry_core_071;
  wire popcount27_6cry_core_072;
  wire popcount27_6cry_core_075;
  wire popcount27_6cry_core_076;
  wire popcount27_6cry_core_079;
  wire popcount27_6cry_core_080;
  wire popcount27_6cry_core_081;
  wire popcount27_6cry_core_082;
  wire popcount27_6cry_core_083;
  wire popcount27_6cry_core_084;
  wire popcount27_6cry_core_086;
  wire popcount27_6cry_core_087;
  wire popcount27_6cry_core_088;
  wire popcount27_6cry_core_090;
  wire popcount27_6cry_core_091;
  wire popcount27_6cry_core_092;
  wire popcount27_6cry_core_093;
  wire popcount27_6cry_core_094;
  wire popcount27_6cry_core_096;
  wire popcount27_6cry_core_099;
  wire popcount27_6cry_core_101;
  wire popcount27_6cry_core_104;
  wire popcount27_6cry_core_106;
  wire popcount27_6cry_core_107;
  wire popcount27_6cry_core_108;
  wire popcount27_6cry_core_113;
  wire popcount27_6cry_core_114;
  wire popcount27_6cry_core_117;
  wire popcount27_6cry_core_118;
  wire popcount27_6cry_core_119;
  wire popcount27_6cry_core_120;
  wire popcount27_6cry_core_121;
  wire popcount27_6cry_core_123;
  wire popcount27_6cry_core_126;
  wire popcount27_6cry_core_127;
  wire popcount27_6cry_core_128;
  wire popcount27_6cry_core_130;
  wire popcount27_6cry_core_131;
  wire popcount27_6cry_core_133;
  wire popcount27_6cry_core_136;
  wire popcount27_6cry_core_137;
  wire popcount27_6cry_core_139;
  wire popcount27_6cry_core_140;
  wire popcount27_6cry_core_142;
  wire popcount27_6cry_core_144;
  wire popcount27_6cry_core_146;
  wire popcount27_6cry_core_147;
  wire popcount27_6cry_core_148;
  wire popcount27_6cry_core_149;
  wire popcount27_6cry_core_154;
  wire popcount27_6cry_core_156;
  wire popcount27_6cry_core_157;
  wire popcount27_6cry_core_158;
  wire popcount27_6cry_core_161;
  wire popcount27_6cry_core_162;
  wire popcount27_6cry_core_163;
  wire popcount27_6cry_core_165;
  wire popcount27_6cry_core_167;
  wire popcount27_6cry_core_168;
  wire popcount27_6cry_core_169;
  wire popcount27_6cry_core_170;
  wire popcount27_6cry_core_171;
  wire popcount27_6cry_core_172;
  wire popcount27_6cry_core_175;
  wire popcount27_6cry_core_176;
  wire popcount27_6cry_core_177;
  wire popcount27_6cry_core_179;
  wire popcount27_6cry_core_182;
  wire popcount27_6cry_core_183;
  wire popcount27_6cry_core_186;
  wire popcount27_6cry_core_187;
  wire popcount27_6cry_core_188;
  wire popcount27_6cry_core_190;
  wire popcount27_6cry_core_192;
  wire popcount27_6cry_core_193;
  wire popcount27_6cry_core_194;
  wire popcount27_6cry_core_195;

  assign popcount27_6cry_core_029 = input_a[16] & input_a[1];
  assign popcount27_6cry_core_032 = input_a[24] & input_a[21];
  assign popcount27_6cry_core_033 = ~(input_a[26] & input_a[7]);
  assign popcount27_6cry_core_034 = input_a[26] | input_a[7];
  assign popcount27_6cry_core_035 = input_a[1] ^ input_a[10];
  assign popcount27_6cry_core_036 = input_a[15] | input_a[1];
  assign popcount27_6cry_core_038_not = ~input_a[10];
  assign popcount27_6cry_core_039 = input_a[16] & input_a[1];
  assign popcount27_6cry_core_040 = input_a[10] & input_a[7];
  assign popcount27_6cry_core_041 = ~(input_a[21] & input_a[20]);
  assign popcount27_6cry_core_043 = input_a[10] & input_a[9];
  assign popcount27_6cry_core_045 = input_a[1] | input_a[23];
  assign popcount27_6cry_core_046 = ~(input_a[21] ^ input_a[2]);
  assign popcount27_6cry_core_048 = ~(input_a[17] | input_a[25]);
  assign popcount27_6cry_core_049 = ~(input_a[1] ^ input_a[20]);
  assign popcount27_6cry_core_050 = ~input_a[1];
  assign popcount27_6cry_core_052 = ~(input_a[5] & input_a[19]);
  assign popcount27_6cry_core_053 = input_a[26] ^ input_a[4];
  assign popcount27_6cry_core_054 = ~input_a[13];
  assign popcount27_6cry_core_055 = ~input_a[24];
  assign popcount27_6cry_core_057 = ~input_a[19];
  assign popcount27_6cry_core_058 = input_a[20] | input_a[7];
  assign popcount27_6cry_core_059 = ~(input_a[17] & input_a[22]);
  assign popcount27_6cry_core_060 = input_a[5] | input_a[17];
  assign popcount27_6cry_core_061 = ~(input_a[4] & input_a[3]);
  assign popcount27_6cry_core_064 = ~(input_a[8] & input_a[1]);
  assign popcount27_6cry_core_065 = input_a[2] & input_a[6];
  assign popcount27_6cry_core_066 = input_a[11] ^ input_a[14];
  assign popcount27_6cry_core_067 = input_a[0] & input_a[16];
  assign popcount27_6cry_core_068 = input_a[24] ^ input_a[9];
  assign popcount27_6cry_core_069 = ~(input_a[19] | input_a[7]);
  assign popcount27_6cry_core_070 = ~input_a[2];
  assign popcount27_6cry_core_071 = ~(input_a[23] & input_a[15]);
  assign popcount27_6cry_core_072 = input_a[17] & input_a[24];
  assign popcount27_6cry_core_075 = input_a[13] & input_a[2];
  assign popcount27_6cry_core_076 = ~(input_a[22] | input_a[12]);
  assign popcount27_6cry_core_079 = input_a[9] ^ input_a[17];
  assign popcount27_6cry_core_080 = input_a[11] & input_a[24];
  assign popcount27_6cry_core_081 = input_a[23] ^ input_a[12];
  assign popcount27_6cry_core_082 = ~(input_a[22] | input_a[13]);
  assign popcount27_6cry_core_083 = input_a[19] & input_a[16];
  assign popcount27_6cry_core_084 = input_a[10] & input_a[15];
  assign popcount27_6cry_core_086 = ~(input_a[16] & input_a[5]);
  assign popcount27_6cry_core_087 = ~(input_a[21] | input_a[21]);
  assign popcount27_6cry_core_088 = ~(input_a[14] ^ input_a[17]);
  assign popcount27_6cry_core_090 = ~(input_a[7] ^ input_a[1]);
  assign popcount27_6cry_core_091 = ~input_a[7];
  assign popcount27_6cry_core_092 = ~(input_a[23] & input_a[18]);
  assign popcount27_6cry_core_093 = input_a[7] ^ input_a[23];
  assign popcount27_6cry_core_094 = ~(input_a[5] & input_a[20]);
  assign popcount27_6cry_core_096 = ~input_a[22];
  assign popcount27_6cry_core_099 = ~(input_a[8] & input_a[24]);
  assign popcount27_6cry_core_101 = input_a[3] ^ input_a[11];
  assign popcount27_6cry_core_104 = input_a[8] | input_a[13];
  assign popcount27_6cry_core_106 = input_a[18] ^ input_a[24];
  assign popcount27_6cry_core_107 = input_a[5] ^ input_a[16];
  assign popcount27_6cry_core_108 = ~input_a[6];
  assign popcount27_6cry_core_113 = input_a[16] & input_a[6];
  assign popcount27_6cry_core_114 = ~(input_a[24] | input_a[5]);
  assign popcount27_6cry_core_117 = ~input_a[10];
  assign popcount27_6cry_core_118 = input_a[10] ^ input_a[15];
  assign popcount27_6cry_core_119 = ~(input_a[20] | input_a[8]);
  assign popcount27_6cry_core_120 = ~(input_a[24] & input_a[18]);
  assign popcount27_6cry_core_121 = ~(input_a[3] & input_a[11]);
  assign popcount27_6cry_core_123 = ~(input_a[3] | input_a[12]);
  assign popcount27_6cry_core_126 = input_a[3] & input_a[5];
  assign popcount27_6cry_core_127 = ~(input_a[18] & input_a[4]);
  assign popcount27_6cry_core_128 = ~input_a[25];
  assign popcount27_6cry_core_130 = ~(input_a[12] & input_a[13]);
  assign popcount27_6cry_core_131 = ~(input_a[23] ^ input_a[15]);
  assign popcount27_6cry_core_133 = ~(input_a[4] | input_a[5]);
  assign popcount27_6cry_core_136 = input_a[13] ^ input_a[25];
  assign popcount27_6cry_core_137 = input_a[25] ^ input_a[26];
  assign popcount27_6cry_core_139 = ~(input_a[11] & input_a[14]);
  assign popcount27_6cry_core_140 = ~(input_a[19] & input_a[2]);
  assign popcount27_6cry_core_142 = ~input_a[13];
  assign popcount27_6cry_core_144 = input_a[3] | input_a[18];
  assign popcount27_6cry_core_146 = input_a[12] ^ input_a[11];
  assign popcount27_6cry_core_147 = input_a[9] ^ input_a[4];
  assign popcount27_6cry_core_148 = input_a[14] | input_a[19];
  assign popcount27_6cry_core_149 = ~(input_a[16] | input_a[6]);
  assign popcount27_6cry_core_154 = ~input_a[1];
  assign popcount27_6cry_core_156 = ~(input_a[2] ^ input_a[15]);
  assign popcount27_6cry_core_157 = ~(input_a[10] | input_a[8]);
  assign popcount27_6cry_core_158 = ~(input_a[18] & input_a[26]);
  assign popcount27_6cry_core_161 = ~(input_a[23] & input_a[6]);
  assign popcount27_6cry_core_162 = ~input_a[5];
  assign popcount27_6cry_core_163 = ~(input_a[13] ^ input_a[2]);
  assign popcount27_6cry_core_165 = input_a[4] & input_a[23];
  assign popcount27_6cry_core_167 = ~(input_a[6] & input_a[9]);
  assign popcount27_6cry_core_168 = ~(input_a[6] ^ input_a[20]);
  assign popcount27_6cry_core_169 = ~(input_a[15] & input_a[14]);
  assign popcount27_6cry_core_170 = ~(input_a[6] ^ input_a[7]);
  assign popcount27_6cry_core_171 = ~input_a[23];
  assign popcount27_6cry_core_172 = input_a[19] & input_a[5];
  assign popcount27_6cry_core_175 = ~(input_a[20] | input_a[10]);
  assign popcount27_6cry_core_176 = ~(input_a[17] ^ input_a[0]);
  assign popcount27_6cry_core_177 = ~input_a[3];
  assign popcount27_6cry_core_179 = ~(input_a[7] & input_a[3]);
  assign popcount27_6cry_core_182 = ~(input_a[10] | input_a[23]);
  assign popcount27_6cry_core_183 = ~(input_a[24] ^ input_a[3]);
  assign popcount27_6cry_core_186 = input_a[24] ^ input_a[22];
  assign popcount27_6cry_core_187 = ~(input_a[11] & input_a[4]);
  assign popcount27_6cry_core_188 = input_a[15] | input_a[5];
  assign popcount27_6cry_core_190 = ~(input_a[2] ^ input_a[13]);
  assign popcount27_6cry_core_192 = ~(input_a[14] ^ input_a[18]);
  assign popcount27_6cry_core_193 = ~input_a[4];
  assign popcount27_6cry_core_194 = input_a[11] | input_a[21];
  assign popcount27_6cry_core_195 = ~(input_a[11] ^ input_a[12]);

  assign popcount27_6cry_out[0] = 1'b1;
  assign popcount27_6cry_out[1] = input_a[26];
  assign popcount27_6cry_out[2] = 1'b0;
  assign popcount27_6cry_out[3] = input_a[14];
  assign popcount27_6cry_out[4] = 1'b0;
endmodule