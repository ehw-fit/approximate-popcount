// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.16973
// WCE=14.0
// EP=0.856089%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_n43g(input [24:0] input_a, output [4:0] popcount25_n43g_out);
  wire popcount25_n43g_core_027;
  wire popcount25_n43g_core_028;
  wire popcount25_n43g_core_029;
  wire popcount25_n43g_core_030;
  wire popcount25_n43g_core_031;
  wire popcount25_n43g_core_032;
  wire popcount25_n43g_core_033;
  wire popcount25_n43g_core_035;
  wire popcount25_n43g_core_038;
  wire popcount25_n43g_core_041;
  wire popcount25_n43g_core_046;
  wire popcount25_n43g_core_047;
  wire popcount25_n43g_core_049;
  wire popcount25_n43g_core_050;
  wire popcount25_n43g_core_051;
  wire popcount25_n43g_core_054;
  wire popcount25_n43g_core_055;
  wire popcount25_n43g_core_057;
  wire popcount25_n43g_core_058;
  wire popcount25_n43g_core_059;
  wire popcount25_n43g_core_060;
  wire popcount25_n43g_core_061;
  wire popcount25_n43g_core_062;
  wire popcount25_n43g_core_064;
  wire popcount25_n43g_core_066;
  wire popcount25_n43g_core_067;
  wire popcount25_n43g_core_068;
  wire popcount25_n43g_core_071_not;
  wire popcount25_n43g_core_072;
  wire popcount25_n43g_core_073;
  wire popcount25_n43g_core_074;
  wire popcount25_n43g_core_076;
  wire popcount25_n43g_core_077;
  wire popcount25_n43g_core_078;
  wire popcount25_n43g_core_079;
  wire popcount25_n43g_core_080;
  wire popcount25_n43g_core_081;
  wire popcount25_n43g_core_086;
  wire popcount25_n43g_core_087;
  wire popcount25_n43g_core_088;
  wire popcount25_n43g_core_089;
  wire popcount25_n43g_core_090;
  wire popcount25_n43g_core_091;
  wire popcount25_n43g_core_092;
  wire popcount25_n43g_core_098;
  wire popcount25_n43g_core_099;
  wire popcount25_n43g_core_100;
  wire popcount25_n43g_core_101;
  wire popcount25_n43g_core_102;
  wire popcount25_n43g_core_104;
  wire popcount25_n43g_core_105;
  wire popcount25_n43g_core_106;
  wire popcount25_n43g_core_107;
  wire popcount25_n43g_core_108;
  wire popcount25_n43g_core_109;
  wire popcount25_n43g_core_110;
  wire popcount25_n43g_core_111;
  wire popcount25_n43g_core_112;
  wire popcount25_n43g_core_113_not;
  wire popcount25_n43g_core_114;
  wire popcount25_n43g_core_115;
  wire popcount25_n43g_core_116;
  wire popcount25_n43g_core_117;
  wire popcount25_n43g_core_118;
  wire popcount25_n43g_core_119;
  wire popcount25_n43g_core_120;
  wire popcount25_n43g_core_122;
  wire popcount25_n43g_core_123;
  wire popcount25_n43g_core_126;
  wire popcount25_n43g_core_129;
  wire popcount25_n43g_core_131_not;
  wire popcount25_n43g_core_133;
  wire popcount25_n43g_core_134;
  wire popcount25_n43g_core_136;
  wire popcount25_n43g_core_137;
  wire popcount25_n43g_core_139;
  wire popcount25_n43g_core_140;
  wire popcount25_n43g_core_142;
  wire popcount25_n43g_core_144;
  wire popcount25_n43g_core_148;
  wire popcount25_n43g_core_150;
  wire popcount25_n43g_core_151;
  wire popcount25_n43g_core_152;
  wire popcount25_n43g_core_153;
  wire popcount25_n43g_core_154;
  wire popcount25_n43g_core_157;
  wire popcount25_n43g_core_158;
  wire popcount25_n43g_core_162;
  wire popcount25_n43g_core_163;
  wire popcount25_n43g_core_164;
  wire popcount25_n43g_core_165;
  wire popcount25_n43g_core_166;
  wire popcount25_n43g_core_168;
  wire popcount25_n43g_core_170;
  wire popcount25_n43g_core_172;
  wire popcount25_n43g_core_173;
  wire popcount25_n43g_core_175;
  wire popcount25_n43g_core_176;
  wire popcount25_n43g_core_178;
  wire popcount25_n43g_core_179;
  wire popcount25_n43g_core_181;
  wire popcount25_n43g_core_183;

  assign popcount25_n43g_core_027 = input_a[4] | input_a[24];
  assign popcount25_n43g_core_028 = ~(input_a[1] | input_a[24]);
  assign popcount25_n43g_core_029 = ~(input_a[13] ^ input_a[0]);
  assign popcount25_n43g_core_030 = ~(input_a[11] ^ input_a[18]);
  assign popcount25_n43g_core_031 = ~input_a[22];
  assign popcount25_n43g_core_032 = ~(input_a[16] & input_a[17]);
  assign popcount25_n43g_core_033 = input_a[23] | input_a[23];
  assign popcount25_n43g_core_035 = input_a[22] & input_a[5];
  assign popcount25_n43g_core_038 = ~(input_a[16] ^ input_a[7]);
  assign popcount25_n43g_core_041 = ~(input_a[2] ^ input_a[8]);
  assign popcount25_n43g_core_046 = ~(input_a[16] | input_a[12]);
  assign popcount25_n43g_core_047 = ~input_a[1];
  assign popcount25_n43g_core_049 = input_a[6] ^ input_a[8];
  assign popcount25_n43g_core_050 = input_a[18] & input_a[24];
  assign popcount25_n43g_core_051 = ~input_a[4];
  assign popcount25_n43g_core_054 = ~input_a[19];
  assign popcount25_n43g_core_055 = ~(input_a[4] | input_a[13]);
  assign popcount25_n43g_core_057 = input_a[15] & input_a[13];
  assign popcount25_n43g_core_058 = input_a[13] | input_a[6];
  assign popcount25_n43g_core_059 = input_a[0] | input_a[12];
  assign popcount25_n43g_core_060 = ~(input_a[4] | input_a[8]);
  assign popcount25_n43g_core_061 = input_a[18] ^ input_a[15];
  assign popcount25_n43g_core_062 = input_a[24] ^ input_a[18];
  assign popcount25_n43g_core_064 = ~input_a[9];
  assign popcount25_n43g_core_066 = ~(input_a[12] & input_a[1]);
  assign popcount25_n43g_core_067 = input_a[15] & input_a[7];
  assign popcount25_n43g_core_068 = input_a[9] | input_a[13];
  assign popcount25_n43g_core_071_not = ~input_a[2];
  assign popcount25_n43g_core_072 = ~input_a[14];
  assign popcount25_n43g_core_073 = ~(input_a[23] ^ input_a[13]);
  assign popcount25_n43g_core_074 = input_a[19] ^ input_a[19];
  assign popcount25_n43g_core_076 = ~(input_a[24] & input_a[1]);
  assign popcount25_n43g_core_077 = input_a[4] ^ input_a[16];
  assign popcount25_n43g_core_078 = ~(input_a[0] ^ input_a[6]);
  assign popcount25_n43g_core_079 = ~(input_a[23] & input_a[13]);
  assign popcount25_n43g_core_080 = input_a[15] | input_a[9];
  assign popcount25_n43g_core_081 = input_a[10] ^ input_a[24];
  assign popcount25_n43g_core_086 = ~input_a[14];
  assign popcount25_n43g_core_087 = input_a[12] | input_a[22];
  assign popcount25_n43g_core_088 = input_a[5] ^ input_a[14];
  assign popcount25_n43g_core_089 = input_a[12] ^ input_a[3];
  assign popcount25_n43g_core_090 = ~(input_a[1] ^ input_a[5]);
  assign popcount25_n43g_core_091 = input_a[0] | input_a[19];
  assign popcount25_n43g_core_092 = ~input_a[10];
  assign popcount25_n43g_core_098 = input_a[19] ^ input_a[22];
  assign popcount25_n43g_core_099 = ~(input_a[14] | input_a[8]);
  assign popcount25_n43g_core_100 = ~(input_a[20] ^ input_a[23]);
  assign popcount25_n43g_core_101 = ~(input_a[3] ^ input_a[11]);
  assign popcount25_n43g_core_102 = input_a[4] | input_a[3];
  assign popcount25_n43g_core_104 = ~(input_a[15] & input_a[6]);
  assign popcount25_n43g_core_105 = input_a[12] ^ input_a[19];
  assign popcount25_n43g_core_106 = ~(input_a[8] ^ input_a[15]);
  assign popcount25_n43g_core_107 = ~(input_a[4] | input_a[1]);
  assign popcount25_n43g_core_108 = input_a[3] ^ input_a[17];
  assign popcount25_n43g_core_109 = ~(input_a[15] & input_a[5]);
  assign popcount25_n43g_core_110 = input_a[9] & input_a[23];
  assign popcount25_n43g_core_111 = input_a[11] ^ input_a[16];
  assign popcount25_n43g_core_112 = ~input_a[8];
  assign popcount25_n43g_core_113_not = ~input_a[11];
  assign popcount25_n43g_core_114 = input_a[11] ^ input_a[14];
  assign popcount25_n43g_core_115 = input_a[20] ^ input_a[13];
  assign popcount25_n43g_core_116 = input_a[11] ^ input_a[15];
  assign popcount25_n43g_core_117 = ~(input_a[8] | input_a[3]);
  assign popcount25_n43g_core_118 = input_a[10] ^ input_a[15];
  assign popcount25_n43g_core_119 = ~input_a[19];
  assign popcount25_n43g_core_120 = input_a[0] | input_a[24];
  assign popcount25_n43g_core_122 = ~input_a[16];
  assign popcount25_n43g_core_123 = input_a[11] & input_a[2];
  assign popcount25_n43g_core_126 = ~(input_a[24] & input_a[19]);
  assign popcount25_n43g_core_129 = ~(input_a[5] | input_a[20]);
  assign popcount25_n43g_core_131_not = ~input_a[0];
  assign popcount25_n43g_core_133 = ~(input_a[12] & input_a[20]);
  assign popcount25_n43g_core_134 = ~input_a[17];
  assign popcount25_n43g_core_136 = ~(input_a[22] & input_a[22]);
  assign popcount25_n43g_core_137 = input_a[1] ^ input_a[6];
  assign popcount25_n43g_core_139 = ~input_a[14];
  assign popcount25_n43g_core_140 = ~input_a[12];
  assign popcount25_n43g_core_142 = ~(input_a[2] | input_a[19]);
  assign popcount25_n43g_core_144 = ~(input_a[8] | input_a[18]);
  assign popcount25_n43g_core_148 = input_a[19] ^ input_a[4];
  assign popcount25_n43g_core_150 = ~(input_a[21] & input_a[19]);
  assign popcount25_n43g_core_151 = input_a[18] ^ input_a[16];
  assign popcount25_n43g_core_152 = ~(input_a[17] & input_a[6]);
  assign popcount25_n43g_core_153 = ~input_a[23];
  assign popcount25_n43g_core_154 = ~(input_a[7] & input_a[17]);
  assign popcount25_n43g_core_157 = input_a[2] ^ input_a[9];
  assign popcount25_n43g_core_158 = input_a[12] | input_a[6];
  assign popcount25_n43g_core_162 = ~(input_a[3] | input_a[7]);
  assign popcount25_n43g_core_163 = input_a[14] | input_a[24];
  assign popcount25_n43g_core_164 = ~input_a[13];
  assign popcount25_n43g_core_165 = ~(input_a[15] ^ input_a[6]);
  assign popcount25_n43g_core_166 = ~input_a[5];
  assign popcount25_n43g_core_168 = ~input_a[23];
  assign popcount25_n43g_core_170 = input_a[12] | input_a[13];
  assign popcount25_n43g_core_172 = input_a[11] & input_a[17];
  assign popcount25_n43g_core_173 = ~(input_a[22] & input_a[15]);
  assign popcount25_n43g_core_175 = ~(input_a[10] ^ input_a[21]);
  assign popcount25_n43g_core_176 = ~(input_a[8] & input_a[0]);
  assign popcount25_n43g_core_178 = input_a[8] & input_a[9];
  assign popcount25_n43g_core_179 = ~(input_a[1] ^ input_a[14]);
  assign popcount25_n43g_core_181 = ~input_a[22];
  assign popcount25_n43g_core_183 = ~(input_a[7] & input_a[18]);

  assign popcount25_n43g_out[0] = 1'b0;
  assign popcount25_n43g_out[1] = input_a[3];
  assign popcount25_n43g_out[2] = 1'b1;
  assign popcount25_n43g_out[3] = 1'b1;
  assign popcount25_n43g_out[4] = 1'b0;
endmodule