// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5032
// WCE=42.0
// EP=0.998396%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_v8o5(input [38:0] input_a, output [5:0] popcount39_v8o5_out);
  wire popcount39_v8o5_core_041_not;
  wire popcount39_v8o5_core_042;
  wire popcount39_v8o5_core_043;
  wire popcount39_v8o5_core_045;
  wire popcount39_v8o5_core_046;
  wire popcount39_v8o5_core_048;
  wire popcount39_v8o5_core_054;
  wire popcount39_v8o5_core_055;
  wire popcount39_v8o5_core_056;
  wire popcount39_v8o5_core_057;
  wire popcount39_v8o5_core_058;
  wire popcount39_v8o5_core_059;
  wire popcount39_v8o5_core_062;
  wire popcount39_v8o5_core_063;
  wire popcount39_v8o5_core_064;
  wire popcount39_v8o5_core_065;
  wire popcount39_v8o5_core_070;
  wire popcount39_v8o5_core_071;
  wire popcount39_v8o5_core_074;
  wire popcount39_v8o5_core_075;
  wire popcount39_v8o5_core_077;
  wire popcount39_v8o5_core_078;
  wire popcount39_v8o5_core_079;
  wire popcount39_v8o5_core_081;
  wire popcount39_v8o5_core_082;
  wire popcount39_v8o5_core_083;
  wire popcount39_v8o5_core_085;
  wire popcount39_v8o5_core_086;
  wire popcount39_v8o5_core_087;
  wire popcount39_v8o5_core_088;
  wire popcount39_v8o5_core_089;
  wire popcount39_v8o5_core_090;
  wire popcount39_v8o5_core_092;
  wire popcount39_v8o5_core_094;
  wire popcount39_v8o5_core_096;
  wire popcount39_v8o5_core_097;
  wire popcount39_v8o5_core_100;
  wire popcount39_v8o5_core_101;
  wire popcount39_v8o5_core_102;
  wire popcount39_v8o5_core_103;
  wire popcount39_v8o5_core_104;
  wire popcount39_v8o5_core_106;
  wire popcount39_v8o5_core_108;
  wire popcount39_v8o5_core_109;
  wire popcount39_v8o5_core_110;
  wire popcount39_v8o5_core_111;
  wire popcount39_v8o5_core_112;
  wire popcount39_v8o5_core_114;
  wire popcount39_v8o5_core_115;
  wire popcount39_v8o5_core_117;
  wire popcount39_v8o5_core_118;
  wire popcount39_v8o5_core_119;
  wire popcount39_v8o5_core_122;
  wire popcount39_v8o5_core_124;
  wire popcount39_v8o5_core_125;
  wire popcount39_v8o5_core_126;
  wire popcount39_v8o5_core_127;
  wire popcount39_v8o5_core_129;
  wire popcount39_v8o5_core_131;
  wire popcount39_v8o5_core_132;
  wire popcount39_v8o5_core_133;
  wire popcount39_v8o5_core_136;
  wire popcount39_v8o5_core_137;
  wire popcount39_v8o5_core_138;
  wire popcount39_v8o5_core_140;
  wire popcount39_v8o5_core_141;
  wire popcount39_v8o5_core_143;
  wire popcount39_v8o5_core_145;
  wire popcount39_v8o5_core_146;
  wire popcount39_v8o5_core_147;
  wire popcount39_v8o5_core_150_not;
  wire popcount39_v8o5_core_151;
  wire popcount39_v8o5_core_152;
  wire popcount39_v8o5_core_153;
  wire popcount39_v8o5_core_155;
  wire popcount39_v8o5_core_156;
  wire popcount39_v8o5_core_158;
  wire popcount39_v8o5_core_160;
  wire popcount39_v8o5_core_161;
  wire popcount39_v8o5_core_165;
  wire popcount39_v8o5_core_166;
  wire popcount39_v8o5_core_168;
  wire popcount39_v8o5_core_169;
  wire popcount39_v8o5_core_170;
  wire popcount39_v8o5_core_171;
  wire popcount39_v8o5_core_172;
  wire popcount39_v8o5_core_173;
  wire popcount39_v8o5_core_174;
  wire popcount39_v8o5_core_176;
  wire popcount39_v8o5_core_177;
  wire popcount39_v8o5_core_178;
  wire popcount39_v8o5_core_179;
  wire popcount39_v8o5_core_180;
  wire popcount39_v8o5_core_182;
  wire popcount39_v8o5_core_185;
  wire popcount39_v8o5_core_186;
  wire popcount39_v8o5_core_187_not;
  wire popcount39_v8o5_core_188;
  wire popcount39_v8o5_core_189;
  wire popcount39_v8o5_core_190;
  wire popcount39_v8o5_core_192;
  wire popcount39_v8o5_core_193;
  wire popcount39_v8o5_core_194;
  wire popcount39_v8o5_core_195;
  wire popcount39_v8o5_core_196;
  wire popcount39_v8o5_core_198;
  wire popcount39_v8o5_core_199;
  wire popcount39_v8o5_core_200;
  wire popcount39_v8o5_core_201;
  wire popcount39_v8o5_core_202;
  wire popcount39_v8o5_core_203;
  wire popcount39_v8o5_core_205;
  wire popcount39_v8o5_core_206;
  wire popcount39_v8o5_core_207;
  wire popcount39_v8o5_core_208;
  wire popcount39_v8o5_core_209;
  wire popcount39_v8o5_core_210;
  wire popcount39_v8o5_core_211;
  wire popcount39_v8o5_core_213;
  wire popcount39_v8o5_core_214;
  wire popcount39_v8o5_core_215;
  wire popcount39_v8o5_core_217;
  wire popcount39_v8o5_core_218;
  wire popcount39_v8o5_core_220;
  wire popcount39_v8o5_core_221;
  wire popcount39_v8o5_core_222;
  wire popcount39_v8o5_core_223;
  wire popcount39_v8o5_core_224;
  wire popcount39_v8o5_core_226;
  wire popcount39_v8o5_core_227;
  wire popcount39_v8o5_core_230;
  wire popcount39_v8o5_core_232;
  wire popcount39_v8o5_core_233;
  wire popcount39_v8o5_core_234;
  wire popcount39_v8o5_core_235;
  wire popcount39_v8o5_core_236;
  wire popcount39_v8o5_core_237;
  wire popcount39_v8o5_core_238;
  wire popcount39_v8o5_core_239;
  wire popcount39_v8o5_core_240;
  wire popcount39_v8o5_core_242;
  wire popcount39_v8o5_core_243;
  wire popcount39_v8o5_core_244;
  wire popcount39_v8o5_core_245;
  wire popcount39_v8o5_core_246;
  wire popcount39_v8o5_core_247;
  wire popcount39_v8o5_core_248;
  wire popcount39_v8o5_core_251;
  wire popcount39_v8o5_core_252;
  wire popcount39_v8o5_core_255;
  wire popcount39_v8o5_core_257;
  wire popcount39_v8o5_core_258;
  wire popcount39_v8o5_core_261;
  wire popcount39_v8o5_core_263;
  wire popcount39_v8o5_core_264;
  wire popcount39_v8o5_core_265;
  wire popcount39_v8o5_core_267;
  wire popcount39_v8o5_core_268;
  wire popcount39_v8o5_core_273;
  wire popcount39_v8o5_core_275;
  wire popcount39_v8o5_core_276;
  wire popcount39_v8o5_core_277;
  wire popcount39_v8o5_core_278;
  wire popcount39_v8o5_core_279;
  wire popcount39_v8o5_core_280;
  wire popcount39_v8o5_core_281;
  wire popcount39_v8o5_core_283;
  wire popcount39_v8o5_core_284_not;
  wire popcount39_v8o5_core_286;
  wire popcount39_v8o5_core_287;
  wire popcount39_v8o5_core_290;
  wire popcount39_v8o5_core_295;
  wire popcount39_v8o5_core_296;
  wire popcount39_v8o5_core_297;
  wire popcount39_v8o5_core_298;
  wire popcount39_v8o5_core_300;
  wire popcount39_v8o5_core_303;

  assign popcount39_v8o5_core_041_not = ~input_a[25];
  assign popcount39_v8o5_core_042 = input_a[34] | input_a[37];
  assign popcount39_v8o5_core_043 = input_a[15] | input_a[2];
  assign popcount39_v8o5_core_045 = input_a[21] | input_a[31];
  assign popcount39_v8o5_core_046 = ~(input_a[9] ^ input_a[9]);
  assign popcount39_v8o5_core_048 = ~input_a[4];
  assign popcount39_v8o5_core_054 = ~(input_a[11] ^ input_a[37]);
  assign popcount39_v8o5_core_055 = input_a[29] ^ input_a[37];
  assign popcount39_v8o5_core_056 = ~(input_a[25] | input_a[25]);
  assign popcount39_v8o5_core_057 = ~input_a[32];
  assign popcount39_v8o5_core_058 = ~(input_a[26] ^ input_a[36]);
  assign popcount39_v8o5_core_059 = ~(input_a[1] | input_a[6]);
  assign popcount39_v8o5_core_062 = ~input_a[14];
  assign popcount39_v8o5_core_063 = input_a[23] | input_a[7];
  assign popcount39_v8o5_core_064 = ~(input_a[11] ^ input_a[37]);
  assign popcount39_v8o5_core_065 = input_a[28] ^ input_a[4];
  assign popcount39_v8o5_core_070 = ~(input_a[2] | input_a[5]);
  assign popcount39_v8o5_core_071 = ~(input_a[11] | input_a[23]);
  assign popcount39_v8o5_core_074 = input_a[33] ^ input_a[10];
  assign popcount39_v8o5_core_075 = ~input_a[5];
  assign popcount39_v8o5_core_077 = input_a[2] | input_a[8];
  assign popcount39_v8o5_core_078 = ~input_a[7];
  assign popcount39_v8o5_core_079 = ~(input_a[24] | input_a[18]);
  assign popcount39_v8o5_core_081 = input_a[17] ^ input_a[17];
  assign popcount39_v8o5_core_082 = ~input_a[22];
  assign popcount39_v8o5_core_083 = input_a[28] | input_a[4];
  assign popcount39_v8o5_core_085 = ~(input_a[33] & input_a[23]);
  assign popcount39_v8o5_core_086 = ~(input_a[37] | input_a[12]);
  assign popcount39_v8o5_core_087 = ~(input_a[34] | input_a[16]);
  assign popcount39_v8o5_core_088 = ~(input_a[18] | input_a[27]);
  assign popcount39_v8o5_core_089 = input_a[21] ^ input_a[18];
  assign popcount39_v8o5_core_090 = ~(input_a[34] ^ input_a[30]);
  assign popcount39_v8o5_core_092 = ~(input_a[2] ^ input_a[34]);
  assign popcount39_v8o5_core_094 = ~(input_a[3] & input_a[2]);
  assign popcount39_v8o5_core_096 = ~input_a[4];
  assign popcount39_v8o5_core_097 = input_a[15] | input_a[26];
  assign popcount39_v8o5_core_100 = input_a[17] & input_a[35];
  assign popcount39_v8o5_core_101 = input_a[14] & input_a[23];
  assign popcount39_v8o5_core_102 = input_a[35] & input_a[30];
  assign popcount39_v8o5_core_103 = ~input_a[9];
  assign popcount39_v8o5_core_104 = input_a[8] | input_a[17];
  assign popcount39_v8o5_core_106 = ~(input_a[0] | input_a[7]);
  assign popcount39_v8o5_core_108 = input_a[28] | input_a[11];
  assign popcount39_v8o5_core_109 = ~input_a[31];
  assign popcount39_v8o5_core_110 = ~(input_a[30] & input_a[26]);
  assign popcount39_v8o5_core_111 = ~input_a[19];
  assign popcount39_v8o5_core_112 = ~(input_a[28] | input_a[37]);
  assign popcount39_v8o5_core_114 = ~(input_a[38] & input_a[37]);
  assign popcount39_v8o5_core_115 = ~(input_a[18] ^ input_a[22]);
  assign popcount39_v8o5_core_117 = ~(input_a[22] ^ input_a[1]);
  assign popcount39_v8o5_core_118 = input_a[9] | input_a[38];
  assign popcount39_v8o5_core_119 = ~input_a[34];
  assign popcount39_v8o5_core_122 = ~(input_a[11] & input_a[7]);
  assign popcount39_v8o5_core_124 = input_a[37] & input_a[17];
  assign popcount39_v8o5_core_125 = input_a[17] | input_a[31];
  assign popcount39_v8o5_core_126 = input_a[6] | input_a[1];
  assign popcount39_v8o5_core_127 = ~input_a[18];
  assign popcount39_v8o5_core_129 = input_a[19] & input_a[16];
  assign popcount39_v8o5_core_131 = input_a[15] & input_a[10];
  assign popcount39_v8o5_core_132 = ~(input_a[12] ^ input_a[27]);
  assign popcount39_v8o5_core_133 = ~(input_a[18] | input_a[28]);
  assign popcount39_v8o5_core_136 = ~(input_a[10] ^ input_a[8]);
  assign popcount39_v8o5_core_137 = input_a[2] ^ input_a[19];
  assign popcount39_v8o5_core_138 = ~(input_a[13] & input_a[11]);
  assign popcount39_v8o5_core_140 = input_a[10] | input_a[31];
  assign popcount39_v8o5_core_141 = ~(input_a[32] | input_a[18]);
  assign popcount39_v8o5_core_143 = ~input_a[2];
  assign popcount39_v8o5_core_145 = ~input_a[12];
  assign popcount39_v8o5_core_146 = input_a[37] ^ input_a[19];
  assign popcount39_v8o5_core_147 = ~(input_a[6] ^ input_a[4]);
  assign popcount39_v8o5_core_150_not = ~input_a[12];
  assign popcount39_v8o5_core_151 = ~(input_a[22] & input_a[22]);
  assign popcount39_v8o5_core_152 = ~(input_a[8] & input_a[1]);
  assign popcount39_v8o5_core_153 = input_a[6] ^ input_a[26];
  assign popcount39_v8o5_core_155 = ~(input_a[28] & input_a[12]);
  assign popcount39_v8o5_core_156 = ~input_a[21];
  assign popcount39_v8o5_core_158 = ~(input_a[15] | input_a[34]);
  assign popcount39_v8o5_core_160 = input_a[26] ^ input_a[32];
  assign popcount39_v8o5_core_161 = input_a[28] | input_a[26];
  assign popcount39_v8o5_core_165 = ~(input_a[12] | input_a[28]);
  assign popcount39_v8o5_core_166 = ~(input_a[12] | input_a[5]);
  assign popcount39_v8o5_core_168 = ~(input_a[28] ^ input_a[13]);
  assign popcount39_v8o5_core_169 = ~(input_a[36] | input_a[16]);
  assign popcount39_v8o5_core_170 = ~input_a[4];
  assign popcount39_v8o5_core_171 = input_a[17] ^ input_a[9];
  assign popcount39_v8o5_core_172 = input_a[33] & input_a[30];
  assign popcount39_v8o5_core_173 = ~(input_a[3] | input_a[0]);
  assign popcount39_v8o5_core_174 = input_a[36] & input_a[22];
  assign popcount39_v8o5_core_176 = ~(input_a[32] ^ input_a[16]);
  assign popcount39_v8o5_core_177 = ~input_a[29];
  assign popcount39_v8o5_core_178 = input_a[25] & input_a[36];
  assign popcount39_v8o5_core_179 = ~input_a[12];
  assign popcount39_v8o5_core_180 = ~(input_a[26] & input_a[19]);
  assign popcount39_v8o5_core_182 = ~(input_a[5] & input_a[26]);
  assign popcount39_v8o5_core_185 = ~(input_a[16] & input_a[23]);
  assign popcount39_v8o5_core_186 = ~input_a[15];
  assign popcount39_v8o5_core_187_not = ~input_a[21];
  assign popcount39_v8o5_core_188 = ~input_a[31];
  assign popcount39_v8o5_core_189 = ~(input_a[12] ^ input_a[36]);
  assign popcount39_v8o5_core_190 = ~input_a[4];
  assign popcount39_v8o5_core_192 = input_a[2] | input_a[22];
  assign popcount39_v8o5_core_193 = ~input_a[27];
  assign popcount39_v8o5_core_194 = ~(input_a[18] & input_a[37]);
  assign popcount39_v8o5_core_195 = ~(input_a[28] | input_a[19]);
  assign popcount39_v8o5_core_196 = input_a[36] & input_a[30];
  assign popcount39_v8o5_core_198 = input_a[27] | input_a[36];
  assign popcount39_v8o5_core_199 = ~input_a[32];
  assign popcount39_v8o5_core_200 = ~input_a[10];
  assign popcount39_v8o5_core_201 = input_a[25] & input_a[1];
  assign popcount39_v8o5_core_202 = ~(input_a[21] & input_a[18]);
  assign popcount39_v8o5_core_203 = input_a[37] & input_a[7];
  assign popcount39_v8o5_core_205 = ~input_a[28];
  assign popcount39_v8o5_core_206 = input_a[21] & input_a[21];
  assign popcount39_v8o5_core_207 = ~input_a[27];
  assign popcount39_v8o5_core_208 = ~input_a[31];
  assign popcount39_v8o5_core_209 = ~(input_a[2] & input_a[22]);
  assign popcount39_v8o5_core_210 = input_a[26] | input_a[4];
  assign popcount39_v8o5_core_211 = ~(input_a[31] ^ input_a[28]);
  assign popcount39_v8o5_core_213 = ~input_a[1];
  assign popcount39_v8o5_core_214 = input_a[6] & input_a[35];
  assign popcount39_v8o5_core_215 = input_a[33] & input_a[17];
  assign popcount39_v8o5_core_217 = ~(input_a[6] | input_a[22]);
  assign popcount39_v8o5_core_218 = input_a[1] & input_a[30];
  assign popcount39_v8o5_core_220 = ~input_a[23];
  assign popcount39_v8o5_core_221 = ~(input_a[3] & input_a[31]);
  assign popcount39_v8o5_core_222 = input_a[8] | input_a[7];
  assign popcount39_v8o5_core_223 = ~(input_a[9] ^ input_a[1]);
  assign popcount39_v8o5_core_224 = ~input_a[6];
  assign popcount39_v8o5_core_226 = ~input_a[12];
  assign popcount39_v8o5_core_227 = ~(input_a[15] | input_a[27]);
  assign popcount39_v8o5_core_230 = input_a[28] | input_a[8];
  assign popcount39_v8o5_core_232 = ~input_a[11];
  assign popcount39_v8o5_core_233 = input_a[18] | input_a[24];
  assign popcount39_v8o5_core_234 = ~input_a[15];
  assign popcount39_v8o5_core_235 = input_a[38] ^ input_a[7];
  assign popcount39_v8o5_core_236 = input_a[25] ^ input_a[22];
  assign popcount39_v8o5_core_237 = ~(input_a[10] & input_a[3]);
  assign popcount39_v8o5_core_238 = input_a[19] | input_a[16];
  assign popcount39_v8o5_core_239 = ~(input_a[10] ^ input_a[20]);
  assign popcount39_v8o5_core_240 = ~(input_a[37] ^ input_a[7]);
  assign popcount39_v8o5_core_242 = ~(input_a[16] ^ input_a[14]);
  assign popcount39_v8o5_core_243 = ~input_a[7];
  assign popcount39_v8o5_core_244 = input_a[6] | input_a[34];
  assign popcount39_v8o5_core_245 = input_a[15] ^ input_a[35];
  assign popcount39_v8o5_core_246 = ~input_a[3];
  assign popcount39_v8o5_core_247 = input_a[1] ^ input_a[22];
  assign popcount39_v8o5_core_248 = input_a[1] & input_a[10];
  assign popcount39_v8o5_core_251 = ~(input_a[30] ^ input_a[19]);
  assign popcount39_v8o5_core_252 = ~input_a[20];
  assign popcount39_v8o5_core_255 = ~input_a[22];
  assign popcount39_v8o5_core_257 = ~(input_a[16] & input_a[2]);
  assign popcount39_v8o5_core_258 = ~(input_a[17] ^ input_a[4]);
  assign popcount39_v8o5_core_261 = ~(input_a[2] & input_a[5]);
  assign popcount39_v8o5_core_263 = input_a[32] | input_a[32];
  assign popcount39_v8o5_core_264 = input_a[36] | input_a[32];
  assign popcount39_v8o5_core_265 = ~(input_a[6] | input_a[12]);
  assign popcount39_v8o5_core_267 = input_a[8] | input_a[18];
  assign popcount39_v8o5_core_268 = ~(input_a[31] ^ input_a[3]);
  assign popcount39_v8o5_core_273 = ~(input_a[8] ^ input_a[14]);
  assign popcount39_v8o5_core_275 = ~(input_a[1] ^ input_a[29]);
  assign popcount39_v8o5_core_276 = ~input_a[4];
  assign popcount39_v8o5_core_277 = input_a[6] | input_a[4];
  assign popcount39_v8o5_core_278 = ~input_a[28];
  assign popcount39_v8o5_core_279 = input_a[6] & input_a[23];
  assign popcount39_v8o5_core_280 = input_a[2] ^ input_a[32];
  assign popcount39_v8o5_core_281 = ~(input_a[14] & input_a[32]);
  assign popcount39_v8o5_core_283 = ~(input_a[3] & input_a[4]);
  assign popcount39_v8o5_core_284_not = ~input_a[5];
  assign popcount39_v8o5_core_286 = input_a[32] & input_a[16];
  assign popcount39_v8o5_core_287 = input_a[16] ^ input_a[4];
  assign popcount39_v8o5_core_290 = input_a[20] ^ input_a[15];
  assign popcount39_v8o5_core_295 = ~(input_a[11] ^ input_a[1]);
  assign popcount39_v8o5_core_296 = input_a[10] ^ input_a[25];
  assign popcount39_v8o5_core_297 = input_a[13] ^ input_a[37];
  assign popcount39_v8o5_core_298 = input_a[33] ^ input_a[15];
  assign popcount39_v8o5_core_300 = input_a[31] | input_a[13];
  assign popcount39_v8o5_core_303 = ~input_a[4];

  assign popcount39_v8o5_out[0] = input_a[34];
  assign popcount39_v8o5_out[1] = input_a[1];
  assign popcount39_v8o5_out[2] = input_a[0];
  assign popcount39_v8o5_out[3] = input_a[17];
  assign popcount39_v8o5_out[4] = 1'b0;
  assign popcount39_v8o5_out[5] = input_a[20];
endmodule