// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.20746
// WCE=18.0
// EP=0.902659%
// Printed PDK parameters:
//  Area=53903702.0
//  Delay=71612168.0
//  Power=2573200.0

module popcount35_g3qe(input [34:0] input_a, output [5:0] popcount35_g3qe_out);
  wire popcount35_g3qe_core_037;
  wire popcount35_g3qe_core_038;
  wire popcount35_g3qe_core_039;
  wire popcount35_g3qe_core_040;
  wire popcount35_g3qe_core_042;
  wire popcount35_g3qe_core_043;
  wire popcount35_g3qe_core_044;
  wire popcount35_g3qe_core_045;
  wire popcount35_g3qe_core_049;
  wire popcount35_g3qe_core_051;
  wire popcount35_g3qe_core_052;
  wire popcount35_g3qe_core_053;
  wire popcount35_g3qe_core_054;
  wire popcount35_g3qe_core_055;
  wire popcount35_g3qe_core_056;
  wire popcount35_g3qe_core_057;
  wire popcount35_g3qe_core_060;
  wire popcount35_g3qe_core_061;
  wire popcount35_g3qe_core_062;
  wire popcount35_g3qe_core_063;
  wire popcount35_g3qe_core_064;
  wire popcount35_g3qe_core_065;
  wire popcount35_g3qe_core_066;
  wire popcount35_g3qe_core_067;
  wire popcount35_g3qe_core_068;
  wire popcount35_g3qe_core_069;
  wire popcount35_g3qe_core_070;
  wire popcount35_g3qe_core_071;
  wire popcount35_g3qe_core_072;
  wire popcount35_g3qe_core_073;
  wire popcount35_g3qe_core_074;
  wire popcount35_g3qe_core_078;
  wire popcount35_g3qe_core_081;
  wire popcount35_g3qe_core_082;
  wire popcount35_g3qe_core_085;
  wire popcount35_g3qe_core_087;
  wire popcount35_g3qe_core_088;
  wire popcount35_g3qe_core_089;
  wire popcount35_g3qe_core_091;
  wire popcount35_g3qe_core_092;
  wire popcount35_g3qe_core_093;
  wire popcount35_g3qe_core_094;
  wire popcount35_g3qe_core_095;
  wire popcount35_g3qe_core_096;
  wire popcount35_g3qe_core_097;
  wire popcount35_g3qe_core_101_not;
  wire popcount35_g3qe_core_106;
  wire popcount35_g3qe_core_107;
  wire popcount35_g3qe_core_108;
  wire popcount35_g3qe_core_109;
  wire popcount35_g3qe_core_110;
  wire popcount35_g3qe_core_113_not;
  wire popcount35_g3qe_core_115;
  wire popcount35_g3qe_core_117;
  wire popcount35_g3qe_core_118;
  wire popcount35_g3qe_core_119;
  wire popcount35_g3qe_core_120;
  wire popcount35_g3qe_core_121;
  wire popcount35_g3qe_core_123;
  wire popcount35_g3qe_core_125;
  wire popcount35_g3qe_core_126;
  wire popcount35_g3qe_core_127;
  wire popcount35_g3qe_core_128;
  wire popcount35_g3qe_core_129;
  wire popcount35_g3qe_core_131;
  wire popcount35_g3qe_core_134;
  wire popcount35_g3qe_core_135;
  wire popcount35_g3qe_core_136;
  wire popcount35_g3qe_core_137;
  wire popcount35_g3qe_core_139;
  wire popcount35_g3qe_core_141;
  wire popcount35_g3qe_core_143;
  wire popcount35_g3qe_core_144;
  wire popcount35_g3qe_core_145;
  wire popcount35_g3qe_core_146;
  wire popcount35_g3qe_core_149;
  wire popcount35_g3qe_core_151;
  wire popcount35_g3qe_core_153;
  wire popcount35_g3qe_core_154;
  wire popcount35_g3qe_core_155;
  wire popcount35_g3qe_core_156;
  wire popcount35_g3qe_core_157;
  wire popcount35_g3qe_core_158;
  wire popcount35_g3qe_core_162;
  wire popcount35_g3qe_core_164;
  wire popcount35_g3qe_core_170;
  wire popcount35_g3qe_core_174;
  wire popcount35_g3qe_core_177;
  wire popcount35_g3qe_core_178;
  wire popcount35_g3qe_core_180;
  wire popcount35_g3qe_core_185;
  wire popcount35_g3qe_core_187;
  wire popcount35_g3qe_core_188;
  wire popcount35_g3qe_core_193;
  wire popcount35_g3qe_core_195;
  wire popcount35_g3qe_core_196;
  wire popcount35_g3qe_core_199;
  wire popcount35_g3qe_core_200;
  wire popcount35_g3qe_core_202;
  wire popcount35_g3qe_core_203;
  wire popcount35_g3qe_core_204;
  wire popcount35_g3qe_core_205;
  wire popcount35_g3qe_core_206;
  wire popcount35_g3qe_core_207;
  wire popcount35_g3qe_core_208;
  wire popcount35_g3qe_core_211;
  wire popcount35_g3qe_core_212;
  wire popcount35_g3qe_core_215;
  wire popcount35_g3qe_core_217;
  wire popcount35_g3qe_core_218;
  wire popcount35_g3qe_core_219;
  wire popcount35_g3qe_core_220;
  wire popcount35_g3qe_core_221;
  wire popcount35_g3qe_core_222;
  wire popcount35_g3qe_core_223;
  wire popcount35_g3qe_core_224;
  wire popcount35_g3qe_core_225;
  wire popcount35_g3qe_core_226;
  wire popcount35_g3qe_core_227;
  wire popcount35_g3qe_core_230;
  wire popcount35_g3qe_core_234;
  wire popcount35_g3qe_core_237;
  wire popcount35_g3qe_core_238;
  wire popcount35_g3qe_core_239;
  wire popcount35_g3qe_core_240;
  wire popcount35_g3qe_core_241;
  wire popcount35_g3qe_core_242;
  wire popcount35_g3qe_core_243;
  wire popcount35_g3qe_core_244;
  wire popcount35_g3qe_core_245;
  wire popcount35_g3qe_core_246;
  wire popcount35_g3qe_core_247;
  wire popcount35_g3qe_core_248;
  wire popcount35_g3qe_core_249;
  wire popcount35_g3qe_core_250;
  wire popcount35_g3qe_core_251;
  wire popcount35_g3qe_core_252;
  wire popcount35_g3qe_core_253;
  wire popcount35_g3qe_core_254;
  wire popcount35_g3qe_core_257;
  wire popcount35_g3qe_core_258;
  wire popcount35_g3qe_core_261;
  wire popcount35_g3qe_core_263;
  wire popcount35_g3qe_core_264;

  assign popcount35_g3qe_core_037 = input_a[31] ^ input_a[18];
  assign popcount35_g3qe_core_038 = input_a[26] & input_a[24];
  assign popcount35_g3qe_core_039 = input_a[2] ^ input_a[3];
  assign popcount35_g3qe_core_040 = input_a[2] & input_a[3];
  assign popcount35_g3qe_core_042 = input_a[25] & popcount35_g3qe_core_039;
  assign popcount35_g3qe_core_043 = popcount35_g3qe_core_038 ^ popcount35_g3qe_core_040;
  assign popcount35_g3qe_core_044 = popcount35_g3qe_core_038 & popcount35_g3qe_core_040;
  assign popcount35_g3qe_core_045 = popcount35_g3qe_core_043 | popcount35_g3qe_core_042;
  assign popcount35_g3qe_core_049 = input_a[32] & input_a[5];
  assign popcount35_g3qe_core_051 = input_a[19] & input_a[5];
  assign popcount35_g3qe_core_052 = ~input_a[21];
  assign popcount35_g3qe_core_053 = input_a[5] & input_a[18];
  assign popcount35_g3qe_core_054 = popcount35_g3qe_core_049 ^ popcount35_g3qe_core_051;
  assign popcount35_g3qe_core_055 = popcount35_g3qe_core_049 & popcount35_g3qe_core_051;
  assign popcount35_g3qe_core_056 = popcount35_g3qe_core_054 | popcount35_g3qe_core_053;
  assign popcount35_g3qe_core_057 = ~input_a[11];
  assign popcount35_g3qe_core_060 = input_a[8] & input_a[20];
  assign popcount35_g3qe_core_061 = popcount35_g3qe_core_045 ^ popcount35_g3qe_core_056;
  assign popcount35_g3qe_core_062 = popcount35_g3qe_core_045 & popcount35_g3qe_core_056;
  assign popcount35_g3qe_core_063 = popcount35_g3qe_core_061 ^ popcount35_g3qe_core_060;
  assign popcount35_g3qe_core_064 = popcount35_g3qe_core_061 & popcount35_g3qe_core_060;
  assign popcount35_g3qe_core_065 = popcount35_g3qe_core_062 | popcount35_g3qe_core_064;
  assign popcount35_g3qe_core_066 = popcount35_g3qe_core_044 ^ popcount35_g3qe_core_055;
  assign popcount35_g3qe_core_067 = popcount35_g3qe_core_044 & popcount35_g3qe_core_055;
  assign popcount35_g3qe_core_068 = popcount35_g3qe_core_066 ^ popcount35_g3qe_core_065;
  assign popcount35_g3qe_core_069 = popcount35_g3qe_core_066 & popcount35_g3qe_core_065;
  assign popcount35_g3qe_core_070 = popcount35_g3qe_core_067 | popcount35_g3qe_core_069;
  assign popcount35_g3qe_core_071 = ~(input_a[12] | input_a[6]);
  assign popcount35_g3qe_core_072 = input_a[7] & input_a[21];
  assign popcount35_g3qe_core_073 = ~input_a[32];
  assign popcount35_g3qe_core_074 = input_a[33] & input_a[11];
  assign popcount35_g3qe_core_078 = input_a[33] & popcount35_g3qe_core_074;
  assign popcount35_g3qe_core_081 = popcount35_g3qe_core_078 | popcount35_g3qe_core_072;
  assign popcount35_g3qe_core_082 = ~input_a[4];
  assign popcount35_g3qe_core_085 = input_a[15] & input_a[16];
  assign popcount35_g3qe_core_087 = input_a[14] & input_a[1];
  assign popcount35_g3qe_core_088 = popcount35_g3qe_core_085 | popcount35_g3qe_core_087;
  assign popcount35_g3qe_core_089 = popcount35_g3qe_core_085 & popcount35_g3qe_core_087;
  assign popcount35_g3qe_core_091 = input_a[34] & input_a[28];
  assign popcount35_g3qe_core_092 = input_a[12] ^ popcount35_g3qe_core_088;
  assign popcount35_g3qe_core_093 = input_a[12] & popcount35_g3qe_core_088;
  assign popcount35_g3qe_core_094 = popcount35_g3qe_core_092 ^ popcount35_g3qe_core_091;
  assign popcount35_g3qe_core_095 = popcount35_g3qe_core_092 & popcount35_g3qe_core_091;
  assign popcount35_g3qe_core_096 = popcount35_g3qe_core_093 | popcount35_g3qe_core_095;
  assign popcount35_g3qe_core_097 = popcount35_g3qe_core_089 | popcount35_g3qe_core_096;
  assign popcount35_g3qe_core_101_not = ~popcount35_g3qe_core_094;
  assign popcount35_g3qe_core_106 = popcount35_g3qe_core_081 ^ popcount35_g3qe_core_097;
  assign popcount35_g3qe_core_107 = popcount35_g3qe_core_081 & popcount35_g3qe_core_097;
  assign popcount35_g3qe_core_108 = popcount35_g3qe_core_106 ^ popcount35_g3qe_core_094;
  assign popcount35_g3qe_core_109 = popcount35_g3qe_core_106 & popcount35_g3qe_core_094;
  assign popcount35_g3qe_core_110 = popcount35_g3qe_core_107 | popcount35_g3qe_core_109;
  assign popcount35_g3qe_core_113_not = ~input_a[29];
  assign popcount35_g3qe_core_115 = popcount35_g3qe_core_063 ^ popcount35_g3qe_core_101_not;
  assign popcount35_g3qe_core_117 = popcount35_g3qe_core_115 ^ input_a[29];
  assign popcount35_g3qe_core_118 = input_a[4] | input_a[31];
  assign popcount35_g3qe_core_119 = input_a[6] ^ input_a[32];
  assign popcount35_g3qe_core_120 = popcount35_g3qe_core_068 ^ popcount35_g3qe_core_108;
  assign popcount35_g3qe_core_121 = popcount35_g3qe_core_068 & popcount35_g3qe_core_108;
  assign popcount35_g3qe_core_123 = ~(input_a[32] | input_a[32]);
  assign popcount35_g3qe_core_125 = popcount35_g3qe_core_070 ^ popcount35_g3qe_core_110;
  assign popcount35_g3qe_core_126 = popcount35_g3qe_core_070 & popcount35_g3qe_core_110;
  assign popcount35_g3qe_core_127 = popcount35_g3qe_core_125 ^ popcount35_g3qe_core_121;
  assign popcount35_g3qe_core_128 = popcount35_g3qe_core_125 & popcount35_g3qe_core_121;
  assign popcount35_g3qe_core_129 = popcount35_g3qe_core_126 | popcount35_g3qe_core_128;
  assign popcount35_g3qe_core_131 = input_a[22] & input_a[9];
  assign popcount35_g3qe_core_134 = ~(input_a[17] & input_a[29]);
  assign popcount35_g3qe_core_135 = input_a[30] & input_a[10];
  assign popcount35_g3qe_core_136 = ~input_a[8];
  assign popcount35_g3qe_core_137 = ~input_a[6];
  assign popcount35_g3qe_core_139 = ~input_a[23];
  assign popcount35_g3qe_core_141 = input_a[30] & input_a[34];
  assign popcount35_g3qe_core_143 = ~(input_a[14] | input_a[3]);
  assign popcount35_g3qe_core_144 = ~(input_a[24] | input_a[21]);
  assign popcount35_g3qe_core_145 = input_a[26] & input_a[4];
  assign popcount35_g3qe_core_146 = ~input_a[30];
  assign popcount35_g3qe_core_149 = input_a[32] | input_a[9];
  assign popcount35_g3qe_core_151 = ~input_a[20];
  assign popcount35_g3qe_core_153 = input_a[1] ^ input_a[3];
  assign popcount35_g3qe_core_154 = input_a[15] ^ input_a[22];
  assign popcount35_g3qe_core_155 = input_a[3] ^ input_a[3];
  assign popcount35_g3qe_core_156 = ~input_a[28];
  assign popcount35_g3qe_core_157 = input_a[2] & input_a[10];
  assign popcount35_g3qe_core_158 = ~(input_a[1] | input_a[0]);
  assign popcount35_g3qe_core_162 = ~(input_a[18] | input_a[27]);
  assign popcount35_g3qe_core_164 = ~(input_a[11] | input_a[28]);
  assign popcount35_g3qe_core_170 = input_a[34] ^ input_a[3];
  assign popcount35_g3qe_core_174 = input_a[19] & input_a[34];
  assign popcount35_g3qe_core_177 = ~(input_a[6] | input_a[32]);
  assign popcount35_g3qe_core_178 = input_a[21] | input_a[32];
  assign popcount35_g3qe_core_180 = input_a[1] | input_a[1];
  assign popcount35_g3qe_core_185 = ~(input_a[8] | input_a[3]);
  assign popcount35_g3qe_core_187 = ~(input_a[17] ^ input_a[33]);
  assign popcount35_g3qe_core_188 = ~input_a[30];
  assign popcount35_g3qe_core_193 = ~(input_a[20] ^ input_a[28]);
  assign popcount35_g3qe_core_195 = input_a[17] | input_a[11];
  assign popcount35_g3qe_core_196 = input_a[0] ^ input_a[26];
  assign popcount35_g3qe_core_199 = input_a[23] | input_a[23];
  assign popcount35_g3qe_core_200 = input_a[30] | input_a[23];
  assign popcount35_g3qe_core_202 = ~(input_a[13] & input_a[12]);
  assign popcount35_g3qe_core_203 = input_a[9] ^ input_a[31];
  assign popcount35_g3qe_core_204 = input_a[15] & input_a[31];
  assign popcount35_g3qe_core_205 = popcount35_g3qe_core_180 & input_a[23];
  assign popcount35_g3qe_core_206 = ~input_a[16];
  assign popcount35_g3qe_core_207 = ~input_a[4];
  assign popcount35_g3qe_core_208 = popcount35_g3qe_core_205 | input_a[12];
  assign popcount35_g3qe_core_211 = input_a[0] ^ popcount35_g3qe_core_208;
  assign popcount35_g3qe_core_212 = input_a[0] & popcount35_g3qe_core_208;
  assign popcount35_g3qe_core_215 = ~(input_a[24] & input_a[7]);
  assign popcount35_g3qe_core_217 = ~(input_a[34] | input_a[3]);
  assign popcount35_g3qe_core_218 = ~(input_a[2] | input_a[16]);
  assign popcount35_g3qe_core_219 = ~(input_a[5] & input_a[21]);
  assign popcount35_g3qe_core_220 = ~(input_a[10] & input_a[5]);
  assign popcount35_g3qe_core_221 = ~(input_a[31] & input_a[17]);
  assign popcount35_g3qe_core_222 = ~(input_a[12] | input_a[1]);
  assign popcount35_g3qe_core_223 = popcount35_g3qe_core_135 ^ popcount35_g3qe_core_211;
  assign popcount35_g3qe_core_224 = popcount35_g3qe_core_135 & popcount35_g3qe_core_211;
  assign popcount35_g3qe_core_225 = popcount35_g3qe_core_223 ^ popcount35_g3qe_core_222;
  assign popcount35_g3qe_core_226 = popcount35_g3qe_core_223 & popcount35_g3qe_core_222;
  assign popcount35_g3qe_core_227 = popcount35_g3qe_core_224 | popcount35_g3qe_core_226;
  assign popcount35_g3qe_core_230 = popcount35_g3qe_core_212 ^ popcount35_g3qe_core_227;
  assign popcount35_g3qe_core_234 = input_a[13] & input_a[18];
  assign popcount35_g3qe_core_237 = input_a[29] & input_a[14];
  assign popcount35_g3qe_core_238 = ~popcount35_g3qe_core_113_not;
  assign popcount35_g3qe_core_239 = popcount35_g3qe_core_113_not & popcount35_g3qe_core_202;
  assign popcount35_g3qe_core_240 = popcount35_g3qe_core_117 ^ popcount35_g3qe_core_220;
  assign popcount35_g3qe_core_241 = popcount35_g3qe_core_117 & popcount35_g3qe_core_220;
  assign popcount35_g3qe_core_242 = popcount35_g3qe_core_240 ^ popcount35_g3qe_core_239;
  assign popcount35_g3qe_core_243 = popcount35_g3qe_core_240 & popcount35_g3qe_core_239;
  assign popcount35_g3qe_core_244 = popcount35_g3qe_core_241 | popcount35_g3qe_core_243;
  assign popcount35_g3qe_core_245 = popcount35_g3qe_core_120 ^ popcount35_g3qe_core_225;
  assign popcount35_g3qe_core_246 = popcount35_g3qe_core_120 & popcount35_g3qe_core_225;
  assign popcount35_g3qe_core_247 = popcount35_g3qe_core_245 ^ popcount35_g3qe_core_244;
  assign popcount35_g3qe_core_248 = popcount35_g3qe_core_245 & popcount35_g3qe_core_244;
  assign popcount35_g3qe_core_249 = popcount35_g3qe_core_246 | popcount35_g3qe_core_248;
  assign popcount35_g3qe_core_250 = popcount35_g3qe_core_127 ^ popcount35_g3qe_core_230;
  assign popcount35_g3qe_core_251 = popcount35_g3qe_core_127 & popcount35_g3qe_core_230;
  assign popcount35_g3qe_core_252 = popcount35_g3qe_core_250 ^ popcount35_g3qe_core_249;
  assign popcount35_g3qe_core_253 = popcount35_g3qe_core_250 & popcount35_g3qe_core_249;
  assign popcount35_g3qe_core_254 = popcount35_g3qe_core_251 | popcount35_g3qe_core_253;
  assign popcount35_g3qe_core_257 = popcount35_g3qe_core_129 ^ popcount35_g3qe_core_254;
  assign popcount35_g3qe_core_258 = popcount35_g3qe_core_129 & popcount35_g3qe_core_254;
  assign popcount35_g3qe_core_261 = ~(input_a[27] ^ input_a[29]);
  assign popcount35_g3qe_core_263 = input_a[14] | input_a[6];
  assign popcount35_g3qe_core_264 = input_a[15] & input_a[1];

  assign popcount35_g3qe_out[0] = popcount35_g3qe_core_238;
  assign popcount35_g3qe_out[1] = popcount35_g3qe_core_242;
  assign popcount35_g3qe_out[2] = popcount35_g3qe_core_247;
  assign popcount35_g3qe_out[3] = popcount35_g3qe_core_252;
  assign popcount35_g3qe_out[4] = popcount35_g3qe_core_257;
  assign popcount35_g3qe_out[5] = popcount35_g3qe_core_258;
endmodule