// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.47028
// WCE=53.0
// EP=0.908513%
// Printed PDK parameters:
//  Area=49365095.0
//  Delay=69493248.0
//  Power=1874200.0

module popcount35_hxy9(input [34:0] input_a, output [5:0] popcount35_hxy9_out);
  wire popcount35_hxy9_core_037;
  wire popcount35_hxy9_core_038;
  wire popcount35_hxy9_core_040;
  wire popcount35_hxy9_core_041;
  wire popcount35_hxy9_core_042;
  wire popcount35_hxy9_core_043;
  wire popcount35_hxy9_core_044;
  wire popcount35_hxy9_core_046;
  wire popcount35_hxy9_core_047;
  wire popcount35_hxy9_core_048;
  wire popcount35_hxy9_core_049;
  wire popcount35_hxy9_core_053;
  wire popcount35_hxy9_core_060;
  wire popcount35_hxy9_core_068;
  wire popcount35_hxy9_core_069;
  wire popcount35_hxy9_core_071;
  wire popcount35_hxy9_core_073;
  wire popcount35_hxy9_core_075;
  wire popcount35_hxy9_core_079_not;
  wire popcount35_hxy9_core_082;
  wire popcount35_hxy9_core_084;
  wire popcount35_hxy9_core_085;
  wire popcount35_hxy9_core_086;
  wire popcount35_hxy9_core_087;
  wire popcount35_hxy9_core_088;
  wire popcount35_hxy9_core_089;
  wire popcount35_hxy9_core_090;
  wire popcount35_hxy9_core_091;
  wire popcount35_hxy9_core_092;
  wire popcount35_hxy9_core_094;
  wire popcount35_hxy9_core_095;
  wire popcount35_hxy9_core_097;
  wire popcount35_hxy9_core_098;
  wire popcount35_hxy9_core_099;
  wire popcount35_hxy9_core_101;
  wire popcount35_hxy9_core_102;
  wire popcount35_hxy9_core_103;
  wire popcount35_hxy9_core_104;
  wire popcount35_hxy9_core_105;
  wire popcount35_hxy9_core_108;
  wire popcount35_hxy9_core_109;
  wire popcount35_hxy9_core_111;
  wire popcount35_hxy9_core_112;
  wire popcount35_hxy9_core_115;
  wire popcount35_hxy9_core_120;
  wire popcount35_hxy9_core_121;
  wire popcount35_hxy9_core_125;
  wire popcount35_hxy9_core_126;
  wire popcount35_hxy9_core_127;
  wire popcount35_hxy9_core_128;
  wire popcount35_hxy9_core_129;
  wire popcount35_hxy9_core_133;
  wire popcount35_hxy9_core_135;
  wire popcount35_hxy9_core_136;
  wire popcount35_hxy9_core_138;
  wire popcount35_hxy9_core_139;
  wire popcount35_hxy9_core_140;
  wire popcount35_hxy9_core_141_not;
  wire popcount35_hxy9_core_142;
  wire popcount35_hxy9_core_146;
  wire popcount35_hxy9_core_148;
  wire popcount35_hxy9_core_149;
  wire popcount35_hxy9_core_150;
  wire popcount35_hxy9_core_153;
  wire popcount35_hxy9_core_155;
  wire popcount35_hxy9_core_157;
  wire popcount35_hxy9_core_158;
  wire popcount35_hxy9_core_160;
  wire popcount35_hxy9_core_162;
  wire popcount35_hxy9_core_163;
  wire popcount35_hxy9_core_164;
  wire popcount35_hxy9_core_167;
  wire popcount35_hxy9_core_169;
  wire popcount35_hxy9_core_170;
  wire popcount35_hxy9_core_174;
  wire popcount35_hxy9_core_177;
  wire popcount35_hxy9_core_182;
  wire popcount35_hxy9_core_183;
  wire popcount35_hxy9_core_185;
  wire popcount35_hxy9_core_186;
  wire popcount35_hxy9_core_187;
  wire popcount35_hxy9_core_188;
  wire popcount35_hxy9_core_189;
  wire popcount35_hxy9_core_190;
  wire popcount35_hxy9_core_191;
  wire popcount35_hxy9_core_192;
  wire popcount35_hxy9_core_193;
  wire popcount35_hxy9_core_194;
  wire popcount35_hxy9_core_195;
  wire popcount35_hxy9_core_196;
  wire popcount35_hxy9_core_197;
  wire popcount35_hxy9_core_198;
  wire popcount35_hxy9_core_199;
  wire popcount35_hxy9_core_200;
  wire popcount35_hxy9_core_201;
  wire popcount35_hxy9_core_202;
  wire popcount35_hxy9_core_203;
  wire popcount35_hxy9_core_204;
  wire popcount35_hxy9_core_205;
  wire popcount35_hxy9_core_206;
  wire popcount35_hxy9_core_207_not;
  wire popcount35_hxy9_core_208;
  wire popcount35_hxy9_core_209;
  wire popcount35_hxy9_core_210;
  wire popcount35_hxy9_core_211;
  wire popcount35_hxy9_core_212;
  wire popcount35_hxy9_core_213;
  wire popcount35_hxy9_core_214;
  wire popcount35_hxy9_core_215;
  wire popcount35_hxy9_core_216;
  wire popcount35_hxy9_core_217;
  wire popcount35_hxy9_core_219;
  wire popcount35_hxy9_core_220_not;
  wire popcount35_hxy9_core_222;
  wire popcount35_hxy9_core_223;
  wire popcount35_hxy9_core_225;
  wire popcount35_hxy9_core_226;
  wire popcount35_hxy9_core_230;
  wire popcount35_hxy9_core_231;
  wire popcount35_hxy9_core_234;
  wire popcount35_hxy9_core_238;
  wire popcount35_hxy9_core_239;
  wire popcount35_hxy9_core_240;
  wire popcount35_hxy9_core_241;
  wire popcount35_hxy9_core_243;
  wire popcount35_hxy9_core_245;
  wire popcount35_hxy9_core_246;
  wire popcount35_hxy9_core_247_not;
  wire popcount35_hxy9_core_249;
  wire popcount35_hxy9_core_250;
  wire popcount35_hxy9_core_251;
  wire popcount35_hxy9_core_252;
  wire popcount35_hxy9_core_253;
  wire popcount35_hxy9_core_254;
  wire popcount35_hxy9_core_255;
  wire popcount35_hxy9_core_257;
  wire popcount35_hxy9_core_258;
  wire popcount35_hxy9_core_259;
  wire popcount35_hxy9_core_260;
  wire popcount35_hxy9_core_262;
  wire popcount35_hxy9_core_263;
  wire popcount35_hxy9_core_264;

  assign popcount35_hxy9_core_037 = input_a[0] | input_a[21];
  assign popcount35_hxy9_core_038 = input_a[0] & input_a[17];
  assign popcount35_hxy9_core_040 = input_a[2] & input_a[27];
  assign popcount35_hxy9_core_041 = ~(input_a[10] & input_a[10]);
  assign popcount35_hxy9_core_042 = popcount35_hxy9_core_037 & input_a[2];
  assign popcount35_hxy9_core_043 = popcount35_hxy9_core_038 ^ popcount35_hxy9_core_040;
  assign popcount35_hxy9_core_044 = popcount35_hxy9_core_038 & input_a[33];
  assign popcount35_hxy9_core_046 = input_a[31] & popcount35_hxy9_core_042;
  assign popcount35_hxy9_core_047 = popcount35_hxy9_core_044 | popcount35_hxy9_core_046;
  assign popcount35_hxy9_core_048 = ~input_a[4];
  assign popcount35_hxy9_core_049 = input_a[4] & input_a[6];
  assign popcount35_hxy9_core_053 = popcount35_hxy9_core_048 & input_a[24];
  assign popcount35_hxy9_core_060 = input_a[24] & input_a[29];
  assign popcount35_hxy9_core_068 = popcount35_hxy9_core_047 ^ popcount35_hxy9_core_043;
  assign popcount35_hxy9_core_069 = popcount35_hxy9_core_047 & popcount35_hxy9_core_043;
  assign popcount35_hxy9_core_071 = input_a[23] ^ input_a[7];
  assign popcount35_hxy9_core_073 = input_a[10] ^ input_a[13];
  assign popcount35_hxy9_core_075 = popcount35_hxy9_core_071 ^ input_a[3];
  assign popcount35_hxy9_core_079_not = ~popcount35_hxy9_core_071;
  assign popcount35_hxy9_core_082 = input_a[12] & input_a[13];
  assign popcount35_hxy9_core_084 = ~(input_a[3] | input_a[19]);
  assign popcount35_hxy9_core_085 = input_a[23] & input_a[16];
  assign popcount35_hxy9_core_086 = input_a[33] ^ input_a[11];
  assign popcount35_hxy9_core_087 = input_a[14] & popcount35_hxy9_core_084;
  assign popcount35_hxy9_core_088 = popcount35_hxy9_core_085 ^ popcount35_hxy9_core_087;
  assign popcount35_hxy9_core_089 = popcount35_hxy9_core_085 & popcount35_hxy9_core_087;
  assign popcount35_hxy9_core_090 = input_a[5] ^ popcount35_hxy9_core_086;
  assign popcount35_hxy9_core_091 = popcount35_hxy9_core_082 & popcount35_hxy9_core_086;
  assign popcount35_hxy9_core_092 = input_a[22] | popcount35_hxy9_core_088;
  assign popcount35_hxy9_core_094 = popcount35_hxy9_core_092 ^ popcount35_hxy9_core_091;
  assign popcount35_hxy9_core_095 = popcount35_hxy9_core_092 & popcount35_hxy9_core_091;
  assign popcount35_hxy9_core_097 = popcount35_hxy9_core_089 ^ popcount35_hxy9_core_095;
  assign popcount35_hxy9_core_098 = popcount35_hxy9_core_089 & popcount35_hxy9_core_095;
  assign popcount35_hxy9_core_099 = popcount35_hxy9_core_075 ^ popcount35_hxy9_core_090;
  assign popcount35_hxy9_core_101 = popcount35_hxy9_core_079_not ^ popcount35_hxy9_core_094;
  assign popcount35_hxy9_core_102 = popcount35_hxy9_core_079_not & popcount35_hxy9_core_094;
  assign popcount35_hxy9_core_103 = popcount35_hxy9_core_101 | input_a[22];
  assign popcount35_hxy9_core_104 = popcount35_hxy9_core_101 & input_a[22];
  assign popcount35_hxy9_core_105 = popcount35_hxy9_core_102 | popcount35_hxy9_core_104;
  assign popcount35_hxy9_core_108 = popcount35_hxy9_core_097 ^ popcount35_hxy9_core_105;
  assign popcount35_hxy9_core_109 = popcount35_hxy9_core_097 & popcount35_hxy9_core_105;
  assign popcount35_hxy9_core_111 = popcount35_hxy9_core_098 ^ popcount35_hxy9_core_109;
  assign popcount35_hxy9_core_112 = popcount35_hxy9_core_098 & input_a[29];
  assign popcount35_hxy9_core_115 = input_a[8] | input_a[29];
  assign popcount35_hxy9_core_120 = popcount35_hxy9_core_068 ^ popcount35_hxy9_core_108;
  assign popcount35_hxy9_core_121 = popcount35_hxy9_core_068 & popcount35_hxy9_core_108;
  assign popcount35_hxy9_core_125 = popcount35_hxy9_core_069 & popcount35_hxy9_core_111;
  assign popcount35_hxy9_core_126 = input_a[5] & input_a[1];
  assign popcount35_hxy9_core_127 = popcount35_hxy9_core_125 ^ popcount35_hxy9_core_121;
  assign popcount35_hxy9_core_128 = input_a[20] & input_a[11];
  assign popcount35_hxy9_core_129 = ~popcount35_hxy9_core_126;
  assign popcount35_hxy9_core_133 = ~(input_a[17] & input_a[18]);
  assign popcount35_hxy9_core_135 = ~(input_a[34] | input_a[9]);
  assign popcount35_hxy9_core_136 = ~(input_a[9] & input_a[19]);
  assign popcount35_hxy9_core_138 = ~popcount35_hxy9_core_133;
  assign popcount35_hxy9_core_139 = ~input_a[28];
  assign popcount35_hxy9_core_140 = popcount35_hxy9_core_138 & input_a[28];
  assign popcount35_hxy9_core_141_not = ~popcount35_hxy9_core_138;
  assign popcount35_hxy9_core_142 = input_a[5] | input_a[28];
  assign popcount35_hxy9_core_146 = ~(input_a[15] ^ input_a[12]);
  assign popcount35_hxy9_core_148 = input_a[21] & input_a[24];
  assign popcount35_hxy9_core_149 = ~(input_a[27] | input_a[5]);
  assign popcount35_hxy9_core_150 = popcount35_hxy9_core_146 & input_a[21];
  assign popcount35_hxy9_core_153 = ~(input_a[16] ^ input_a[32]);
  assign popcount35_hxy9_core_155 = input_a[21] | input_a[20];
  assign popcount35_hxy9_core_157 = input_a[0] | input_a[30];
  assign popcount35_hxy9_core_158 = input_a[32] ^ input_a[21];
  assign popcount35_hxy9_core_160 = ~(popcount35_hxy9_core_136 | input_a[31]);
  assign popcount35_hxy9_core_162 = ~popcount35_hxy9_core_140;
  assign popcount35_hxy9_core_163 = input_a[18] & popcount35_hxy9_core_155;
  assign popcount35_hxy9_core_164 = input_a[29] ^ input_a[5];
  assign popcount35_hxy9_core_167 = input_a[24] | popcount35_hxy9_core_158;
  assign popcount35_hxy9_core_169 = input_a[18] ^ popcount35_hxy9_core_163;
  assign popcount35_hxy9_core_170 = ~(popcount35_hxy9_core_167 | input_a[14]);
  assign popcount35_hxy9_core_174 = ~(input_a[26] & input_a[27]);
  assign popcount35_hxy9_core_177 = input_a[28] & input_a[25];
  assign popcount35_hxy9_core_182 = ~(popcount35_hxy9_core_177 & input_a[29]);
  assign popcount35_hxy9_core_183 = popcount35_hxy9_core_177 & input_a[14];
  assign popcount35_hxy9_core_185 = input_a[1] | input_a[15];
  assign popcount35_hxy9_core_186 = input_a[30] & input_a[19];
  assign popcount35_hxy9_core_187 = input_a[33] ^ input_a[34];
  assign popcount35_hxy9_core_188 = input_a[33] & input_a[34];
  assign popcount35_hxy9_core_189 = ~input_a[9];
  assign popcount35_hxy9_core_190 = input_a[21] & popcount35_hxy9_core_187;
  assign popcount35_hxy9_core_191 = popcount35_hxy9_core_188 | popcount35_hxy9_core_190;
  assign popcount35_hxy9_core_192 = popcount35_hxy9_core_188 & popcount35_hxy9_core_190;
  assign popcount35_hxy9_core_193 = input_a[13] ^ input_a[28];
  assign popcount35_hxy9_core_194 = popcount35_hxy9_core_185 & input_a[23];
  assign popcount35_hxy9_core_195 = popcount35_hxy9_core_186 ^ popcount35_hxy9_core_191;
  assign popcount35_hxy9_core_196 = popcount35_hxy9_core_186 & popcount35_hxy9_core_191;
  assign popcount35_hxy9_core_197 = popcount35_hxy9_core_195 ^ popcount35_hxy9_core_194;
  assign popcount35_hxy9_core_198 = popcount35_hxy9_core_195 & popcount35_hxy9_core_194;
  assign popcount35_hxy9_core_199 = popcount35_hxy9_core_196 | popcount35_hxy9_core_198;
  assign popcount35_hxy9_core_200 = popcount35_hxy9_core_192 ^ popcount35_hxy9_core_199;
  assign popcount35_hxy9_core_201 = popcount35_hxy9_core_192 & input_a[8];
  assign popcount35_hxy9_core_202 = input_a[12] ^ input_a[13];
  assign popcount35_hxy9_core_203 = input_a[2] ^ input_a[18];
  assign popcount35_hxy9_core_204 = ~popcount35_hxy9_core_182;
  assign popcount35_hxy9_core_205 = popcount35_hxy9_core_182 & popcount35_hxy9_core_197;
  assign popcount35_hxy9_core_206 = input_a[1] ^ input_a[19];
  assign popcount35_hxy9_core_207_not = ~popcount35_hxy9_core_203;
  assign popcount35_hxy9_core_208 = popcount35_hxy9_core_205 | input_a[11];
  assign popcount35_hxy9_core_209 = popcount35_hxy9_core_183 ^ popcount35_hxy9_core_200;
  assign popcount35_hxy9_core_210 = popcount35_hxy9_core_183 & popcount35_hxy9_core_200;
  assign popcount35_hxy9_core_211 = popcount35_hxy9_core_209 ^ popcount35_hxy9_core_208;
  assign popcount35_hxy9_core_212 = popcount35_hxy9_core_209 & popcount35_hxy9_core_208;
  assign popcount35_hxy9_core_213 = popcount35_hxy9_core_210 | popcount35_hxy9_core_212;
  assign popcount35_hxy9_core_214 = popcount35_hxy9_core_201 ^ popcount35_hxy9_core_213;
  assign popcount35_hxy9_core_215 = popcount35_hxy9_core_201 & input_a[24];
  assign popcount35_hxy9_core_216 = input_a[23] & popcount35_hxy9_core_202;
  assign popcount35_hxy9_core_217 = input_a[20] & input_a[2];
  assign popcount35_hxy9_core_219 = input_a[5] & popcount35_hxy9_core_206;
  assign popcount35_hxy9_core_220_not = ~popcount35_hxy9_core_217;
  assign popcount35_hxy9_core_222 = input_a[3] | input_a[24];
  assign popcount35_hxy9_core_223 = popcount35_hxy9_core_169 ^ popcount35_hxy9_core_211;
  assign popcount35_hxy9_core_225 = popcount35_hxy9_core_223 ^ popcount35_hxy9_core_222;
  assign popcount35_hxy9_core_226 = popcount35_hxy9_core_223 & popcount35_hxy9_core_222;
  assign popcount35_hxy9_core_230 = popcount35_hxy9_core_214 ^ popcount35_hxy9_core_226;
  assign popcount35_hxy9_core_231 = popcount35_hxy9_core_214 & popcount35_hxy9_core_226;
  assign popcount35_hxy9_core_234 = input_a[31] & popcount35_hxy9_core_215;
  assign popcount35_hxy9_core_238 = input_a[7] ^ input_a[4];
  assign popcount35_hxy9_core_239 = input_a[26] & popcount35_hxy9_core_216;
  assign popcount35_hxy9_core_240 = input_a[6] ^ input_a[34];
  assign popcount35_hxy9_core_241 = input_a[6] & popcount35_hxy9_core_220_not;
  assign popcount35_hxy9_core_243 = ~input_a[22];
  assign popcount35_hxy9_core_245 = popcount35_hxy9_core_120 ^ popcount35_hxy9_core_225;
  assign popcount35_hxy9_core_246 = popcount35_hxy9_core_120 & popcount35_hxy9_core_225;
  assign popcount35_hxy9_core_247_not = ~popcount35_hxy9_core_245;
  assign popcount35_hxy9_core_249 = popcount35_hxy9_core_246 | popcount35_hxy9_core_245;
  assign popcount35_hxy9_core_250 = popcount35_hxy9_core_127 ^ popcount35_hxy9_core_230;
  assign popcount35_hxy9_core_251 = popcount35_hxy9_core_127 & popcount35_hxy9_core_230;
  assign popcount35_hxy9_core_252 = popcount35_hxy9_core_250 ^ popcount35_hxy9_core_249;
  assign popcount35_hxy9_core_253 = popcount35_hxy9_core_250 & popcount35_hxy9_core_249;
  assign popcount35_hxy9_core_254 = popcount35_hxy9_core_251 | popcount35_hxy9_core_253;
  assign popcount35_hxy9_core_255 = popcount35_hxy9_core_112 ^ popcount35_hxy9_core_231;
  assign popcount35_hxy9_core_257 = popcount35_hxy9_core_255 ^ popcount35_hxy9_core_254;
  assign popcount35_hxy9_core_258 = popcount35_hxy9_core_255 & popcount35_hxy9_core_254;
  assign popcount35_hxy9_core_259 = popcount35_hxy9_core_112 | popcount35_hxy9_core_258;
  assign popcount35_hxy9_core_260 = popcount35_hxy9_core_112 ^ popcount35_hxy9_core_234;
  assign popcount35_hxy9_core_262 = popcount35_hxy9_core_260 | popcount35_hxy9_core_259;
  assign popcount35_hxy9_core_263 = ~(popcount35_hxy9_core_260 | popcount35_hxy9_core_259);
  assign popcount35_hxy9_core_264 = input_a[27] | input_a[13];

  assign popcount35_hxy9_out[0] = popcount35_hxy9_core_044;
  assign popcount35_hxy9_out[1] = popcount35_hxy9_core_103;
  assign popcount35_hxy9_out[2] = popcount35_hxy9_core_247_not;
  assign popcount35_hxy9_out[3] = popcount35_hxy9_core_252;
  assign popcount35_hxy9_out[4] = popcount35_hxy9_core_257;
  assign popcount35_hxy9_out[5] = popcount35_hxy9_core_262;
endmodule