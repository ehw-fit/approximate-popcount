// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.74882
// WCE=27.0
// EP=0.951668%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_4bty(input [28:0] input_a, output [4:0] popcount29_4bty_out);
  wire popcount29_4bty_core_031;
  wire popcount29_4bty_core_032;
  wire popcount29_4bty_core_033;
  wire popcount29_4bty_core_034;
  wire popcount29_4bty_core_035;
  wire popcount29_4bty_core_036;
  wire popcount29_4bty_core_039;
  wire popcount29_4bty_core_040;
  wire popcount29_4bty_core_041;
  wire popcount29_4bty_core_043;
  wire popcount29_4bty_core_046;
  wire popcount29_4bty_core_050;
  wire popcount29_4bty_core_052;
  wire popcount29_4bty_core_053;
  wire popcount29_4bty_core_054;
  wire popcount29_4bty_core_056;
  wire popcount29_4bty_core_057;
  wire popcount29_4bty_core_059;
  wire popcount29_4bty_core_060;
  wire popcount29_4bty_core_061;
  wire popcount29_4bty_core_062;
  wire popcount29_4bty_core_064;
  wire popcount29_4bty_core_068;
  wire popcount29_4bty_core_070;
  wire popcount29_4bty_core_071;
  wire popcount29_4bty_core_073;
  wire popcount29_4bty_core_074;
  wire popcount29_4bty_core_075;
  wire popcount29_4bty_core_077;
  wire popcount29_4bty_core_078;
  wire popcount29_4bty_core_079;
  wire popcount29_4bty_core_080;
  wire popcount29_4bty_core_081;
  wire popcount29_4bty_core_082;
  wire popcount29_4bty_core_083;
  wire popcount29_4bty_core_085;
  wire popcount29_4bty_core_086;
  wire popcount29_4bty_core_087;
  wire popcount29_4bty_core_088;
  wire popcount29_4bty_core_090;
  wire popcount29_4bty_core_092;
  wire popcount29_4bty_core_093;
  wire popcount29_4bty_core_094;
  wire popcount29_4bty_core_095;
  wire popcount29_4bty_core_096;
  wire popcount29_4bty_core_097;
  wire popcount29_4bty_core_099;
  wire popcount29_4bty_core_101;
  wire popcount29_4bty_core_102;
  wire popcount29_4bty_core_105;
  wire popcount29_4bty_core_106;
  wire popcount29_4bty_core_107;
  wire popcount29_4bty_core_109;
  wire popcount29_4bty_core_110;
  wire popcount29_4bty_core_111;
  wire popcount29_4bty_core_115;
  wire popcount29_4bty_core_117;
  wire popcount29_4bty_core_118;
  wire popcount29_4bty_core_119;
  wire popcount29_4bty_core_123;
  wire popcount29_4bty_core_126;
  wire popcount29_4bty_core_128;
  wire popcount29_4bty_core_131_not;
  wire popcount29_4bty_core_133;
  wire popcount29_4bty_core_134;
  wire popcount29_4bty_core_136;
  wire popcount29_4bty_core_138;
  wire popcount29_4bty_core_140;
  wire popcount29_4bty_core_142;
  wire popcount29_4bty_core_143;
  wire popcount29_4bty_core_145;
  wire popcount29_4bty_core_146;
  wire popcount29_4bty_core_147;
  wire popcount29_4bty_core_148;
  wire popcount29_4bty_core_149;
  wire popcount29_4bty_core_152;
  wire popcount29_4bty_core_153;
  wire popcount29_4bty_core_154;
  wire popcount29_4bty_core_155;
  wire popcount29_4bty_core_156;
  wire popcount29_4bty_core_160;
  wire popcount29_4bty_core_161;
  wire popcount29_4bty_core_162;
  wire popcount29_4bty_core_163;
  wire popcount29_4bty_core_164;
  wire popcount29_4bty_core_165;
  wire popcount29_4bty_core_166;
  wire popcount29_4bty_core_168;
  wire popcount29_4bty_core_170;
  wire popcount29_4bty_core_171;
  wire popcount29_4bty_core_172_not;
  wire popcount29_4bty_core_173;
  wire popcount29_4bty_core_174;
  wire popcount29_4bty_core_176;
  wire popcount29_4bty_core_178;
  wire popcount29_4bty_core_182;
  wire popcount29_4bty_core_184;
  wire popcount29_4bty_core_185;
  wire popcount29_4bty_core_187;
  wire popcount29_4bty_core_190;
  wire popcount29_4bty_core_191_not;
  wire popcount29_4bty_core_192;
  wire popcount29_4bty_core_194;
  wire popcount29_4bty_core_195;
  wire popcount29_4bty_core_196;
  wire popcount29_4bty_core_203;
  wire popcount29_4bty_core_204;
  wire popcount29_4bty_core_205;
  wire popcount29_4bty_core_206;
  wire popcount29_4bty_core_207;

  assign popcount29_4bty_core_031 = ~input_a[0];
  assign popcount29_4bty_core_032 = input_a[9] & input_a[18];
  assign popcount29_4bty_core_033 = ~(input_a[4] ^ input_a[17]);
  assign popcount29_4bty_core_034 = input_a[3] ^ input_a[5];
  assign popcount29_4bty_core_035 = input_a[2] & input_a[6];
  assign popcount29_4bty_core_036 = input_a[24] ^ input_a[0];
  assign popcount29_4bty_core_039 = ~input_a[15];
  assign popcount29_4bty_core_040 = input_a[6] ^ input_a[19];
  assign popcount29_4bty_core_041 = input_a[26] | input_a[26];
  assign popcount29_4bty_core_043 = ~(input_a[0] & input_a[15]);
  assign popcount29_4bty_core_046 = ~(input_a[9] | input_a[12]);
  assign popcount29_4bty_core_050 = ~(input_a[22] ^ input_a[27]);
  assign popcount29_4bty_core_052 = ~(input_a[21] & input_a[28]);
  assign popcount29_4bty_core_053 = ~(input_a[27] | input_a[24]);
  assign popcount29_4bty_core_054 = ~(input_a[13] | input_a[10]);
  assign popcount29_4bty_core_056 = input_a[12] | input_a[9];
  assign popcount29_4bty_core_057 = ~(input_a[23] ^ input_a[11]);
  assign popcount29_4bty_core_059 = input_a[13] & input_a[11];
  assign popcount29_4bty_core_060 = ~input_a[2];
  assign popcount29_4bty_core_061 = input_a[23] & input_a[27];
  assign popcount29_4bty_core_062 = ~(input_a[23] ^ input_a[11]);
  assign popcount29_4bty_core_064 = ~(input_a[14] & input_a[18]);
  assign popcount29_4bty_core_068 = input_a[28] | input_a[21];
  assign popcount29_4bty_core_070 = input_a[6] ^ input_a[26];
  assign popcount29_4bty_core_071 = ~(input_a[11] ^ input_a[15]);
  assign popcount29_4bty_core_073 = input_a[9] | input_a[9];
  assign popcount29_4bty_core_074 = input_a[3] | input_a[10];
  assign popcount29_4bty_core_075 = ~input_a[6];
  assign popcount29_4bty_core_077 = ~(input_a[28] | input_a[11]);
  assign popcount29_4bty_core_078 = input_a[15] | input_a[4];
  assign popcount29_4bty_core_079 = input_a[6] ^ input_a[15];
  assign popcount29_4bty_core_080 = ~input_a[23];
  assign popcount29_4bty_core_081 = ~(input_a[17] ^ input_a[4]);
  assign popcount29_4bty_core_082 = ~(input_a[1] | input_a[21]);
  assign popcount29_4bty_core_083 = input_a[0] | input_a[8];
  assign popcount29_4bty_core_085 = input_a[3] ^ input_a[6];
  assign popcount29_4bty_core_086 = ~(input_a[6] & input_a[14]);
  assign popcount29_4bty_core_087 = input_a[3] ^ input_a[2];
  assign popcount29_4bty_core_088 = input_a[21] & input_a[15];
  assign popcount29_4bty_core_090 = input_a[6] | input_a[1];
  assign popcount29_4bty_core_092 = ~input_a[17];
  assign popcount29_4bty_core_093 = ~(input_a[11] | input_a[9]);
  assign popcount29_4bty_core_094 = ~(input_a[13] ^ input_a[20]);
  assign popcount29_4bty_core_095 = ~(input_a[8] | input_a[10]);
  assign popcount29_4bty_core_096 = ~(input_a[26] ^ input_a[22]);
  assign popcount29_4bty_core_097 = ~(input_a[6] ^ input_a[3]);
  assign popcount29_4bty_core_099 = input_a[14] | input_a[16];
  assign popcount29_4bty_core_101 = input_a[15] ^ input_a[9];
  assign popcount29_4bty_core_102 = input_a[5] | input_a[2];
  assign popcount29_4bty_core_105 = input_a[27] & input_a[5];
  assign popcount29_4bty_core_106 = ~(input_a[9] ^ input_a[8]);
  assign popcount29_4bty_core_107 = ~input_a[8];
  assign popcount29_4bty_core_109 = ~(input_a[19] ^ input_a[15]);
  assign popcount29_4bty_core_110 = ~(input_a[14] | input_a[7]);
  assign popcount29_4bty_core_111 = input_a[25] | input_a[27];
  assign popcount29_4bty_core_115 = ~(input_a[5] | input_a[23]);
  assign popcount29_4bty_core_117 = input_a[9] ^ input_a[28];
  assign popcount29_4bty_core_118 = ~(input_a[22] & input_a[23]);
  assign popcount29_4bty_core_119 = ~(input_a[21] ^ input_a[22]);
  assign popcount29_4bty_core_123 = input_a[18] & input_a[28];
  assign popcount29_4bty_core_126 = ~input_a[23];
  assign popcount29_4bty_core_128 = ~(input_a[8] | input_a[6]);
  assign popcount29_4bty_core_131_not = ~input_a[8];
  assign popcount29_4bty_core_133 = ~(input_a[16] ^ input_a[18]);
  assign popcount29_4bty_core_134 = input_a[9] | input_a[17];
  assign popcount29_4bty_core_136 = ~input_a[2];
  assign popcount29_4bty_core_138 = input_a[9] ^ input_a[0];
  assign popcount29_4bty_core_140 = ~(input_a[7] ^ input_a[2]);
  assign popcount29_4bty_core_142 = input_a[2] | input_a[11];
  assign popcount29_4bty_core_143 = input_a[22] & input_a[18];
  assign popcount29_4bty_core_145 = ~input_a[22];
  assign popcount29_4bty_core_146 = ~input_a[2];
  assign popcount29_4bty_core_147 = input_a[17] & input_a[21];
  assign popcount29_4bty_core_148 = ~(input_a[21] ^ input_a[18]);
  assign popcount29_4bty_core_149 = ~(input_a[3] ^ input_a[12]);
  assign popcount29_4bty_core_152 = ~(input_a[1] & input_a[19]);
  assign popcount29_4bty_core_153 = ~(input_a[23] | input_a[3]);
  assign popcount29_4bty_core_154 = ~(input_a[4] & input_a[12]);
  assign popcount29_4bty_core_155 = input_a[16] | input_a[24];
  assign popcount29_4bty_core_156 = ~(input_a[13] & input_a[11]);
  assign popcount29_4bty_core_160 = ~(input_a[14] & input_a[14]);
  assign popcount29_4bty_core_161 = ~(input_a[12] | input_a[7]);
  assign popcount29_4bty_core_162 = input_a[18] | input_a[24];
  assign popcount29_4bty_core_163 = ~(input_a[22] | input_a[1]);
  assign popcount29_4bty_core_164 = ~(input_a[1] ^ input_a[14]);
  assign popcount29_4bty_core_165 = input_a[27] ^ input_a[13];
  assign popcount29_4bty_core_166 = ~(input_a[13] | input_a[6]);
  assign popcount29_4bty_core_168 = ~(input_a[6] ^ input_a[24]);
  assign popcount29_4bty_core_170 = input_a[27] & input_a[0];
  assign popcount29_4bty_core_171 = input_a[17] ^ input_a[20];
  assign popcount29_4bty_core_172_not = ~input_a[0];
  assign popcount29_4bty_core_173 = ~(input_a[5] | input_a[6]);
  assign popcount29_4bty_core_174 = ~(input_a[15] | input_a[10]);
  assign popcount29_4bty_core_176 = ~(input_a[25] & input_a[27]);
  assign popcount29_4bty_core_178 = input_a[0] | input_a[5];
  assign popcount29_4bty_core_182 = ~input_a[23];
  assign popcount29_4bty_core_184 = ~(input_a[15] | input_a[4]);
  assign popcount29_4bty_core_185 = ~(input_a[10] & input_a[12]);
  assign popcount29_4bty_core_187 = ~(input_a[16] ^ input_a[21]);
  assign popcount29_4bty_core_190 = ~input_a[21];
  assign popcount29_4bty_core_191_not = ~input_a[14];
  assign popcount29_4bty_core_192 = ~(input_a[22] & input_a[2]);
  assign popcount29_4bty_core_194 = ~(input_a[1] & input_a[28]);
  assign popcount29_4bty_core_195 = input_a[25] | input_a[8];
  assign popcount29_4bty_core_196 = ~(input_a[27] | input_a[16]);
  assign popcount29_4bty_core_203 = ~(input_a[22] ^ input_a[27]);
  assign popcount29_4bty_core_204 = ~(input_a[13] ^ input_a[8]);
  assign popcount29_4bty_core_205 = ~input_a[12];
  assign popcount29_4bty_core_206 = ~(input_a[6] & input_a[26]);
  assign popcount29_4bty_core_207 = input_a[6] ^ input_a[18];

  assign popcount29_4bty_out[0] = 1'b1;
  assign popcount29_4bty_out[1] = input_a[3];
  assign popcount29_4bty_out[2] = 1'b0;
  assign popcount29_4bty_out[3] = 1'b0;
  assign popcount29_4bty_out[4] = input_a[2];
endmodule