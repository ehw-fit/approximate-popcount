// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.58726
// WCE=11.0
// EP=0.80441%
// Printed PDK parameters:
//  Area=31367463.0
//  Delay=64410472.0
//  Power=1299200.0

module popcount32_0itb(input [31:0] input_a, output [5:0] popcount32_0itb_out);
  wire popcount32_0itb_core_034;
  wire popcount32_0itb_core_036;
  wire popcount32_0itb_core_037;
  wire popcount32_0itb_core_038;
  wire popcount32_0itb_core_041;
  wire popcount32_0itb_core_044_not;
  wire popcount32_0itb_core_045;
  wire popcount32_0itb_core_046;
  wire popcount32_0itb_core_048;
  wire popcount32_0itb_core_049;
  wire popcount32_0itb_core_050;
  wire popcount32_0itb_core_051;
  wire popcount32_0itb_core_053;
  wire popcount32_0itb_core_055;
  wire popcount32_0itb_core_056;
  wire popcount32_0itb_core_058;
  wire popcount32_0itb_core_059;
  wire popcount32_0itb_core_060;
  wire popcount32_0itb_core_061;
  wire popcount32_0itb_core_062;
  wire popcount32_0itb_core_064;
  wire popcount32_0itb_core_067;
  wire popcount32_0itb_core_068;
  wire popcount32_0itb_core_069;
  wire popcount32_0itb_core_070;
  wire popcount32_0itb_core_071;
  wire popcount32_0itb_core_072;
  wire popcount32_0itb_core_073;
  wire popcount32_0itb_core_074;
  wire popcount32_0itb_core_075;
  wire popcount32_0itb_core_076;
  wire popcount32_0itb_core_080;
  wire popcount32_0itb_core_081;
  wire popcount32_0itb_core_082;
  wire popcount32_0itb_core_083;
  wire popcount32_0itb_core_086;
  wire popcount32_0itb_core_087;
  wire popcount32_0itb_core_088;
  wire popcount32_0itb_core_089_not;
  wire popcount32_0itb_core_091;
  wire popcount32_0itb_core_092;
  wire popcount32_0itb_core_093;
  wire popcount32_0itb_core_095;
  wire popcount32_0itb_core_099;
  wire popcount32_0itb_core_100;
  wire popcount32_0itb_core_101;
  wire popcount32_0itb_core_103;
  wire popcount32_0itb_core_104;
  wire popcount32_0itb_core_105;
  wire popcount32_0itb_core_106;
  wire popcount32_0itb_core_107;
  wire popcount32_0itb_core_108;
  wire popcount32_0itb_core_109;
  wire popcount32_0itb_core_110;
  wire popcount32_0itb_core_111;
  wire popcount32_0itb_core_112;
  wire popcount32_0itb_core_113;
  wire popcount32_0itb_core_115;
  wire popcount32_0itb_core_117;
  wire popcount32_0itb_core_118_not;
  wire popcount32_0itb_core_119;
  wire popcount32_0itb_core_120;
  wire popcount32_0itb_core_121;
  wire popcount32_0itb_core_123;
  wire popcount32_0itb_core_128;
  wire popcount32_0itb_core_130;
  wire popcount32_0itb_core_131;
  wire popcount32_0itb_core_132;
  wire popcount32_0itb_core_133;
  wire popcount32_0itb_core_134;
  wire popcount32_0itb_core_135;
  wire popcount32_0itb_core_136;
  wire popcount32_0itb_core_139;
  wire popcount32_0itb_core_140;
  wire popcount32_0itb_core_141;
  wire popcount32_0itb_core_142;
  wire popcount32_0itb_core_143_not;
  wire popcount32_0itb_core_145;
  wire popcount32_0itb_core_146;
  wire popcount32_0itb_core_147;
  wire popcount32_0itb_core_157;
  wire popcount32_0itb_core_158;
  wire popcount32_0itb_core_160;
  wire popcount32_0itb_core_162;
  wire popcount32_0itb_core_163;
  wire popcount32_0itb_core_165;
  wire popcount32_0itb_core_166;
  wire popcount32_0itb_core_167;
  wire popcount32_0itb_core_169;
  wire popcount32_0itb_core_170;
  wire popcount32_0itb_core_171;
  wire popcount32_0itb_core_172;
  wire popcount32_0itb_core_174;
  wire popcount32_0itb_core_175;
  wire popcount32_0itb_core_176;
  wire popcount32_0itb_core_179;
  wire popcount32_0itb_core_183;
  wire popcount32_0itb_core_186;
  wire popcount32_0itb_core_189;
  wire popcount32_0itb_core_190;
  wire popcount32_0itb_core_194;
  wire popcount32_0itb_core_195;
  wire popcount32_0itb_core_196;
  wire popcount32_0itb_core_197;
  wire popcount32_0itb_core_198;
  wire popcount32_0itb_core_203;
  wire popcount32_0itb_core_204;
  wire popcount32_0itb_core_205;
  wire popcount32_0itb_core_206;
  wire popcount32_0itb_core_208;
  wire popcount32_0itb_core_210;
  wire popcount32_0itb_core_211;
  wire popcount32_0itb_core_212;
  wire popcount32_0itb_core_213;
  wire popcount32_0itb_core_214;
  wire popcount32_0itb_core_215;
  wire popcount32_0itb_core_216;
  wire popcount32_0itb_core_217;
  wire popcount32_0itb_core_218;
  wire popcount32_0itb_core_219;
  wire popcount32_0itb_core_220;
  wire popcount32_0itb_core_221;
  wire popcount32_0itb_core_222;

  assign popcount32_0itb_core_034 = ~(input_a[21] ^ input_a[2]);
  assign popcount32_0itb_core_036 = ~(input_a[25] ^ input_a[26]);
  assign popcount32_0itb_core_037 = input_a[2] & input_a[24];
  assign popcount32_0itb_core_038 = input_a[28] | input_a[0];
  assign popcount32_0itb_core_041 = input_a[9] ^ input_a[13];
  assign popcount32_0itb_core_044_not = ~input_a[24];
  assign popcount32_0itb_core_045 = input_a[28] | input_a[3];
  assign popcount32_0itb_core_046 = input_a[13] & input_a[27];
  assign popcount32_0itb_core_048 = input_a[14] & input_a[9];
  assign popcount32_0itb_core_049 = input_a[26] | input_a[25];
  assign popcount32_0itb_core_050 = input_a[3] & input_a[8];
  assign popcount32_0itb_core_051 = popcount32_0itb_core_046 | popcount32_0itb_core_048;
  assign popcount32_0itb_core_053 = popcount32_0itb_core_051 | popcount32_0itb_core_050;
  assign popcount32_0itb_core_055 = ~(input_a[26] ^ input_a[13]);
  assign popcount32_0itb_core_056 = ~(input_a[15] ^ input_a[28]);
  assign popcount32_0itb_core_058 = popcount32_0itb_core_037 ^ popcount32_0itb_core_053;
  assign popcount32_0itb_core_059 = popcount32_0itb_core_037 & popcount32_0itb_core_053;
  assign popcount32_0itb_core_060 = popcount32_0itb_core_058 ^ popcount32_0itb_core_038;
  assign popcount32_0itb_core_061 = popcount32_0itb_core_058 & popcount32_0itb_core_038;
  assign popcount32_0itb_core_062 = popcount32_0itb_core_059 | popcount32_0itb_core_061;
  assign popcount32_0itb_core_064 = input_a[27] ^ input_a[28];
  assign popcount32_0itb_core_067 = ~(input_a[10] | input_a[15]);
  assign popcount32_0itb_core_068 = input_a[7] ^ input_a[0];
  assign popcount32_0itb_core_069 = input_a[5] & input_a[31];
  assign popcount32_0itb_core_070 = ~input_a[10];
  assign popcount32_0itb_core_071 = ~(input_a[11] ^ input_a[3]);
  assign popcount32_0itb_core_072 = input_a[29] & input_a[13];
  assign popcount32_0itb_core_073 = input_a[19] & popcount32_0itb_core_070;
  assign popcount32_0itb_core_074 = popcount32_0itb_core_069 ^ input_a[10];
  assign popcount32_0itb_core_075 = popcount32_0itb_core_069 & input_a[10];
  assign popcount32_0itb_core_076 = popcount32_0itb_core_074 | popcount32_0itb_core_073;
  assign popcount32_0itb_core_080 = ~(input_a[31] ^ input_a[11]);
  assign popcount32_0itb_core_081 = ~input_a[26];
  assign popcount32_0itb_core_082 = ~(input_a[13] & input_a[23]);
  assign popcount32_0itb_core_083 = ~(input_a[6] | input_a[27]);
  assign popcount32_0itb_core_086 = input_a[5] ^ input_a[31];
  assign popcount32_0itb_core_087 = input_a[1] | input_a[26];
  assign popcount32_0itb_core_088 = input_a[10] | input_a[12];
  assign popcount32_0itb_core_089_not = ~input_a[0];
  assign popcount32_0itb_core_091 = ~(input_a[26] & input_a[4]);
  assign popcount32_0itb_core_092 = ~(popcount32_0itb_core_076 & popcount32_0itb_core_087);
  assign popcount32_0itb_core_093 = popcount32_0itb_core_076 & popcount32_0itb_core_087;
  assign popcount32_0itb_core_095 = input_a[10] | input_a[6];
  assign popcount32_0itb_core_099 = popcount32_0itb_core_075 | popcount32_0itb_core_093;
  assign popcount32_0itb_core_100 = ~(input_a[16] | input_a[4]);
  assign popcount32_0itb_core_101 = ~(input_a[3] & input_a[21]);
  assign popcount32_0itb_core_103 = input_a[25] & input_a[17];
  assign popcount32_0itb_core_104 = popcount32_0itb_core_060 ^ popcount32_0itb_core_092;
  assign popcount32_0itb_core_105 = popcount32_0itb_core_060 & popcount32_0itb_core_092;
  assign popcount32_0itb_core_106 = popcount32_0itb_core_104 ^ popcount32_0itb_core_103;
  assign popcount32_0itb_core_107 = popcount32_0itb_core_104 & popcount32_0itb_core_103;
  assign popcount32_0itb_core_108 = popcount32_0itb_core_105 | popcount32_0itb_core_107;
  assign popcount32_0itb_core_109 = popcount32_0itb_core_062 ^ popcount32_0itb_core_099;
  assign popcount32_0itb_core_110 = popcount32_0itb_core_062 & popcount32_0itb_core_099;
  assign popcount32_0itb_core_111 = popcount32_0itb_core_109 ^ popcount32_0itb_core_108;
  assign popcount32_0itb_core_112 = popcount32_0itb_core_109 & popcount32_0itb_core_108;
  assign popcount32_0itb_core_113 = popcount32_0itb_core_110 | popcount32_0itb_core_112;
  assign popcount32_0itb_core_115 = input_a[27] ^ input_a[18];
  assign popcount32_0itb_core_117 = ~input_a[26];
  assign popcount32_0itb_core_118_not = ~input_a[27];
  assign popcount32_0itb_core_119 = ~input_a[22];
  assign popcount32_0itb_core_120 = ~(input_a[18] ^ input_a[18]);
  assign popcount32_0itb_core_121 = input_a[7] ^ input_a[2];
  assign popcount32_0itb_core_123 = input_a[24] & input_a[7];
  assign popcount32_0itb_core_128 = input_a[6] & input_a[3];
  assign popcount32_0itb_core_130 = ~(input_a[26] | input_a[14]);
  assign popcount32_0itb_core_131 = input_a[4] & input_a[21];
  assign popcount32_0itb_core_132 = input_a[5] & input_a[31];
  assign popcount32_0itb_core_133 = input_a[15] & input_a[11];
  assign popcount32_0itb_core_134 = ~input_a[24];
  assign popcount32_0itb_core_135 = input_a[28] ^ input_a[28];
  assign popcount32_0itb_core_136 = popcount32_0itb_core_131 | popcount32_0itb_core_133;
  assign popcount32_0itb_core_139 = ~input_a[12];
  assign popcount32_0itb_core_140 = ~(input_a[2] ^ input_a[14]);
  assign popcount32_0itb_core_141 = ~(input_a[30] ^ input_a[5]);
  assign popcount32_0itb_core_142 = input_a[20] & input_a[22];
  assign popcount32_0itb_core_143_not = ~popcount32_0itb_core_136;
  assign popcount32_0itb_core_145 = popcount32_0itb_core_143_not ^ popcount32_0itb_core_142;
  assign popcount32_0itb_core_146 = input_a[20] & input_a[22];
  assign popcount32_0itb_core_147 = popcount32_0itb_core_136 | popcount32_0itb_core_146;
  assign popcount32_0itb_core_157 = input_a[2] | input_a[9];
  assign popcount32_0itb_core_158 = input_a[8] ^ input_a[19];
  assign popcount32_0itb_core_160 = ~(input_a[14] & input_a[16]);
  assign popcount32_0itb_core_162 = input_a[9] & input_a[26];
  assign popcount32_0itb_core_163 = ~input_a[3];
  assign popcount32_0itb_core_165 = input_a[23] & input_a[7];
  assign popcount32_0itb_core_166 = ~input_a[27];
  assign popcount32_0itb_core_167 = input_a[30] & input_a[29];
  assign popcount32_0itb_core_169 = input_a[16] & input_a[6];
  assign popcount32_0itb_core_170 = popcount32_0itb_core_165 | popcount32_0itb_core_167;
  assign popcount32_0itb_core_171 = input_a[13] ^ input_a[25];
  assign popcount32_0itb_core_172 = popcount32_0itb_core_170 | popcount32_0itb_core_169;
  assign popcount32_0itb_core_174 = ~(input_a[26] | input_a[15]);
  assign popcount32_0itb_core_175 = input_a[31] ^ input_a[22];
  assign popcount32_0itb_core_176 = ~(input_a[9] ^ input_a[25]);
  assign popcount32_0itb_core_179 = ~popcount32_0itb_core_172;
  assign popcount32_0itb_core_183 = ~(input_a[1] ^ input_a[29]);
  assign popcount32_0itb_core_186 = ~(input_a[22] & input_a[29]);
  assign popcount32_0itb_core_189 = popcount32_0itb_core_145 ^ popcount32_0itb_core_179;
  assign popcount32_0itb_core_190 = popcount32_0itb_core_145 & popcount32_0itb_core_179;
  assign popcount32_0itb_core_194 = popcount32_0itb_core_147 ^ popcount32_0itb_core_172;
  assign popcount32_0itb_core_195 = popcount32_0itb_core_147 & popcount32_0itb_core_172;
  assign popcount32_0itb_core_196 = popcount32_0itb_core_194 ^ popcount32_0itb_core_190;
  assign popcount32_0itb_core_197 = popcount32_0itb_core_194 & popcount32_0itb_core_190;
  assign popcount32_0itb_core_198 = popcount32_0itb_core_195 | popcount32_0itb_core_197;
  assign popcount32_0itb_core_203 = ~input_a[11];
  assign popcount32_0itb_core_204 = ~(input_a[29] | input_a[7]);
  assign popcount32_0itb_core_205 = input_a[31] ^ input_a[2];
  assign popcount32_0itb_core_206 = popcount32_0itb_core_106 ^ popcount32_0itb_core_189;
  assign popcount32_0itb_core_208 = ~popcount32_0itb_core_206;
  assign popcount32_0itb_core_210 = popcount32_0itb_core_106 | popcount32_0itb_core_206;
  assign popcount32_0itb_core_211 = popcount32_0itb_core_111 ^ popcount32_0itb_core_196;
  assign popcount32_0itb_core_212 = popcount32_0itb_core_111 & popcount32_0itb_core_196;
  assign popcount32_0itb_core_213 = popcount32_0itb_core_211 ^ popcount32_0itb_core_210;
  assign popcount32_0itb_core_214 = popcount32_0itb_core_211 & popcount32_0itb_core_210;
  assign popcount32_0itb_core_215 = popcount32_0itb_core_212 | popcount32_0itb_core_214;
  assign popcount32_0itb_core_216 = popcount32_0itb_core_113 ^ popcount32_0itb_core_198;
  assign popcount32_0itb_core_217 = popcount32_0itb_core_113 & popcount32_0itb_core_198;
  assign popcount32_0itb_core_218 = popcount32_0itb_core_216 ^ popcount32_0itb_core_215;
  assign popcount32_0itb_core_219 = popcount32_0itb_core_216 & popcount32_0itb_core_215;
  assign popcount32_0itb_core_220 = popcount32_0itb_core_217 | popcount32_0itb_core_219;
  assign popcount32_0itb_core_221 = ~(input_a[17] | input_a[4]);
  assign popcount32_0itb_core_222 = input_a[14] & input_a[9];

  assign popcount32_0itb_out[0] = popcount32_0itb_core_218;
  assign popcount32_0itb_out[1] = popcount32_0itb_core_208;
  assign popcount32_0itb_out[2] = popcount32_0itb_core_213;
  assign popcount32_0itb_out[3] = popcount32_0itb_core_218;
  assign popcount32_0itb_out[4] = popcount32_0itb_core_220;
  assign popcount32_0itb_out[5] = 1'b0;
endmodule