// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.19996
// WCE=10.0
// EP=0.996658%
// Printed PDK parameters:
//  Area=19067625.0
//  Delay=40574652.0
//  Power=848140.0

module popcount20_bv09(input [19:0] input_a, output [4:0] popcount20_bv09_out);
  wire popcount20_bv09_core_022_not;
  wire popcount20_bv09_core_023;
  wire popcount20_bv09_core_024;
  wire popcount20_bv09_core_025;
  wire popcount20_bv09_core_026_not;
  wire popcount20_bv09_core_027;
  wire popcount20_bv09_core_028;
  wire popcount20_bv09_core_029;
  wire popcount20_bv09_core_031;
  wire popcount20_bv09_core_033;
  wire popcount20_bv09_core_036;
  wire popcount20_bv09_core_038;
  wire popcount20_bv09_core_045;
  wire popcount20_bv09_core_046;
  wire popcount20_bv09_core_047;
  wire popcount20_bv09_core_048;
  wire popcount20_bv09_core_049;
  wire popcount20_bv09_core_050;
  wire popcount20_bv09_core_054;
  wire popcount20_bv09_core_055;
  wire popcount20_bv09_core_056;
  wire popcount20_bv09_core_057;
  wire popcount20_bv09_core_058;
  wire popcount20_bv09_core_059;
  wire popcount20_bv09_core_061;
  wire popcount20_bv09_core_066;
  wire popcount20_bv09_core_068;
  wire popcount20_bv09_core_070;
  wire popcount20_bv09_core_071;
  wire popcount20_bv09_core_072;
  wire popcount20_bv09_core_073;
  wire popcount20_bv09_core_074;
  wire popcount20_bv09_core_076;
  wire popcount20_bv09_core_077;
  wire popcount20_bv09_core_083;
  wire popcount20_bv09_core_084;
  wire popcount20_bv09_core_086;
  wire popcount20_bv09_core_090;
  wire popcount20_bv09_core_091;
  wire popcount20_bv09_core_092;
  wire popcount20_bv09_core_093;
  wire popcount20_bv09_core_095;
  wire popcount20_bv09_core_096;
  wire popcount20_bv09_core_099;
  wire popcount20_bv09_core_100;
  wire popcount20_bv09_core_101;
  wire popcount20_bv09_core_102;
  wire popcount20_bv09_core_103;
  wire popcount20_bv09_core_104;
  wire popcount20_bv09_core_107;
  wire popcount20_bv09_core_108;
  wire popcount20_bv09_core_111;
  wire popcount20_bv09_core_112;
  wire popcount20_bv09_core_114;
  wire popcount20_bv09_core_115;
  wire popcount20_bv09_core_116;
  wire popcount20_bv09_core_117;
  wire popcount20_bv09_core_118;
  wire popcount20_bv09_core_120;
  wire popcount20_bv09_core_122;
  wire popcount20_bv09_core_124;
  wire popcount20_bv09_core_125;
  wire popcount20_bv09_core_128;
  wire popcount20_bv09_core_129;
  wire popcount20_bv09_core_131;
  wire popcount20_bv09_core_132;
  wire popcount20_bv09_core_133;
  wire popcount20_bv09_core_134;
  wire popcount20_bv09_core_135;
  wire popcount20_bv09_core_137;
  wire popcount20_bv09_core_138;
  wire popcount20_bv09_core_140;
  wire popcount20_bv09_core_141;
  wire popcount20_bv09_core_142;
  wire popcount20_bv09_core_143;
  wire popcount20_bv09_core_144;

  assign popcount20_bv09_core_022_not = ~input_a[19];
  assign popcount20_bv09_core_023 = input_a[8] ^ input_a[2];
  assign popcount20_bv09_core_024 = input_a[14] ^ input_a[2];
  assign popcount20_bv09_core_025 = input_a[11] ^ input_a[13];
  assign popcount20_bv09_core_026_not = ~input_a[5];
  assign popcount20_bv09_core_027 = ~(input_a[7] & input_a[6]);
  assign popcount20_bv09_core_028 = ~(input_a[6] | input_a[6]);
  assign popcount20_bv09_core_029 = input_a[19] ^ input_a[7];
  assign popcount20_bv09_core_031 = ~(input_a[15] | input_a[7]);
  assign popcount20_bv09_core_033 = ~(input_a[7] & input_a[13]);
  assign popcount20_bv09_core_036 = input_a[9] ^ input_a[6];
  assign popcount20_bv09_core_038 = input_a[12] | input_a[10];
  assign popcount20_bv09_core_045 = input_a[13] | input_a[8];
  assign popcount20_bv09_core_046 = input_a[0] & input_a[10];
  assign popcount20_bv09_core_047 = ~(input_a[7] | input_a[14]);
  assign popcount20_bv09_core_048 = ~(input_a[17] ^ input_a[11]);
  assign popcount20_bv09_core_049 = ~(input_a[1] | input_a[14]);
  assign popcount20_bv09_core_050 = input_a[12] & input_a[13];
  assign popcount20_bv09_core_054 = popcount20_bv09_core_046 | popcount20_bv09_core_050;
  assign popcount20_bv09_core_055 = ~(input_a[12] & input_a[13]);
  assign popcount20_bv09_core_056 = ~input_a[19];
  assign popcount20_bv09_core_057 = input_a[0] | input_a[14];
  assign popcount20_bv09_core_058 = ~input_a[6];
  assign popcount20_bv09_core_059 = ~input_a[2];
  assign popcount20_bv09_core_061 = input_a[15] & input_a[14];
  assign popcount20_bv09_core_066 = ~(input_a[5] ^ input_a[0]);
  assign popcount20_bv09_core_068 = ~(input_a[15] ^ input_a[14]);
  assign popcount20_bv09_core_070 = input_a[8] & input_a[8];
  assign popcount20_bv09_core_071 = input_a[9] & input_a[14];
  assign popcount20_bv09_core_072 = input_a[15] & input_a[2];
  assign popcount20_bv09_core_073 = input_a[7] | input_a[15];
  assign popcount20_bv09_core_074 = input_a[14] & input_a[3];
  assign popcount20_bv09_core_076 = input_a[11] & input_a[8];
  assign popcount20_bv09_core_077 = ~input_a[7];
  assign popcount20_bv09_core_083 = ~input_a[18];
  assign popcount20_bv09_core_084 = popcount20_bv09_core_074 & popcount20_bv09_core_076;
  assign popcount20_bv09_core_086 = ~input_a[13];
  assign popcount20_bv09_core_090 = input_a[15] ^ input_a[16];
  assign popcount20_bv09_core_091 = input_a[15] & input_a[16];
  assign popcount20_bv09_core_092 = ~(input_a[8] ^ input_a[9]);
  assign popcount20_bv09_core_093 = input_a[18] & input_a[19];
  assign popcount20_bv09_core_095 = input_a[17] & input_a[6];
  assign popcount20_bv09_core_096 = popcount20_bv09_core_093 | popcount20_bv09_core_095;
  assign popcount20_bv09_core_099 = popcount20_bv09_core_090 & input_a[9];
  assign popcount20_bv09_core_100 = popcount20_bv09_core_091 ^ popcount20_bv09_core_096;
  assign popcount20_bv09_core_101 = popcount20_bv09_core_091 & popcount20_bv09_core_096;
  assign popcount20_bv09_core_102 = popcount20_bv09_core_100 ^ popcount20_bv09_core_099;
  assign popcount20_bv09_core_103 = popcount20_bv09_core_100 & popcount20_bv09_core_099;
  assign popcount20_bv09_core_104 = popcount20_bv09_core_101 | popcount20_bv09_core_103;
  assign popcount20_bv09_core_107 = input_a[6] ^ input_a[16];
  assign popcount20_bv09_core_108 = input_a[5] & input_a[1];
  assign popcount20_bv09_core_111 = popcount20_bv09_core_102 ^ popcount20_bv09_core_108;
  assign popcount20_bv09_core_112 = popcount20_bv09_core_102 & popcount20_bv09_core_108;
  assign popcount20_bv09_core_114 = popcount20_bv09_core_084 ^ popcount20_bv09_core_104;
  assign popcount20_bv09_core_115 = popcount20_bv09_core_084 & popcount20_bv09_core_104;
  assign popcount20_bv09_core_116 = popcount20_bv09_core_114 ^ popcount20_bv09_core_112;
  assign popcount20_bv09_core_117 = popcount20_bv09_core_114 & popcount20_bv09_core_112;
  assign popcount20_bv09_core_118 = popcount20_bv09_core_115 | popcount20_bv09_core_117;
  assign popcount20_bv09_core_120 = input_a[16] ^ input_a[6];
  assign popcount20_bv09_core_122 = ~(input_a[17] | input_a[4]);
  assign popcount20_bv09_core_124 = ~input_a[12];
  assign popcount20_bv09_core_125 = input_a[4] & input_a[7];
  assign popcount20_bv09_core_128 = popcount20_bv09_core_111 ^ popcount20_bv09_core_125;
  assign popcount20_bv09_core_129 = popcount20_bv09_core_111 & popcount20_bv09_core_125;
  assign popcount20_bv09_core_131 = popcount20_bv09_core_054 ^ popcount20_bv09_core_116;
  assign popcount20_bv09_core_132 = popcount20_bv09_core_054 & popcount20_bv09_core_116;
  assign popcount20_bv09_core_133 = popcount20_bv09_core_131 ^ popcount20_bv09_core_129;
  assign popcount20_bv09_core_134 = popcount20_bv09_core_131 & popcount20_bv09_core_129;
  assign popcount20_bv09_core_135 = popcount20_bv09_core_132 | popcount20_bv09_core_134;
  assign popcount20_bv09_core_137 = input_a[11] & popcount20_bv09_core_118;
  assign popcount20_bv09_core_138 = input_a[8] ^ input_a[7];
  assign popcount20_bv09_core_140 = popcount20_bv09_core_137 | popcount20_bv09_core_135;
  assign popcount20_bv09_core_141 = ~(input_a[17] | input_a[6]);
  assign popcount20_bv09_core_142 = input_a[15] | input_a[13];
  assign popcount20_bv09_core_143 = input_a[12] ^ input_a[5];
  assign popcount20_bv09_core_144 = input_a[13] | input_a[16];

  assign popcount20_bv09_out[0] = input_a[2];
  assign popcount20_bv09_out[1] = popcount20_bv09_core_128;
  assign popcount20_bv09_out[2] = popcount20_bv09_core_133;
  assign popcount20_bv09_out[3] = 1'b0;
  assign popcount20_bv09_out[4] = popcount20_bv09_core_140;
endmodule