// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.50741
// WCE=20.0
// EP=0.874629%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount40_txyt(input [39:0] input_a, output [5:0] popcount40_txyt_out);
  wire popcount40_txyt_core_043;
  wire popcount40_txyt_core_044;
  wire popcount40_txyt_core_048;
  wire popcount40_txyt_core_050;
  wire popcount40_txyt_core_051;
  wire popcount40_txyt_core_053;
  wire popcount40_txyt_core_055;
  wire popcount40_txyt_core_056;
  wire popcount40_txyt_core_057;
  wire popcount40_txyt_core_058;
  wire popcount40_txyt_core_059;
  wire popcount40_txyt_core_061;
  wire popcount40_txyt_core_063;
  wire popcount40_txyt_core_065;
  wire popcount40_txyt_core_068;
  wire popcount40_txyt_core_071;
  wire popcount40_txyt_core_073;
  wire popcount40_txyt_core_074;
  wire popcount40_txyt_core_075;
  wire popcount40_txyt_core_076;
  wire popcount40_txyt_core_077;
  wire popcount40_txyt_core_078;
  wire popcount40_txyt_core_081;
  wire popcount40_txyt_core_083;
  wire popcount40_txyt_core_084;
  wire popcount40_txyt_core_086;
  wire popcount40_txyt_core_087;
  wire popcount40_txyt_core_089;
  wire popcount40_txyt_core_090_not;
  wire popcount40_txyt_core_091;
  wire popcount40_txyt_core_092;
  wire popcount40_txyt_core_094;
  wire popcount40_txyt_core_095;
  wire popcount40_txyt_core_099;
  wire popcount40_txyt_core_100;
  wire popcount40_txyt_core_101;
  wire popcount40_txyt_core_103;
  wire popcount40_txyt_core_104;
  wire popcount40_txyt_core_106;
  wire popcount40_txyt_core_108;
  wire popcount40_txyt_core_109;
  wire popcount40_txyt_core_110;
  wire popcount40_txyt_core_111;
  wire popcount40_txyt_core_112;
  wire popcount40_txyt_core_113;
  wire popcount40_txyt_core_114;
  wire popcount40_txyt_core_115;
  wire popcount40_txyt_core_116;
  wire popcount40_txyt_core_117;
  wire popcount40_txyt_core_118;
  wire popcount40_txyt_core_119;
  wire popcount40_txyt_core_120_not;
  wire popcount40_txyt_core_122;
  wire popcount40_txyt_core_123;
  wire popcount40_txyt_core_124;
  wire popcount40_txyt_core_125;
  wire popcount40_txyt_core_126_not;
  wire popcount40_txyt_core_128;
  wire popcount40_txyt_core_130;
  wire popcount40_txyt_core_132;
  wire popcount40_txyt_core_133;
  wire popcount40_txyt_core_135;
  wire popcount40_txyt_core_136;
  wire popcount40_txyt_core_138;
  wire popcount40_txyt_core_139;
  wire popcount40_txyt_core_141;
  wire popcount40_txyt_core_142;
  wire popcount40_txyt_core_144;
  wire popcount40_txyt_core_145;
  wire popcount40_txyt_core_146;
  wire popcount40_txyt_core_147;
  wire popcount40_txyt_core_152;
  wire popcount40_txyt_core_153;
  wire popcount40_txyt_core_155;
  wire popcount40_txyt_core_156;
  wire popcount40_txyt_core_157_not;
  wire popcount40_txyt_core_158;
  wire popcount40_txyt_core_159;
  wire popcount40_txyt_core_161;
  wire popcount40_txyt_core_162;
  wire popcount40_txyt_core_164;
  wire popcount40_txyt_core_165;
  wire popcount40_txyt_core_166;
  wire popcount40_txyt_core_167;
  wire popcount40_txyt_core_169;
  wire popcount40_txyt_core_172;
  wire popcount40_txyt_core_173;
  wire popcount40_txyt_core_174;
  wire popcount40_txyt_core_175;
  wire popcount40_txyt_core_176;
  wire popcount40_txyt_core_177;
  wire popcount40_txyt_core_178;
  wire popcount40_txyt_core_180;
  wire popcount40_txyt_core_181;
  wire popcount40_txyt_core_182;
  wire popcount40_txyt_core_183;
  wire popcount40_txyt_core_184;
  wire popcount40_txyt_core_186;
  wire popcount40_txyt_core_187;
  wire popcount40_txyt_core_190;
  wire popcount40_txyt_core_194;
  wire popcount40_txyt_core_195;
  wire popcount40_txyt_core_196;
  wire popcount40_txyt_core_198_not;
  wire popcount40_txyt_core_199;
  wire popcount40_txyt_core_200;
  wire popcount40_txyt_core_202;
  wire popcount40_txyt_core_203;
  wire popcount40_txyt_core_204;
  wire popcount40_txyt_core_205;
  wire popcount40_txyt_core_206;
  wire popcount40_txyt_core_207;
  wire popcount40_txyt_core_208;
  wire popcount40_txyt_core_210;
  wire popcount40_txyt_core_211;
  wire popcount40_txyt_core_212;
  wire popcount40_txyt_core_213;
  wire popcount40_txyt_core_214;
  wire popcount40_txyt_core_215;
  wire popcount40_txyt_core_216;
  wire popcount40_txyt_core_219;
  wire popcount40_txyt_core_222;
  wire popcount40_txyt_core_223;
  wire popcount40_txyt_core_225;
  wire popcount40_txyt_core_226;
  wire popcount40_txyt_core_227;
  wire popcount40_txyt_core_229;
  wire popcount40_txyt_core_230;
  wire popcount40_txyt_core_231;
  wire popcount40_txyt_core_232;
  wire popcount40_txyt_core_234;
  wire popcount40_txyt_core_235;
  wire popcount40_txyt_core_236;
  wire popcount40_txyt_core_238;
  wire popcount40_txyt_core_239;
  wire popcount40_txyt_core_240;
  wire popcount40_txyt_core_241;
  wire popcount40_txyt_core_242;
  wire popcount40_txyt_core_244;
  wire popcount40_txyt_core_245;
  wire popcount40_txyt_core_246;
  wire popcount40_txyt_core_248;
  wire popcount40_txyt_core_251;
  wire popcount40_txyt_core_252;
  wire popcount40_txyt_core_254;
  wire popcount40_txyt_core_255;
  wire popcount40_txyt_core_256;
  wire popcount40_txyt_core_257;
  wire popcount40_txyt_core_260;
  wire popcount40_txyt_core_261;
  wire popcount40_txyt_core_262;
  wire popcount40_txyt_core_263;
  wire popcount40_txyt_core_264;
  wire popcount40_txyt_core_266;
  wire popcount40_txyt_core_267;
  wire popcount40_txyt_core_269;
  wire popcount40_txyt_core_271;
  wire popcount40_txyt_core_272;
  wire popcount40_txyt_core_274;
  wire popcount40_txyt_core_275;
  wire popcount40_txyt_core_276;
  wire popcount40_txyt_core_277;
  wire popcount40_txyt_core_278;
  wire popcount40_txyt_core_280;
  wire popcount40_txyt_core_282;
  wire popcount40_txyt_core_283;
  wire popcount40_txyt_core_285;
  wire popcount40_txyt_core_286;
  wire popcount40_txyt_core_287;
  wire popcount40_txyt_core_289;
  wire popcount40_txyt_core_290;
  wire popcount40_txyt_core_292;
  wire popcount40_txyt_core_293;
  wire popcount40_txyt_core_294;
  wire popcount40_txyt_core_295;
  wire popcount40_txyt_core_296;
  wire popcount40_txyt_core_298;
  wire popcount40_txyt_core_300;
  wire popcount40_txyt_core_303;
  wire popcount40_txyt_core_304;
  wire popcount40_txyt_core_305;
  wire popcount40_txyt_core_306;
  wire popcount40_txyt_core_307;
  wire popcount40_txyt_core_308;
  wire popcount40_txyt_core_309;
  wire popcount40_txyt_core_310;
  wire popcount40_txyt_core_311;
  wire popcount40_txyt_core_312;
  wire popcount40_txyt_core_313;
  wire popcount40_txyt_core_314;
  wire popcount40_txyt_core_316;

  assign popcount40_txyt_core_043 = ~input_a[27];
  assign popcount40_txyt_core_044 = input_a[20] & input_a[21];
  assign popcount40_txyt_core_048 = input_a[9] ^ input_a[14];
  assign popcount40_txyt_core_050 = input_a[22] | input_a[3];
  assign popcount40_txyt_core_051 = input_a[29] ^ input_a[9];
  assign popcount40_txyt_core_053 = ~(input_a[33] | input_a[2]);
  assign popcount40_txyt_core_055 = ~(input_a[1] | input_a[38]);
  assign popcount40_txyt_core_056 = input_a[5] | input_a[39];
  assign popcount40_txyt_core_057 = ~input_a[15];
  assign popcount40_txyt_core_058 = ~(input_a[3] | input_a[21]);
  assign popcount40_txyt_core_059 = input_a[22] & input_a[6];
  assign popcount40_txyt_core_061 = ~(input_a[29] ^ input_a[39]);
  assign popcount40_txyt_core_063 = input_a[24] & input_a[36];
  assign popcount40_txyt_core_065 = ~(input_a[3] & input_a[35]);
  assign popcount40_txyt_core_068 = input_a[35] & input_a[6];
  assign popcount40_txyt_core_071 = input_a[22] ^ input_a[11];
  assign popcount40_txyt_core_073 = ~(input_a[8] | input_a[13]);
  assign popcount40_txyt_core_074 = ~(input_a[18] & input_a[6]);
  assign popcount40_txyt_core_075 = ~(input_a[37] ^ input_a[4]);
  assign popcount40_txyt_core_076 = ~(input_a[11] & input_a[28]);
  assign popcount40_txyt_core_077 = ~input_a[5];
  assign popcount40_txyt_core_078 = input_a[0] | input_a[39];
  assign popcount40_txyt_core_081 = input_a[31] & input_a[27];
  assign popcount40_txyt_core_083 = ~(input_a[2] & input_a[5]);
  assign popcount40_txyt_core_084 = ~input_a[38];
  assign popcount40_txyt_core_086 = ~(input_a[21] ^ input_a[31]);
  assign popcount40_txyt_core_087 = ~(input_a[36] & input_a[17]);
  assign popcount40_txyt_core_089 = input_a[1] ^ input_a[10];
  assign popcount40_txyt_core_090_not = ~input_a[12];
  assign popcount40_txyt_core_091 = ~(input_a[10] ^ input_a[3]);
  assign popcount40_txyt_core_092 = ~input_a[23];
  assign popcount40_txyt_core_094 = input_a[6] ^ input_a[22];
  assign popcount40_txyt_core_095 = ~(input_a[5] ^ input_a[15]);
  assign popcount40_txyt_core_099 = input_a[27] | input_a[34];
  assign popcount40_txyt_core_100 = input_a[36] ^ input_a[9];
  assign popcount40_txyt_core_101 = input_a[3] & input_a[38];
  assign popcount40_txyt_core_103 = input_a[8] & input_a[30];
  assign popcount40_txyt_core_104 = ~(input_a[31] ^ input_a[13]);
  assign popcount40_txyt_core_106 = ~(input_a[9] | input_a[5]);
  assign popcount40_txyt_core_108 = input_a[25] | input_a[35];
  assign popcount40_txyt_core_109 = input_a[32] & input_a[9];
  assign popcount40_txyt_core_110 = ~(input_a[10] | input_a[12]);
  assign popcount40_txyt_core_111 = ~(input_a[5] | input_a[37]);
  assign popcount40_txyt_core_112 = ~(input_a[25] & input_a[15]);
  assign popcount40_txyt_core_113 = ~input_a[24];
  assign popcount40_txyt_core_114 = ~input_a[27];
  assign popcount40_txyt_core_115 = ~(input_a[13] ^ input_a[15]);
  assign popcount40_txyt_core_116 = ~(input_a[12] & input_a[16]);
  assign popcount40_txyt_core_117 = input_a[16] | input_a[1];
  assign popcount40_txyt_core_118 = ~(input_a[28] ^ input_a[21]);
  assign popcount40_txyt_core_119 = input_a[31] | input_a[25];
  assign popcount40_txyt_core_120_not = ~input_a[25];
  assign popcount40_txyt_core_122 = input_a[22] & input_a[37];
  assign popcount40_txyt_core_123 = ~input_a[33];
  assign popcount40_txyt_core_124 = input_a[6] ^ input_a[4];
  assign popcount40_txyt_core_125 = ~input_a[34];
  assign popcount40_txyt_core_126_not = ~input_a[9];
  assign popcount40_txyt_core_128 = input_a[39] | input_a[15];
  assign popcount40_txyt_core_130 = ~input_a[31];
  assign popcount40_txyt_core_132 = ~(input_a[12] | input_a[10]);
  assign popcount40_txyt_core_133 = ~(input_a[36] & input_a[10]);
  assign popcount40_txyt_core_135 = ~(input_a[5] ^ input_a[25]);
  assign popcount40_txyt_core_136 = ~(input_a[28] | input_a[32]);
  assign popcount40_txyt_core_138 = input_a[20] | input_a[21];
  assign popcount40_txyt_core_139 = input_a[15] & input_a[28];
  assign popcount40_txyt_core_141 = ~(input_a[29] ^ input_a[23]);
  assign popcount40_txyt_core_142 = input_a[11] & input_a[0];
  assign popcount40_txyt_core_144 = input_a[33] & input_a[13];
  assign popcount40_txyt_core_145 = input_a[0] | input_a[24];
  assign popcount40_txyt_core_146 = ~(input_a[33] ^ input_a[0]);
  assign popcount40_txyt_core_147 = input_a[7] ^ input_a[20];
  assign popcount40_txyt_core_152 = ~input_a[7];
  assign popcount40_txyt_core_153 = ~(input_a[26] & input_a[30]);
  assign popcount40_txyt_core_155 = input_a[0] ^ input_a[28];
  assign popcount40_txyt_core_156 = input_a[1] & input_a[5];
  assign popcount40_txyt_core_157_not = ~input_a[18];
  assign popcount40_txyt_core_158 = ~input_a[13];
  assign popcount40_txyt_core_159 = input_a[30] ^ input_a[8];
  assign popcount40_txyt_core_161 = ~input_a[35];
  assign popcount40_txyt_core_162 = ~(input_a[33] ^ input_a[2]);
  assign popcount40_txyt_core_164 = input_a[9] & input_a[10];
  assign popcount40_txyt_core_165 = ~(input_a[1] & input_a[18]);
  assign popcount40_txyt_core_166 = input_a[28] & input_a[1];
  assign popcount40_txyt_core_167 = ~input_a[20];
  assign popcount40_txyt_core_169 = ~(input_a[0] | input_a[11]);
  assign popcount40_txyt_core_172 = input_a[11] ^ input_a[3];
  assign popcount40_txyt_core_173 = input_a[20] ^ input_a[33];
  assign popcount40_txyt_core_174 = input_a[39] & input_a[14];
  assign popcount40_txyt_core_175 = input_a[1] & input_a[2];
  assign popcount40_txyt_core_176 = input_a[21] | input_a[23];
  assign popcount40_txyt_core_177 = input_a[39] & input_a[18];
  assign popcount40_txyt_core_178 = ~(input_a[18] | input_a[38]);
  assign popcount40_txyt_core_180 = ~input_a[39];
  assign popcount40_txyt_core_181 = ~input_a[39];
  assign popcount40_txyt_core_182 = ~input_a[26];
  assign popcount40_txyt_core_183 = ~input_a[28];
  assign popcount40_txyt_core_184 = ~(input_a[39] ^ input_a[8]);
  assign popcount40_txyt_core_186 = ~input_a[33];
  assign popcount40_txyt_core_187 = input_a[4] | input_a[32];
  assign popcount40_txyt_core_190 = input_a[35] & input_a[27];
  assign popcount40_txyt_core_194 = ~(input_a[15] ^ input_a[2]);
  assign popcount40_txyt_core_195 = ~(input_a[39] & input_a[30]);
  assign popcount40_txyt_core_196 = input_a[4] | input_a[24];
  assign popcount40_txyt_core_198_not = ~input_a[18];
  assign popcount40_txyt_core_199 = input_a[21] | input_a[19];
  assign popcount40_txyt_core_200 = ~(input_a[27] ^ input_a[22]);
  assign popcount40_txyt_core_202 = input_a[11] | input_a[33];
  assign popcount40_txyt_core_203 = input_a[10] ^ input_a[19];
  assign popcount40_txyt_core_204 = ~(input_a[17] | input_a[3]);
  assign popcount40_txyt_core_205 = input_a[32] ^ input_a[20];
  assign popcount40_txyt_core_206 = ~(input_a[21] & input_a[39]);
  assign popcount40_txyt_core_207 = ~(input_a[0] ^ input_a[3]);
  assign popcount40_txyt_core_208 = input_a[22] | input_a[6];
  assign popcount40_txyt_core_210 = ~(input_a[8] ^ input_a[35]);
  assign popcount40_txyt_core_211 = input_a[15] ^ input_a[20];
  assign popcount40_txyt_core_212 = input_a[28] ^ input_a[7];
  assign popcount40_txyt_core_213 = input_a[10] ^ input_a[38];
  assign popcount40_txyt_core_214 = input_a[24] | input_a[18];
  assign popcount40_txyt_core_215 = input_a[26] | input_a[9];
  assign popcount40_txyt_core_216 = ~(input_a[26] & input_a[34]);
  assign popcount40_txyt_core_219 = input_a[39] | input_a[30];
  assign popcount40_txyt_core_222 = input_a[21] | input_a[22];
  assign popcount40_txyt_core_223 = ~(input_a[14] ^ input_a[16]);
  assign popcount40_txyt_core_225 = input_a[9] ^ input_a[24];
  assign popcount40_txyt_core_226 = input_a[20] ^ input_a[34];
  assign popcount40_txyt_core_227 = ~(input_a[5] ^ input_a[15]);
  assign popcount40_txyt_core_229 = ~(input_a[30] | input_a[7]);
  assign popcount40_txyt_core_230 = input_a[3] & input_a[36];
  assign popcount40_txyt_core_231 = input_a[37] & input_a[12];
  assign popcount40_txyt_core_232 = input_a[2] & input_a[23];
  assign popcount40_txyt_core_234 = input_a[13] ^ input_a[7];
  assign popcount40_txyt_core_235 = ~input_a[0];
  assign popcount40_txyt_core_236 = input_a[30] & input_a[29];
  assign popcount40_txyt_core_238 = input_a[20] & input_a[28];
  assign popcount40_txyt_core_239 = ~(input_a[39] & input_a[29]);
  assign popcount40_txyt_core_240 = input_a[25] | input_a[3];
  assign popcount40_txyt_core_241 = input_a[4] | input_a[16];
  assign popcount40_txyt_core_242 = ~(input_a[26] ^ input_a[21]);
  assign popcount40_txyt_core_244 = input_a[17] ^ input_a[17];
  assign popcount40_txyt_core_245 = ~(input_a[27] & input_a[36]);
  assign popcount40_txyt_core_246 = input_a[7] | input_a[24];
  assign popcount40_txyt_core_248 = ~(input_a[1] ^ input_a[19]);
  assign popcount40_txyt_core_251 = ~(input_a[32] & input_a[38]);
  assign popcount40_txyt_core_252 = input_a[36] ^ input_a[7];
  assign popcount40_txyt_core_254 = ~input_a[34];
  assign popcount40_txyt_core_255 = input_a[17] | input_a[21];
  assign popcount40_txyt_core_256 = input_a[1] | input_a[11];
  assign popcount40_txyt_core_257 = input_a[6] & input_a[10];
  assign popcount40_txyt_core_260 = input_a[33] | input_a[5];
  assign popcount40_txyt_core_261 = ~input_a[20];
  assign popcount40_txyt_core_262 = ~(input_a[13] ^ input_a[11]);
  assign popcount40_txyt_core_263 = input_a[34] & input_a[39];
  assign popcount40_txyt_core_264 = ~(input_a[32] & input_a[28]);
  assign popcount40_txyt_core_266 = input_a[1] | input_a[32];
  assign popcount40_txyt_core_267 = input_a[38] ^ input_a[0];
  assign popcount40_txyt_core_269 = input_a[33] | input_a[36];
  assign popcount40_txyt_core_271 = ~(input_a[33] & input_a[34]);
  assign popcount40_txyt_core_272 = ~input_a[21];
  assign popcount40_txyt_core_274 = ~input_a[4];
  assign popcount40_txyt_core_275 = ~(input_a[18] & input_a[32]);
  assign popcount40_txyt_core_276 = input_a[13] ^ input_a[3];
  assign popcount40_txyt_core_277 = ~(input_a[9] ^ input_a[0]);
  assign popcount40_txyt_core_278 = input_a[38] & input_a[29];
  assign popcount40_txyt_core_280 = ~(input_a[29] | input_a[15]);
  assign popcount40_txyt_core_282 = ~input_a[21];
  assign popcount40_txyt_core_283 = input_a[22] & input_a[23];
  assign popcount40_txyt_core_285 = input_a[4] ^ input_a[17];
  assign popcount40_txyt_core_286 = ~input_a[13];
  assign popcount40_txyt_core_287 = input_a[12] ^ input_a[5];
  assign popcount40_txyt_core_289 = ~(input_a[34] & input_a[11]);
  assign popcount40_txyt_core_290 = ~(input_a[7] | input_a[26]);
  assign popcount40_txyt_core_292 = ~(input_a[31] & input_a[20]);
  assign popcount40_txyt_core_293 = input_a[35] ^ input_a[9];
  assign popcount40_txyt_core_294 = input_a[20] ^ input_a[2];
  assign popcount40_txyt_core_295 = input_a[13] | input_a[25];
  assign popcount40_txyt_core_296 = ~(input_a[9] | input_a[24]);
  assign popcount40_txyt_core_298 = ~input_a[19];
  assign popcount40_txyt_core_300 = input_a[22] | input_a[14];
  assign popcount40_txyt_core_303 = ~(input_a[22] ^ input_a[37]);
  assign popcount40_txyt_core_304 = input_a[31] ^ input_a[15];
  assign popcount40_txyt_core_305 = ~input_a[8];
  assign popcount40_txyt_core_306 = ~input_a[12];
  assign popcount40_txyt_core_307 = ~(input_a[12] & input_a[29]);
  assign popcount40_txyt_core_308 = ~(input_a[20] & input_a[11]);
  assign popcount40_txyt_core_309 = ~(input_a[26] | input_a[27]);
  assign popcount40_txyt_core_310 = ~input_a[1];
  assign popcount40_txyt_core_311 = input_a[26] | input_a[3];
  assign popcount40_txyt_core_312 = ~input_a[30];
  assign popcount40_txyt_core_313 = ~(input_a[27] | input_a[1]);
  assign popcount40_txyt_core_314 = ~(input_a[15] & input_a[13]);
  assign popcount40_txyt_core_316 = ~(input_a[27] ^ input_a[28]);

  assign popcount40_txyt_out[0] = input_a[33];
  assign popcount40_txyt_out[1] = popcount40_txyt_core_305;
  assign popcount40_txyt_out[2] = input_a[8];
  assign popcount40_txyt_out[3] = 1'b0;
  assign popcount40_txyt_out[4] = 1'b1;
  assign popcount40_txyt_out[5] = 1'b0;
endmodule