// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=9.5126
// WCE=30.0
// EP=0.993924%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_ssce(input [35:0] input_a, output [5:0] popcount36_ssce_out);
  wire popcount36_ssce_core_038;
  wire popcount36_ssce_core_039;
  wire popcount36_ssce_core_040;
  wire popcount36_ssce_core_041;
  wire popcount36_ssce_core_042;
  wire popcount36_ssce_core_046;
  wire popcount36_ssce_core_047;
  wire popcount36_ssce_core_048;
  wire popcount36_ssce_core_049;
  wire popcount36_ssce_core_050;
  wire popcount36_ssce_core_052;
  wire popcount36_ssce_core_053;
  wire popcount36_ssce_core_054;
  wire popcount36_ssce_core_056;
  wire popcount36_ssce_core_057;
  wire popcount36_ssce_core_058;
  wire popcount36_ssce_core_060;
  wire popcount36_ssce_core_062;
  wire popcount36_ssce_core_064;
  wire popcount36_ssce_core_065;
  wire popcount36_ssce_core_066;
  wire popcount36_ssce_core_068_not;
  wire popcount36_ssce_core_070;
  wire popcount36_ssce_core_071;
  wire popcount36_ssce_core_072_not;
  wire popcount36_ssce_core_074;
  wire popcount36_ssce_core_075;
  wire popcount36_ssce_core_076;
  wire popcount36_ssce_core_077;
  wire popcount36_ssce_core_078;
  wire popcount36_ssce_core_079;
  wire popcount36_ssce_core_080;
  wire popcount36_ssce_core_081;
  wire popcount36_ssce_core_085;
  wire popcount36_ssce_core_087;
  wire popcount36_ssce_core_088;
  wire popcount36_ssce_core_089;
  wire popcount36_ssce_core_090;
  wire popcount36_ssce_core_091;
  wire popcount36_ssce_core_092;
  wire popcount36_ssce_core_093;
  wire popcount36_ssce_core_097;
  wire popcount36_ssce_core_098;
  wire popcount36_ssce_core_099;
  wire popcount36_ssce_core_100;
  wire popcount36_ssce_core_111;
  wire popcount36_ssce_core_112;
  wire popcount36_ssce_core_113;
  wire popcount36_ssce_core_116;
  wire popcount36_ssce_core_118;
  wire popcount36_ssce_core_119;
  wire popcount36_ssce_core_122;
  wire popcount36_ssce_core_124;
  wire popcount36_ssce_core_125;
  wire popcount36_ssce_core_126;
  wire popcount36_ssce_core_128;
  wire popcount36_ssce_core_129;
  wire popcount36_ssce_core_130;
  wire popcount36_ssce_core_131;
  wire popcount36_ssce_core_132;
  wire popcount36_ssce_core_134;
  wire popcount36_ssce_core_135;
  wire popcount36_ssce_core_138;
  wire popcount36_ssce_core_140;
  wire popcount36_ssce_core_142;
  wire popcount36_ssce_core_143;
  wire popcount36_ssce_core_144;
  wire popcount36_ssce_core_145;
  wire popcount36_ssce_core_146;
  wire popcount36_ssce_core_147;
  wire popcount36_ssce_core_148;
  wire popcount36_ssce_core_150;
  wire popcount36_ssce_core_151;
  wire popcount36_ssce_core_152;
  wire popcount36_ssce_core_154;
  wire popcount36_ssce_core_155;
  wire popcount36_ssce_core_160;
  wire popcount36_ssce_core_161;
  wire popcount36_ssce_core_163;
  wire popcount36_ssce_core_164;
  wire popcount36_ssce_core_166;
  wire popcount36_ssce_core_167;
  wire popcount36_ssce_core_168;
  wire popcount36_ssce_core_169;
  wire popcount36_ssce_core_170;
  wire popcount36_ssce_core_171;
  wire popcount36_ssce_core_174;
  wire popcount36_ssce_core_176;
  wire popcount36_ssce_core_179;
  wire popcount36_ssce_core_181;
  wire popcount36_ssce_core_182;
  wire popcount36_ssce_core_183_not;
  wire popcount36_ssce_core_185;
  wire popcount36_ssce_core_186;
  wire popcount36_ssce_core_187;
  wire popcount36_ssce_core_189;
  wire popcount36_ssce_core_190;
  wire popcount36_ssce_core_191;
  wire popcount36_ssce_core_193;
  wire popcount36_ssce_core_195;
  wire popcount36_ssce_core_197;
  wire popcount36_ssce_core_198;
  wire popcount36_ssce_core_199;
  wire popcount36_ssce_core_201;
  wire popcount36_ssce_core_202;
  wire popcount36_ssce_core_203;
  wire popcount36_ssce_core_204;
  wire popcount36_ssce_core_208;
  wire popcount36_ssce_core_209;
  wire popcount36_ssce_core_211;
  wire popcount36_ssce_core_213;
  wire popcount36_ssce_core_214;
  wire popcount36_ssce_core_215;
  wire popcount36_ssce_core_219;
  wire popcount36_ssce_core_220;
  wire popcount36_ssce_core_222_not;
  wire popcount36_ssce_core_225;
  wire popcount36_ssce_core_226;
  wire popcount36_ssce_core_227;
  wire popcount36_ssce_core_228;
  wire popcount36_ssce_core_229;
  wire popcount36_ssce_core_230;
  wire popcount36_ssce_core_231;
  wire popcount36_ssce_core_232;
  wire popcount36_ssce_core_233;
  wire popcount36_ssce_core_236;
  wire popcount36_ssce_core_237;
  wire popcount36_ssce_core_238;
  wire popcount36_ssce_core_242;
  wire popcount36_ssce_core_243;
  wire popcount36_ssce_core_244;
  wire popcount36_ssce_core_245;
  wire popcount36_ssce_core_246;
  wire popcount36_ssce_core_247;
  wire popcount36_ssce_core_248;
  wire popcount36_ssce_core_249;
  wire popcount36_ssce_core_250;
  wire popcount36_ssce_core_251_not;
  wire popcount36_ssce_core_254;
  wire popcount36_ssce_core_255;
  wire popcount36_ssce_core_256;
  wire popcount36_ssce_core_257;
  wire popcount36_ssce_core_258;
  wire popcount36_ssce_core_260;
  wire popcount36_ssce_core_261;
  wire popcount36_ssce_core_263;
  wire popcount36_ssce_core_265;
  wire popcount36_ssce_core_267;
  wire popcount36_ssce_core_269;
  wire popcount36_ssce_core_270;
  wire popcount36_ssce_core_273;
  wire popcount36_ssce_core_274;

  assign popcount36_ssce_core_038 = input_a[9] | input_a[33];
  assign popcount36_ssce_core_039 = input_a[24] ^ input_a[27];
  assign popcount36_ssce_core_040 = input_a[23] & input_a[11];
  assign popcount36_ssce_core_041 = ~(input_a[18] & input_a[8]);
  assign popcount36_ssce_core_042 = ~(input_a[33] & input_a[10]);
  assign popcount36_ssce_core_046 = ~(input_a[15] | input_a[13]);
  assign popcount36_ssce_core_047 = input_a[18] & input_a[14];
  assign popcount36_ssce_core_048 = ~input_a[19];
  assign popcount36_ssce_core_049 = ~input_a[20];
  assign popcount36_ssce_core_050 = input_a[11] ^ input_a[30];
  assign popcount36_ssce_core_052 = ~input_a[20];
  assign popcount36_ssce_core_053 = ~(input_a[20] ^ input_a[26]);
  assign popcount36_ssce_core_054 = input_a[27] ^ input_a[34];
  assign popcount36_ssce_core_056 = input_a[31] & input_a[28];
  assign popcount36_ssce_core_057 = ~(input_a[8] & input_a[26]);
  assign popcount36_ssce_core_058 = ~input_a[17];
  assign popcount36_ssce_core_060 = input_a[19] & input_a[9];
  assign popcount36_ssce_core_062 = ~input_a[13];
  assign popcount36_ssce_core_064 = input_a[22] ^ input_a[31];
  assign popcount36_ssce_core_065 = ~input_a[25];
  assign popcount36_ssce_core_066 = ~(input_a[1] | input_a[12]);
  assign popcount36_ssce_core_068_not = ~input_a[7];
  assign popcount36_ssce_core_070 = ~(input_a[23] ^ input_a[25]);
  assign popcount36_ssce_core_071 = ~(input_a[21] & input_a[31]);
  assign popcount36_ssce_core_072_not = ~input_a[25];
  assign popcount36_ssce_core_074 = ~input_a[32];
  assign popcount36_ssce_core_075 = ~(input_a[20] & input_a[32]);
  assign popcount36_ssce_core_076 = ~(input_a[7] | input_a[2]);
  assign popcount36_ssce_core_077 = ~input_a[17];
  assign popcount36_ssce_core_078 = input_a[3] | input_a[18];
  assign popcount36_ssce_core_079 = ~input_a[4];
  assign popcount36_ssce_core_080 = ~(input_a[30] | input_a[17]);
  assign popcount36_ssce_core_081 = ~input_a[0];
  assign popcount36_ssce_core_085 = ~(input_a[2] ^ input_a[8]);
  assign popcount36_ssce_core_087 = input_a[34] ^ input_a[21];
  assign popcount36_ssce_core_088 = ~(input_a[35] ^ input_a[6]);
  assign popcount36_ssce_core_089 = ~input_a[22];
  assign popcount36_ssce_core_090 = ~(input_a[27] ^ input_a[12]);
  assign popcount36_ssce_core_091 = ~input_a[19];
  assign popcount36_ssce_core_092 = ~(input_a[31] | input_a[34]);
  assign popcount36_ssce_core_093 = input_a[7] ^ input_a[24];
  assign popcount36_ssce_core_097 = ~(input_a[33] ^ input_a[30]);
  assign popcount36_ssce_core_098 = ~input_a[3];
  assign popcount36_ssce_core_099 = input_a[0] ^ input_a[17];
  assign popcount36_ssce_core_100 = ~(input_a[26] & input_a[0]);
  assign popcount36_ssce_core_111 = input_a[19] ^ input_a[27];
  assign popcount36_ssce_core_112 = ~(input_a[24] ^ input_a[25]);
  assign popcount36_ssce_core_113 = ~(input_a[26] | input_a[26]);
  assign popcount36_ssce_core_116 = input_a[20] ^ input_a[32];
  assign popcount36_ssce_core_118 = input_a[13] ^ input_a[9];
  assign popcount36_ssce_core_119 = ~input_a[30];
  assign popcount36_ssce_core_122 = ~(input_a[23] ^ input_a[29]);
  assign popcount36_ssce_core_124 = input_a[9] ^ input_a[8];
  assign popcount36_ssce_core_125 = ~(input_a[18] ^ input_a[7]);
  assign popcount36_ssce_core_126 = ~(input_a[33] | input_a[2]);
  assign popcount36_ssce_core_128 = ~(input_a[6] & input_a[19]);
  assign popcount36_ssce_core_129 = input_a[5] & input_a[25];
  assign popcount36_ssce_core_130 = ~(input_a[21] & input_a[19]);
  assign popcount36_ssce_core_131 = ~(input_a[19] ^ input_a[4]);
  assign popcount36_ssce_core_132 = input_a[23] & input_a[5];
  assign popcount36_ssce_core_134 = input_a[11] ^ input_a[7];
  assign popcount36_ssce_core_135 = input_a[27] | input_a[20];
  assign popcount36_ssce_core_138 = ~(input_a[18] | input_a[2]);
  assign popcount36_ssce_core_140 = ~(input_a[2] | input_a[10]);
  assign popcount36_ssce_core_142 = input_a[30] ^ input_a[23];
  assign popcount36_ssce_core_143 = ~input_a[8];
  assign popcount36_ssce_core_144 = input_a[16] | input_a[33];
  assign popcount36_ssce_core_145 = ~(input_a[28] | input_a[29]);
  assign popcount36_ssce_core_146 = ~input_a[7];
  assign popcount36_ssce_core_147 = input_a[25] | input_a[0];
  assign popcount36_ssce_core_148 = ~input_a[5];
  assign popcount36_ssce_core_150 = ~(input_a[22] | input_a[27]);
  assign popcount36_ssce_core_151 = ~(input_a[17] ^ input_a[21]);
  assign popcount36_ssce_core_152 = ~(input_a[7] ^ input_a[28]);
  assign popcount36_ssce_core_154 = input_a[6] ^ input_a[6];
  assign popcount36_ssce_core_155 = ~(input_a[34] ^ input_a[5]);
  assign popcount36_ssce_core_160 = input_a[31] | input_a[13];
  assign popcount36_ssce_core_161 = ~(input_a[32] | input_a[3]);
  assign popcount36_ssce_core_163 = ~(input_a[0] | input_a[20]);
  assign popcount36_ssce_core_164 = ~(input_a[23] ^ input_a[1]);
  assign popcount36_ssce_core_166 = input_a[15] ^ input_a[35];
  assign popcount36_ssce_core_167 = input_a[18] & input_a[4];
  assign popcount36_ssce_core_168 = input_a[15] | input_a[29];
  assign popcount36_ssce_core_169 = input_a[34] | input_a[25];
  assign popcount36_ssce_core_170 = input_a[6] | input_a[29];
  assign popcount36_ssce_core_171 = input_a[7] ^ input_a[34];
  assign popcount36_ssce_core_174 = ~(input_a[24] & input_a[13]);
  assign popcount36_ssce_core_176 = ~input_a[2];
  assign popcount36_ssce_core_179 = ~(input_a[7] | input_a[20]);
  assign popcount36_ssce_core_181 = ~input_a[26];
  assign popcount36_ssce_core_182 = ~(input_a[14] ^ input_a[12]);
  assign popcount36_ssce_core_183_not = ~input_a[14];
  assign popcount36_ssce_core_185 = input_a[1] | input_a[1];
  assign popcount36_ssce_core_186 = input_a[30] ^ input_a[25];
  assign popcount36_ssce_core_187 = ~(input_a[25] | input_a[4]);
  assign popcount36_ssce_core_189 = ~(input_a[6] & input_a[6]);
  assign popcount36_ssce_core_190 = ~input_a[33];
  assign popcount36_ssce_core_191 = ~input_a[6];
  assign popcount36_ssce_core_193 = ~(input_a[6] & input_a[26]);
  assign popcount36_ssce_core_195 = ~(input_a[0] | input_a[7]);
  assign popcount36_ssce_core_197 = ~(input_a[13] ^ input_a[34]);
  assign popcount36_ssce_core_198 = ~(input_a[25] & input_a[7]);
  assign popcount36_ssce_core_199 = ~(input_a[24] | input_a[6]);
  assign popcount36_ssce_core_201 = input_a[35] | input_a[31];
  assign popcount36_ssce_core_202 = ~(input_a[4] | input_a[21]);
  assign popcount36_ssce_core_203 = ~(input_a[11] & input_a[1]);
  assign popcount36_ssce_core_204 = input_a[34] | input_a[5];
  assign popcount36_ssce_core_208 = input_a[17] | input_a[0];
  assign popcount36_ssce_core_209 = ~(input_a[30] ^ input_a[15]);
  assign popcount36_ssce_core_211 = ~(input_a[12] ^ input_a[11]);
  assign popcount36_ssce_core_213 = ~(input_a[35] & input_a[0]);
  assign popcount36_ssce_core_214 = ~(input_a[20] & input_a[14]);
  assign popcount36_ssce_core_215 = ~(input_a[5] & input_a[6]);
  assign popcount36_ssce_core_219 = ~(input_a[10] | input_a[11]);
  assign popcount36_ssce_core_220 = ~(input_a[34] & input_a[12]);
  assign popcount36_ssce_core_222_not = ~input_a[2];
  assign popcount36_ssce_core_225 = ~input_a[34];
  assign popcount36_ssce_core_226 = input_a[10] ^ input_a[9];
  assign popcount36_ssce_core_227 = ~input_a[8];
  assign popcount36_ssce_core_228 = ~(input_a[13] & input_a[16]);
  assign popcount36_ssce_core_229 = input_a[26] ^ input_a[13];
  assign popcount36_ssce_core_230 = ~(input_a[14] | input_a[28]);
  assign popcount36_ssce_core_231 = input_a[12] | input_a[13];
  assign popcount36_ssce_core_232 = input_a[17] ^ input_a[16];
  assign popcount36_ssce_core_233 = ~(input_a[23] | input_a[28]);
  assign popcount36_ssce_core_236 = input_a[31] | input_a[30];
  assign popcount36_ssce_core_237 = ~(input_a[16] & input_a[31]);
  assign popcount36_ssce_core_238 = input_a[0] ^ input_a[5];
  assign popcount36_ssce_core_242 = input_a[35] | input_a[0];
  assign popcount36_ssce_core_243 = ~(input_a[5] & input_a[20]);
  assign popcount36_ssce_core_244 = input_a[10] ^ input_a[23];
  assign popcount36_ssce_core_245 = ~input_a[22];
  assign popcount36_ssce_core_246 = ~(input_a[9] & input_a[34]);
  assign popcount36_ssce_core_247 = input_a[23] ^ input_a[7];
  assign popcount36_ssce_core_248 = ~(input_a[8] | input_a[23]);
  assign popcount36_ssce_core_249 = input_a[7] & input_a[16];
  assign popcount36_ssce_core_250 = ~(input_a[21] & input_a[19]);
  assign popcount36_ssce_core_251_not = ~input_a[14];
  assign popcount36_ssce_core_254 = ~(input_a[20] | input_a[0]);
  assign popcount36_ssce_core_255 = ~(input_a[31] & input_a[35]);
  assign popcount36_ssce_core_256 = ~(input_a[7] ^ input_a[26]);
  assign popcount36_ssce_core_257 = ~(input_a[25] | input_a[28]);
  assign popcount36_ssce_core_258 = ~(input_a[0] ^ input_a[3]);
  assign popcount36_ssce_core_260 = ~(input_a[34] & input_a[33]);
  assign popcount36_ssce_core_261 = ~(input_a[34] | input_a[17]);
  assign popcount36_ssce_core_263 = ~input_a[1];
  assign popcount36_ssce_core_265 = input_a[7] & input_a[22];
  assign popcount36_ssce_core_267 = ~input_a[2];
  assign popcount36_ssce_core_269 = input_a[8] | input_a[20];
  assign popcount36_ssce_core_270 = ~input_a[15];
  assign popcount36_ssce_core_273 = input_a[25] | input_a[7];
  assign popcount36_ssce_core_274 = input_a[10] & input_a[0];

  assign popcount36_ssce_out[0] = 1'b1;
  assign popcount36_ssce_out[1] = 1'b1;
  assign popcount36_ssce_out[2] = input_a[12];
  assign popcount36_ssce_out[3] = 1'b1;
  assign popcount36_ssce_out[4] = input_a[12];
  assign popcount36_ssce_out[5] = 1'b0;
endmodule