// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.2915
// WCE=18.0
// EP=0.932187%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_cmon(input [21:0] input_a, output [4:0] popcount22_cmon_out);
  wire popcount22_cmon_core_025;
  wire popcount22_cmon_core_027;
  wire popcount22_cmon_core_029;
  wire popcount22_cmon_core_030;
  wire popcount22_cmon_core_031;
  wire popcount22_cmon_core_032;
  wire popcount22_cmon_core_033;
  wire popcount22_cmon_core_034;
  wire popcount22_cmon_core_036;
  wire popcount22_cmon_core_037;
  wire popcount22_cmon_core_039;
  wire popcount22_cmon_core_041;
  wire popcount22_cmon_core_042;
  wire popcount22_cmon_core_043;
  wire popcount22_cmon_core_044;
  wire popcount22_cmon_core_045;
  wire popcount22_cmon_core_046;
  wire popcount22_cmon_core_047;
  wire popcount22_cmon_core_050;
  wire popcount22_cmon_core_051;
  wire popcount22_cmon_core_053;
  wire popcount22_cmon_core_055;
  wire popcount22_cmon_core_057;
  wire popcount22_cmon_core_059;
  wire popcount22_cmon_core_060;
  wire popcount22_cmon_core_061;
  wire popcount22_cmon_core_063;
  wire popcount22_cmon_core_064;
  wire popcount22_cmon_core_065;
  wire popcount22_cmon_core_066;
  wire popcount22_cmon_core_067;
  wire popcount22_cmon_core_068;
  wire popcount22_cmon_core_069;
  wire popcount22_cmon_core_072;
  wire popcount22_cmon_core_073;
  wire popcount22_cmon_core_074;
  wire popcount22_cmon_core_077;
  wire popcount22_cmon_core_078;
  wire popcount22_cmon_core_081;
  wire popcount22_cmon_core_082;
  wire popcount22_cmon_core_083;
  wire popcount22_cmon_core_085;
  wire popcount22_cmon_core_086;
  wire popcount22_cmon_core_087;
  wire popcount22_cmon_core_088;
  wire popcount22_cmon_core_089;
  wire popcount22_cmon_core_092;
  wire popcount22_cmon_core_094;
  wire popcount22_cmon_core_098;
  wire popcount22_cmon_core_099;
  wire popcount22_cmon_core_101;
  wire popcount22_cmon_core_102;
  wire popcount22_cmon_core_103;
  wire popcount22_cmon_core_107_not;
  wire popcount22_cmon_core_108;
  wire popcount22_cmon_core_109;
  wire popcount22_cmon_core_110;
  wire popcount22_cmon_core_111;
  wire popcount22_cmon_core_113;
  wire popcount22_cmon_core_114;
  wire popcount22_cmon_core_115;
  wire popcount22_cmon_core_116;
  wire popcount22_cmon_core_118;
  wire popcount22_cmon_core_119;
  wire popcount22_cmon_core_123;
  wire popcount22_cmon_core_124;
  wire popcount22_cmon_core_125;
  wire popcount22_cmon_core_126;
  wire popcount22_cmon_core_127;
  wire popcount22_cmon_core_128;
  wire popcount22_cmon_core_131;
  wire popcount22_cmon_core_132;
  wire popcount22_cmon_core_133;
  wire popcount22_cmon_core_134;
  wire popcount22_cmon_core_139;
  wire popcount22_cmon_core_140;
  wire popcount22_cmon_core_142_not;
  wire popcount22_cmon_core_144;
  wire popcount22_cmon_core_145;
  wire popcount22_cmon_core_147;
  wire popcount22_cmon_core_148;
  wire popcount22_cmon_core_149;
  wire popcount22_cmon_core_150;
  wire popcount22_cmon_core_152;
  wire popcount22_cmon_core_153;
  wire popcount22_cmon_core_154;
  wire popcount22_cmon_core_155;
  wire popcount22_cmon_core_158;
  wire popcount22_cmon_core_159;
  wire popcount22_cmon_core_161;

  assign popcount22_cmon_core_025 = ~(input_a[17] | input_a[21]);
  assign popcount22_cmon_core_027 = ~input_a[5];
  assign popcount22_cmon_core_029 = ~(input_a[16] ^ input_a[5]);
  assign popcount22_cmon_core_030 = ~(input_a[6] & input_a[5]);
  assign popcount22_cmon_core_031 = ~(input_a[20] & input_a[17]);
  assign popcount22_cmon_core_032 = input_a[3] ^ input_a[17];
  assign popcount22_cmon_core_033 = ~(input_a[16] | input_a[13]);
  assign popcount22_cmon_core_034 = ~(input_a[16] ^ input_a[15]);
  assign popcount22_cmon_core_036 = ~(input_a[15] ^ input_a[9]);
  assign popcount22_cmon_core_037 = input_a[9] | input_a[16];
  assign popcount22_cmon_core_039 = ~input_a[11];
  assign popcount22_cmon_core_041 = ~(input_a[20] & input_a[0]);
  assign popcount22_cmon_core_042 = input_a[2] & input_a[14];
  assign popcount22_cmon_core_043 = ~input_a[16];
  assign popcount22_cmon_core_044 = ~(input_a[2] | input_a[6]);
  assign popcount22_cmon_core_045 = input_a[3] ^ input_a[7];
  assign popcount22_cmon_core_046 = ~input_a[2];
  assign popcount22_cmon_core_047 = input_a[6] & input_a[3];
  assign popcount22_cmon_core_050 = ~input_a[9];
  assign popcount22_cmon_core_051 = ~input_a[4];
  assign popcount22_cmon_core_053 = input_a[16] ^ input_a[7];
  assign popcount22_cmon_core_055 = input_a[1] ^ input_a[14];
  assign popcount22_cmon_core_057 = input_a[0] | input_a[8];
  assign popcount22_cmon_core_059 = input_a[15] | input_a[15];
  assign popcount22_cmon_core_060 = input_a[4] & input_a[9];
  assign popcount22_cmon_core_061 = input_a[9] ^ input_a[11];
  assign popcount22_cmon_core_063 = input_a[0] | input_a[10];
  assign popcount22_cmon_core_064 = input_a[1] | input_a[18];
  assign popcount22_cmon_core_065 = ~(input_a[13] ^ input_a[19]);
  assign popcount22_cmon_core_066 = ~(input_a[6] | input_a[18]);
  assign popcount22_cmon_core_067 = ~(input_a[20] & input_a[12]);
  assign popcount22_cmon_core_068 = ~(input_a[12] | input_a[14]);
  assign popcount22_cmon_core_069 = ~input_a[19];
  assign popcount22_cmon_core_072 = ~(input_a[9] ^ input_a[5]);
  assign popcount22_cmon_core_073 = input_a[6] | input_a[18];
  assign popcount22_cmon_core_074 = input_a[14] & input_a[3];
  assign popcount22_cmon_core_077 = input_a[10] ^ input_a[14];
  assign popcount22_cmon_core_078 = ~(input_a[6] | input_a[0]);
  assign popcount22_cmon_core_081 = ~(input_a[8] & input_a[10]);
  assign popcount22_cmon_core_082 = ~(input_a[12] ^ input_a[0]);
  assign popcount22_cmon_core_083 = ~(input_a[11] & input_a[12]);
  assign popcount22_cmon_core_085 = ~input_a[10];
  assign popcount22_cmon_core_086 = ~input_a[8];
  assign popcount22_cmon_core_087 = input_a[6] ^ input_a[21];
  assign popcount22_cmon_core_088 = ~(input_a[12] | input_a[6]);
  assign popcount22_cmon_core_089 = input_a[3] & input_a[8];
  assign popcount22_cmon_core_092 = input_a[21] ^ input_a[20];
  assign popcount22_cmon_core_094 = ~(input_a[2] & input_a[2]);
  assign popcount22_cmon_core_098 = ~input_a[3];
  assign popcount22_cmon_core_099 = input_a[16] ^ input_a[2];
  assign popcount22_cmon_core_101 = ~input_a[10];
  assign popcount22_cmon_core_102 = ~(input_a[2] | input_a[2]);
  assign popcount22_cmon_core_103 = ~input_a[18];
  assign popcount22_cmon_core_107_not = ~input_a[11];
  assign popcount22_cmon_core_108 = input_a[9] | input_a[11];
  assign popcount22_cmon_core_109 = ~(input_a[7] & input_a[17]);
  assign popcount22_cmon_core_110 = ~input_a[5];
  assign popcount22_cmon_core_111 = ~input_a[19];
  assign popcount22_cmon_core_113 = ~input_a[20];
  assign popcount22_cmon_core_114 = ~(input_a[8] | input_a[17]);
  assign popcount22_cmon_core_115 = input_a[10] | input_a[15];
  assign popcount22_cmon_core_116 = input_a[11] & input_a[2];
  assign popcount22_cmon_core_118 = ~(input_a[11] ^ input_a[5]);
  assign popcount22_cmon_core_119 = input_a[3] ^ input_a[9];
  assign popcount22_cmon_core_123 = input_a[11] ^ input_a[15];
  assign popcount22_cmon_core_124 = input_a[19] | input_a[19];
  assign popcount22_cmon_core_125 = ~(input_a[0] | input_a[8]);
  assign popcount22_cmon_core_126 = input_a[10] | input_a[0];
  assign popcount22_cmon_core_127 = ~input_a[14];
  assign popcount22_cmon_core_128 = input_a[16] ^ input_a[19];
  assign popcount22_cmon_core_131 = input_a[5] ^ input_a[12];
  assign popcount22_cmon_core_132 = ~(input_a[6] & input_a[20]);
  assign popcount22_cmon_core_133 = input_a[8] ^ input_a[8];
  assign popcount22_cmon_core_134 = ~input_a[17];
  assign popcount22_cmon_core_139 = input_a[20] & input_a[18];
  assign popcount22_cmon_core_140 = ~(input_a[7] | input_a[4]);
  assign popcount22_cmon_core_142_not = ~input_a[1];
  assign popcount22_cmon_core_144 = ~(input_a[21] | input_a[2]);
  assign popcount22_cmon_core_145 = ~input_a[2];
  assign popcount22_cmon_core_147 = ~(input_a[8] & input_a[9]);
  assign popcount22_cmon_core_148 = ~(input_a[13] & input_a[3]);
  assign popcount22_cmon_core_149 = ~(input_a[20] & input_a[18]);
  assign popcount22_cmon_core_150 = ~input_a[15];
  assign popcount22_cmon_core_152 = input_a[8] ^ input_a[13];
  assign popcount22_cmon_core_153 = ~(input_a[11] | input_a[3]);
  assign popcount22_cmon_core_154 = ~input_a[0];
  assign popcount22_cmon_core_155 = ~input_a[9];
  assign popcount22_cmon_core_158 = ~(input_a[10] & input_a[8]);
  assign popcount22_cmon_core_159 = ~input_a[21];
  assign popcount22_cmon_core_161 = input_a[19] & input_a[10];

  assign popcount22_cmon_out[0] = input_a[3];
  assign popcount22_cmon_out[1] = 1'b1;
  assign popcount22_cmon_out[2] = 1'b1;
  assign popcount22_cmon_out[3] = input_a[4];
  assign popcount22_cmon_out[4] = 1'b0;
endmodule