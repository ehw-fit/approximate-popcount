// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.16618
// WCE=28.0
// EP=0.973036%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_ez8k(input [27:0] input_a, output [4:0] popcount28_ez8k_out);
  wire popcount28_ez8k_core_031;
  wire popcount28_ez8k_core_034;
  wire popcount28_ez8k_core_035;
  wire popcount28_ez8k_core_036;
  wire popcount28_ez8k_core_039;
  wire popcount28_ez8k_core_040;
  wire popcount28_ez8k_core_041;
  wire popcount28_ez8k_core_042;
  wire popcount28_ez8k_core_045;
  wire popcount28_ez8k_core_046;
  wire popcount28_ez8k_core_047;
  wire popcount28_ez8k_core_048;
  wire popcount28_ez8k_core_050;
  wire popcount28_ez8k_core_051;
  wire popcount28_ez8k_core_052;
  wire popcount28_ez8k_core_054;
  wire popcount28_ez8k_core_055;
  wire popcount28_ez8k_core_056;
  wire popcount28_ez8k_core_058;
  wire popcount28_ez8k_core_059;
  wire popcount28_ez8k_core_061;
  wire popcount28_ez8k_core_063;
  wire popcount28_ez8k_core_064;
  wire popcount28_ez8k_core_068;
  wire popcount28_ez8k_core_069;
  wire popcount28_ez8k_core_070;
  wire popcount28_ez8k_core_071;
  wire popcount28_ez8k_core_073;
  wire popcount28_ez8k_core_074;
  wire popcount28_ez8k_core_076;
  wire popcount28_ez8k_core_077;
  wire popcount28_ez8k_core_079;
  wire popcount28_ez8k_core_080;
  wire popcount28_ez8k_core_083;
  wire popcount28_ez8k_core_084;
  wire popcount28_ez8k_core_085;
  wire popcount28_ez8k_core_086;
  wire popcount28_ez8k_core_088;
  wire popcount28_ez8k_core_089;
  wire popcount28_ez8k_core_090;
  wire popcount28_ez8k_core_091;
  wire popcount28_ez8k_core_092;
  wire popcount28_ez8k_core_093;
  wire popcount28_ez8k_core_094;
  wire popcount28_ez8k_core_095;
  wire popcount28_ez8k_core_096;
  wire popcount28_ez8k_core_097;
  wire popcount28_ez8k_core_098;
  wire popcount28_ez8k_core_102;
  wire popcount28_ez8k_core_103;
  wire popcount28_ez8k_core_104;
  wire popcount28_ez8k_core_105;
  wire popcount28_ez8k_core_106;
  wire popcount28_ez8k_core_108;
  wire popcount28_ez8k_core_109;
  wire popcount28_ez8k_core_110;
  wire popcount28_ez8k_core_112;
  wire popcount28_ez8k_core_113;
  wire popcount28_ez8k_core_114;
  wire popcount28_ez8k_core_116;
  wire popcount28_ez8k_core_117;
  wire popcount28_ez8k_core_118;
  wire popcount28_ez8k_core_119;
  wire popcount28_ez8k_core_121;
  wire popcount28_ez8k_core_123;
  wire popcount28_ez8k_core_124;
  wire popcount28_ez8k_core_125;
  wire popcount28_ez8k_core_127;
  wire popcount28_ez8k_core_128;
  wire popcount28_ez8k_core_129;
  wire popcount28_ez8k_core_130;
  wire popcount28_ez8k_core_132;
  wire popcount28_ez8k_core_134;
  wire popcount28_ez8k_core_135;
  wire popcount28_ez8k_core_136;
  wire popcount28_ez8k_core_139;
  wire popcount28_ez8k_core_140;
  wire popcount28_ez8k_core_141;
  wire popcount28_ez8k_core_143;
  wire popcount28_ez8k_core_144;
  wire popcount28_ez8k_core_145;
  wire popcount28_ez8k_core_146;
  wire popcount28_ez8k_core_149;
  wire popcount28_ez8k_core_151;
  wire popcount28_ez8k_core_152;
  wire popcount28_ez8k_core_153;
  wire popcount28_ez8k_core_155;
  wire popcount28_ez8k_core_159;
  wire popcount28_ez8k_core_160;
  wire popcount28_ez8k_core_161;
  wire popcount28_ez8k_core_164;
  wire popcount28_ez8k_core_167;
  wire popcount28_ez8k_core_168;
  wire popcount28_ez8k_core_173_not;
  wire popcount28_ez8k_core_174;
  wire popcount28_ez8k_core_175;
  wire popcount28_ez8k_core_176;
  wire popcount28_ez8k_core_177;
  wire popcount28_ez8k_core_178;
  wire popcount28_ez8k_core_179;
  wire popcount28_ez8k_core_180;
  wire popcount28_ez8k_core_183;
  wire popcount28_ez8k_core_184;
  wire popcount28_ez8k_core_185;
  wire popcount28_ez8k_core_186;
  wire popcount28_ez8k_core_187;
  wire popcount28_ez8k_core_188;
  wire popcount28_ez8k_core_190;
  wire popcount28_ez8k_core_191;
  wire popcount28_ez8k_core_192;
  wire popcount28_ez8k_core_193;
  wire popcount28_ez8k_core_195;
  wire popcount28_ez8k_core_196;
  wire popcount28_ez8k_core_197;
  wire popcount28_ez8k_core_199;
  wire popcount28_ez8k_core_200;

  assign popcount28_ez8k_core_031 = input_a[10] | input_a[22];
  assign popcount28_ez8k_core_034 = input_a[1] & input_a[23];
  assign popcount28_ez8k_core_035 = ~(input_a[20] & input_a[15]);
  assign popcount28_ez8k_core_036 = ~(input_a[23] ^ input_a[9]);
  assign popcount28_ez8k_core_039 = ~(input_a[22] & input_a[12]);
  assign popcount28_ez8k_core_040 = input_a[14] ^ input_a[27];
  assign popcount28_ez8k_core_041 = ~(input_a[19] ^ input_a[9]);
  assign popcount28_ez8k_core_042 = ~(input_a[3] ^ input_a[18]);
  assign popcount28_ez8k_core_045 = ~(input_a[9] | input_a[2]);
  assign popcount28_ez8k_core_046 = input_a[16] ^ input_a[4];
  assign popcount28_ez8k_core_047 = input_a[20] ^ input_a[26];
  assign popcount28_ez8k_core_048 = input_a[9] & input_a[19];
  assign popcount28_ez8k_core_050 = input_a[7] & input_a[4];
  assign popcount28_ez8k_core_051 = ~(input_a[17] | input_a[23]);
  assign popcount28_ez8k_core_052 = ~(input_a[1] ^ input_a[13]);
  assign popcount28_ez8k_core_054 = input_a[19] & input_a[10];
  assign popcount28_ez8k_core_055 = input_a[3] ^ input_a[23];
  assign popcount28_ez8k_core_056 = ~(input_a[26] | input_a[10]);
  assign popcount28_ez8k_core_058 = input_a[20] ^ input_a[22];
  assign popcount28_ez8k_core_059 = ~input_a[21];
  assign popcount28_ez8k_core_061 = ~input_a[21];
  assign popcount28_ez8k_core_063 = input_a[16] & input_a[24];
  assign popcount28_ez8k_core_064 = input_a[6] ^ input_a[16];
  assign popcount28_ez8k_core_068 = ~(input_a[21] | input_a[3]);
  assign popcount28_ez8k_core_069 = ~(input_a[21] ^ input_a[27]);
  assign popcount28_ez8k_core_070 = ~(input_a[25] & input_a[27]);
  assign popcount28_ez8k_core_071 = ~(input_a[4] | input_a[13]);
  assign popcount28_ez8k_core_073 = input_a[18] ^ input_a[11];
  assign popcount28_ez8k_core_074 = ~input_a[9];
  assign popcount28_ez8k_core_076 = input_a[15] & input_a[11];
  assign popcount28_ez8k_core_077 = ~(input_a[23] & input_a[23]);
  assign popcount28_ez8k_core_079 = ~(input_a[25] | input_a[10]);
  assign popcount28_ez8k_core_080 = ~(input_a[23] & input_a[27]);
  assign popcount28_ez8k_core_083 = ~(input_a[2] | input_a[22]);
  assign popcount28_ez8k_core_084 = input_a[7] & input_a[0];
  assign popcount28_ez8k_core_085 = ~(input_a[16] | input_a[0]);
  assign popcount28_ez8k_core_086 = ~input_a[24];
  assign popcount28_ez8k_core_088 = ~input_a[6];
  assign popcount28_ez8k_core_089 = ~(input_a[4] ^ input_a[20]);
  assign popcount28_ez8k_core_090 = input_a[3] & input_a[5];
  assign popcount28_ez8k_core_091 = input_a[9] ^ input_a[8];
  assign popcount28_ez8k_core_092 = ~input_a[3];
  assign popcount28_ez8k_core_093 = ~input_a[15];
  assign popcount28_ez8k_core_094 = input_a[10] | input_a[17];
  assign popcount28_ez8k_core_095 = ~(input_a[22] ^ input_a[26]);
  assign popcount28_ez8k_core_096 = input_a[6] | input_a[2];
  assign popcount28_ez8k_core_097 = ~(input_a[17] & input_a[2]);
  assign popcount28_ez8k_core_098 = ~(input_a[16] & input_a[4]);
  assign popcount28_ez8k_core_102 = ~(input_a[16] ^ input_a[20]);
  assign popcount28_ez8k_core_103 = input_a[5] | input_a[4];
  assign popcount28_ez8k_core_104 = input_a[16] | input_a[17];
  assign popcount28_ez8k_core_105 = input_a[14] ^ input_a[3];
  assign popcount28_ez8k_core_106 = input_a[2] ^ input_a[16];
  assign popcount28_ez8k_core_108 = ~(input_a[1] ^ input_a[19]);
  assign popcount28_ez8k_core_109 = ~(input_a[15] & input_a[21]);
  assign popcount28_ez8k_core_110 = input_a[23] | input_a[27];
  assign popcount28_ez8k_core_112 = ~input_a[24];
  assign popcount28_ez8k_core_113 = ~(input_a[2] | input_a[14]);
  assign popcount28_ez8k_core_114 = input_a[6] ^ input_a[20];
  assign popcount28_ez8k_core_116 = ~(input_a[7] ^ input_a[12]);
  assign popcount28_ez8k_core_117 = input_a[14] | input_a[22];
  assign popcount28_ez8k_core_118 = ~(input_a[27] ^ input_a[15]);
  assign popcount28_ez8k_core_119 = input_a[6] | input_a[21];
  assign popcount28_ez8k_core_121 = ~input_a[27];
  assign popcount28_ez8k_core_123 = input_a[0] | input_a[22];
  assign popcount28_ez8k_core_124 = ~(input_a[23] | input_a[27]);
  assign popcount28_ez8k_core_125 = ~(input_a[18] | input_a[12]);
  assign popcount28_ez8k_core_127 = input_a[18] | input_a[21];
  assign popcount28_ez8k_core_128 = input_a[21] | input_a[13];
  assign popcount28_ez8k_core_129 = ~input_a[24];
  assign popcount28_ez8k_core_130 = input_a[21] ^ input_a[27];
  assign popcount28_ez8k_core_132 = input_a[26] & input_a[1];
  assign popcount28_ez8k_core_134 = input_a[25] ^ input_a[13];
  assign popcount28_ez8k_core_135 = input_a[22] & input_a[9];
  assign popcount28_ez8k_core_136 = ~(input_a[3] ^ input_a[23]);
  assign popcount28_ez8k_core_139 = input_a[4] & input_a[19];
  assign popcount28_ez8k_core_140 = ~(input_a[14] ^ input_a[3]);
  assign popcount28_ez8k_core_141 = ~(input_a[1] ^ input_a[14]);
  assign popcount28_ez8k_core_143 = input_a[21] ^ input_a[2];
  assign popcount28_ez8k_core_144 = input_a[20] ^ input_a[20];
  assign popcount28_ez8k_core_145 = ~(input_a[14] | input_a[14]);
  assign popcount28_ez8k_core_146 = ~(input_a[19] | input_a[22]);
  assign popcount28_ez8k_core_149 = input_a[6] ^ input_a[16];
  assign popcount28_ez8k_core_151 = ~(input_a[0] & input_a[20]);
  assign popcount28_ez8k_core_152 = ~(input_a[6] | input_a[12]);
  assign popcount28_ez8k_core_153 = ~(input_a[19] | input_a[20]);
  assign popcount28_ez8k_core_155 = ~input_a[20];
  assign popcount28_ez8k_core_159 = input_a[5] ^ input_a[1];
  assign popcount28_ez8k_core_160 = ~(input_a[6] | input_a[17]);
  assign popcount28_ez8k_core_161 = input_a[22] | input_a[2];
  assign popcount28_ez8k_core_164 = ~(input_a[27] | input_a[21]);
  assign popcount28_ez8k_core_167 = ~input_a[18];
  assign popcount28_ez8k_core_168 = ~(input_a[10] | input_a[0]);
  assign popcount28_ez8k_core_173_not = ~input_a[16];
  assign popcount28_ez8k_core_174 = ~input_a[12];
  assign popcount28_ez8k_core_175 = ~(input_a[19] & input_a[3]);
  assign popcount28_ez8k_core_176 = input_a[14] ^ input_a[19];
  assign popcount28_ez8k_core_177 = input_a[12] | input_a[25];
  assign popcount28_ez8k_core_178 = ~(input_a[16] & input_a[11]);
  assign popcount28_ez8k_core_179 = ~(input_a[11] | input_a[14]);
  assign popcount28_ez8k_core_180 = input_a[20] & input_a[13];
  assign popcount28_ez8k_core_183 = input_a[12] & input_a[8];
  assign popcount28_ez8k_core_184 = input_a[20] | input_a[14];
  assign popcount28_ez8k_core_185 = input_a[22] & input_a[17];
  assign popcount28_ez8k_core_186 = input_a[5] ^ input_a[19];
  assign popcount28_ez8k_core_187 = ~(input_a[23] & input_a[23]);
  assign popcount28_ez8k_core_188 = input_a[19] ^ input_a[8];
  assign popcount28_ez8k_core_190 = input_a[16] | input_a[12];
  assign popcount28_ez8k_core_191 = ~(input_a[23] & input_a[16]);
  assign popcount28_ez8k_core_192 = input_a[9] | input_a[0];
  assign popcount28_ez8k_core_193 = ~(input_a[2] ^ input_a[5]);
  assign popcount28_ez8k_core_195 = input_a[4] & input_a[14];
  assign popcount28_ez8k_core_196 = ~(input_a[27] ^ input_a[7]);
  assign popcount28_ez8k_core_197 = ~(input_a[20] & input_a[19]);
  assign popcount28_ez8k_core_199 = input_a[23] & input_a[23];
  assign popcount28_ez8k_core_200 = input_a[0] & input_a[9];

  assign popcount28_ez8k_out[0] = 1'b1;
  assign popcount28_ez8k_out[1] = input_a[1];
  assign popcount28_ez8k_out[2] = input_a[26];
  assign popcount28_ez8k_out[3] = input_a[7];
  assign popcount28_ez8k_out[4] = 1'b1;
endmodule