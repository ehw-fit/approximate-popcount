// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.5385
// WCE=13.0
// EP=0.796093%
// Printed PDK parameters:
//  Area=44023844.0
//  Delay=66198628.0
//  Power=2346000.0

module popcount31_x8ez(input [30:0] input_a, output [4:0] popcount31_x8ez_out);
  wire popcount31_x8ez_core_033;
  wire popcount31_x8ez_core_034;
  wire popcount31_x8ez_core_035;
  wire popcount31_x8ez_core_036;
  wire popcount31_x8ez_core_037;
  wire popcount31_x8ez_core_038;
  wire popcount31_x8ez_core_040;
  wire popcount31_x8ez_core_041;
  wire popcount31_x8ez_core_042;
  wire popcount31_x8ez_core_043;
  wire popcount31_x8ez_core_044;
  wire popcount31_x8ez_core_045;
  wire popcount31_x8ez_core_046;
  wire popcount31_x8ez_core_047;
  wire popcount31_x8ez_core_048;
  wire popcount31_x8ez_core_049;
  wire popcount31_x8ez_core_051;
  wire popcount31_x8ez_core_052;
  wire popcount31_x8ez_core_054;
  wire popcount31_x8ez_core_055;
  wire popcount31_x8ez_core_056;
  wire popcount31_x8ez_core_058;
  wire popcount31_x8ez_core_060;
  wire popcount31_x8ez_core_062;
  wire popcount31_x8ez_core_064;
  wire popcount31_x8ez_core_065;
  wire popcount31_x8ez_core_066;
  wire popcount31_x8ez_core_067;
  wire popcount31_x8ez_core_068;
  wire popcount31_x8ez_core_069;
  wire popcount31_x8ez_core_070;
  wire popcount31_x8ez_core_072;
  wire popcount31_x8ez_core_073;
  wire popcount31_x8ez_core_074;
  wire popcount31_x8ez_core_075;
  wire popcount31_x8ez_core_076;
  wire popcount31_x8ez_core_077;
  wire popcount31_x8ez_core_078;
  wire popcount31_x8ez_core_079;
  wire popcount31_x8ez_core_080;
  wire popcount31_x8ez_core_081;
  wire popcount31_x8ez_core_082;
  wire popcount31_x8ez_core_084;
  wire popcount31_x8ez_core_086;
  wire popcount31_x8ez_core_087;
  wire popcount31_x8ez_core_091;
  wire popcount31_x8ez_core_092_not;
  wire popcount31_x8ez_core_093;
  wire popcount31_x8ez_core_095;
  wire popcount31_x8ez_core_096;
  wire popcount31_x8ez_core_097;
  wire popcount31_x8ez_core_098;
  wire popcount31_x8ez_core_100;
  wire popcount31_x8ez_core_102;
  wire popcount31_x8ez_core_103;
  wire popcount31_x8ez_core_105;
  wire popcount31_x8ez_core_107;
  wire popcount31_x8ez_core_108;
  wire popcount31_x8ez_core_110;
  wire popcount31_x8ez_core_111;
  wire popcount31_x8ez_core_112;
  wire popcount31_x8ez_core_113;
  wire popcount31_x8ez_core_114;
  wire popcount31_x8ez_core_116;
  wire popcount31_x8ez_core_118;
  wire popcount31_x8ez_core_119;
  wire popcount31_x8ez_core_120;
  wire popcount31_x8ez_core_122;
  wire popcount31_x8ez_core_125;
  wire popcount31_x8ez_core_126;
  wire popcount31_x8ez_core_127;
  wire popcount31_x8ez_core_129;
  wire popcount31_x8ez_core_130;
  wire popcount31_x8ez_core_131;
  wire popcount31_x8ez_core_133;
  wire popcount31_x8ez_core_136;
  wire popcount31_x8ez_core_137;
  wire popcount31_x8ez_core_138;
  wire popcount31_x8ez_core_139;
  wire popcount31_x8ez_core_140;
  wire popcount31_x8ez_core_141;
  wire popcount31_x8ez_core_142;
  wire popcount31_x8ez_core_144;
  wire popcount31_x8ez_core_145;
  wire popcount31_x8ez_core_147;
  wire popcount31_x8ez_core_148;
  wire popcount31_x8ez_core_149;
  wire popcount31_x8ez_core_150;
  wire popcount31_x8ez_core_152;
  wire popcount31_x8ez_core_154;
  wire popcount31_x8ez_core_156;
  wire popcount31_x8ez_core_157;
  wire popcount31_x8ez_core_158;
  wire popcount31_x8ez_core_159;
  wire popcount31_x8ez_core_160;
  wire popcount31_x8ez_core_161;
  wire popcount31_x8ez_core_165;
  wire popcount31_x8ez_core_166;
  wire popcount31_x8ez_core_167;
  wire popcount31_x8ez_core_169;
  wire popcount31_x8ez_core_170;
  wire popcount31_x8ez_core_171;
  wire popcount31_x8ez_core_172;
  wire popcount31_x8ez_core_173;
  wire popcount31_x8ez_core_174;
  wire popcount31_x8ez_core_175;
  wire popcount31_x8ez_core_177;
  wire popcount31_x8ez_core_179;
  wire popcount31_x8ez_core_182;
  wire popcount31_x8ez_core_183;
  wire popcount31_x8ez_core_184;
  wire popcount31_x8ez_core_186;
  wire popcount31_x8ez_core_188;
  wire popcount31_x8ez_core_189;
  wire popcount31_x8ez_core_190;
  wire popcount31_x8ez_core_191;
  wire popcount31_x8ez_core_192;
  wire popcount31_x8ez_core_194;
  wire popcount31_x8ez_core_195;
  wire popcount31_x8ez_core_196;
  wire popcount31_x8ez_core_197;
  wire popcount31_x8ez_core_198;
  wire popcount31_x8ez_core_199;
  wire popcount31_x8ez_core_200;
  wire popcount31_x8ez_core_201;
  wire popcount31_x8ez_core_203;
  wire popcount31_x8ez_core_205;
  wire popcount31_x8ez_core_206;
  wire popcount31_x8ez_core_207;
  wire popcount31_x8ez_core_208;
  wire popcount31_x8ez_core_209;
  wire popcount31_x8ez_core_210;
  wire popcount31_x8ez_core_211;
  wire popcount31_x8ez_core_212;
  wire popcount31_x8ez_core_213;
  wire popcount31_x8ez_core_214;
  wire popcount31_x8ez_core_219;

  assign popcount31_x8ez_core_033 = input_a[2] | input_a[1];
  assign popcount31_x8ez_core_034 = input_a[2] & input_a[20];
  assign popcount31_x8ez_core_035 = input_a[25] & input_a[16];
  assign popcount31_x8ez_core_036 = input_a[0] & input_a[1];
  assign popcount31_x8ez_core_037 = popcount31_x8ez_core_034 | popcount31_x8ez_core_036;
  assign popcount31_x8ez_core_038 = input_a[4] | input_a[15];
  assign popcount31_x8ez_core_040 = ~(input_a[8] & input_a[30]);
  assign popcount31_x8ez_core_041 = ~input_a[1];
  assign popcount31_x8ez_core_042 = input_a[10] ^ input_a[30];
  assign popcount31_x8ez_core_043 = ~(input_a[6] & input_a[29]);
  assign popcount31_x8ez_core_044 = ~(input_a[11] | input_a[18]);
  assign popcount31_x8ez_core_045 = ~(input_a[23] & input_a[0]);
  assign popcount31_x8ez_core_046 = ~(input_a[26] | input_a[7]);
  assign popcount31_x8ez_core_047 = ~(input_a[8] ^ input_a[24]);
  assign popcount31_x8ez_core_048 = input_a[6] ^ input_a[14];
  assign popcount31_x8ez_core_049 = ~input_a[15];
  assign popcount31_x8ez_core_051 = input_a[7] & input_a[30];
  assign popcount31_x8ez_core_052 = ~popcount31_x8ez_core_037;
  assign popcount31_x8ez_core_054 = popcount31_x8ez_core_052 ^ popcount31_x8ez_core_051;
  assign popcount31_x8ez_core_055 = input_a[7] & input_a[30];
  assign popcount31_x8ez_core_056 = popcount31_x8ez_core_037 | popcount31_x8ez_core_055;
  assign popcount31_x8ez_core_058 = ~input_a[29];
  assign popcount31_x8ez_core_060 = ~(input_a[13] | input_a[29]);
  assign popcount31_x8ez_core_062 = ~(input_a[1] ^ input_a[0]);
  assign popcount31_x8ez_core_064 = ~input_a[4];
  assign popcount31_x8ez_core_065 = input_a[26] & input_a[22];
  assign popcount31_x8ez_core_066 = input_a[4] ^ input_a[11];
  assign popcount31_x8ez_core_067 = input_a[5] & input_a[1];
  assign popcount31_x8ez_core_068 = input_a[4] | popcount31_x8ez_core_065;
  assign popcount31_x8ez_core_069 = input_a[30] ^ input_a[30];
  assign popcount31_x8ez_core_070 = ~popcount31_x8ez_core_068;
  assign popcount31_x8ez_core_072 = input_a[4] | popcount31_x8ez_core_068;
  assign popcount31_x8ez_core_073 = input_a[11] ^ input_a[12];
  assign popcount31_x8ez_core_074 = input_a[11] & input_a[12];
  assign popcount31_x8ez_core_075 = ~(input_a[2] ^ input_a[12]);
  assign popcount31_x8ez_core_076 = input_a[13] & input_a[14];
  assign popcount31_x8ez_core_077 = input_a[29] | input_a[5];
  assign popcount31_x8ez_core_078 = popcount31_x8ez_core_073 & input_a[24];
  assign popcount31_x8ez_core_079 = popcount31_x8ez_core_074 ^ popcount31_x8ez_core_076;
  assign popcount31_x8ez_core_080 = popcount31_x8ez_core_074 & popcount31_x8ez_core_076;
  assign popcount31_x8ez_core_081 = popcount31_x8ez_core_079 | popcount31_x8ez_core_078;
  assign popcount31_x8ez_core_082 = input_a[22] ^ input_a[27];
  assign popcount31_x8ez_core_084 = input_a[8] & input_a[17];
  assign popcount31_x8ez_core_086 = popcount31_x8ez_core_070 ^ popcount31_x8ez_core_081;
  assign popcount31_x8ez_core_087 = popcount31_x8ez_core_070 & popcount31_x8ez_core_081;
  assign popcount31_x8ez_core_091 = popcount31_x8ez_core_072 ^ popcount31_x8ez_core_080;
  assign popcount31_x8ez_core_092_not = ~input_a[21];
  assign popcount31_x8ez_core_093 = popcount31_x8ez_core_091 | popcount31_x8ez_core_087;
  assign popcount31_x8ez_core_095 = input_a[28] & input_a[1];
  assign popcount31_x8ez_core_096 = ~input_a[15];
  assign popcount31_x8ez_core_097 = ~(input_a[26] | input_a[0]);
  assign popcount31_x8ez_core_098 = popcount31_x8ez_core_054 ^ popcount31_x8ez_core_086;
  assign popcount31_x8ez_core_100 = ~popcount31_x8ez_core_098;
  assign popcount31_x8ez_core_102 = popcount31_x8ez_core_054 | popcount31_x8ez_core_098;
  assign popcount31_x8ez_core_103 = popcount31_x8ez_core_056 ^ popcount31_x8ez_core_093;
  assign popcount31_x8ez_core_105 = popcount31_x8ez_core_103 ^ popcount31_x8ez_core_102;
  assign popcount31_x8ez_core_107 = popcount31_x8ez_core_056 | popcount31_x8ez_core_103;
  assign popcount31_x8ez_core_108 = ~(input_a[12] ^ input_a[6]);
  assign popcount31_x8ez_core_110 = input_a[4] | popcount31_x8ez_core_107;
  assign popcount31_x8ez_core_111 = input_a[1] & input_a[27];
  assign popcount31_x8ez_core_112 = input_a[24] ^ input_a[0];
  assign popcount31_x8ez_core_113 = input_a[12] | input_a[3];
  assign popcount31_x8ez_core_114 = input_a[9] & input_a[25];
  assign popcount31_x8ez_core_116 = input_a[17] & input_a[15];
  assign popcount31_x8ez_core_118 = ~input_a[22];
  assign popcount31_x8ez_core_119 = popcount31_x8ez_core_114 ^ popcount31_x8ez_core_116;
  assign popcount31_x8ez_core_120 = popcount31_x8ez_core_114 & popcount31_x8ez_core_116;
  assign popcount31_x8ez_core_122 = input_a[30] ^ input_a[3];
  assign popcount31_x8ez_core_125 = input_a[19] & input_a[28];
  assign popcount31_x8ez_core_126 = ~input_a[13];
  assign popcount31_x8ez_core_127 = input_a[21] & input_a[5];
  assign popcount31_x8ez_core_129 = input_a[21] & input_a[0];
  assign popcount31_x8ez_core_130 = popcount31_x8ez_core_125 ^ popcount31_x8ez_core_127;
  assign popcount31_x8ez_core_131 = popcount31_x8ez_core_125 & popcount31_x8ez_core_127;
  assign popcount31_x8ez_core_133 = input_a[1] ^ input_a[13];
  assign popcount31_x8ez_core_136 = input_a[3] & input_a[16];
  assign popcount31_x8ez_core_137 = popcount31_x8ez_core_119 ^ popcount31_x8ez_core_130;
  assign popcount31_x8ez_core_138 = popcount31_x8ez_core_119 & popcount31_x8ez_core_130;
  assign popcount31_x8ez_core_139 = popcount31_x8ez_core_137 ^ popcount31_x8ez_core_136;
  assign popcount31_x8ez_core_140 = popcount31_x8ez_core_137 & popcount31_x8ez_core_136;
  assign popcount31_x8ez_core_141 = popcount31_x8ez_core_138 | popcount31_x8ez_core_140;
  assign popcount31_x8ez_core_142 = popcount31_x8ez_core_120 | popcount31_x8ez_core_131;
  assign popcount31_x8ez_core_144 = popcount31_x8ez_core_142 ^ popcount31_x8ez_core_141;
  assign popcount31_x8ez_core_145 = popcount31_x8ez_core_142 & popcount31_x8ez_core_141;
  assign popcount31_x8ez_core_147 = ~(input_a[21] & input_a[29]);
  assign popcount31_x8ez_core_148 = input_a[23] & input_a[18];
  assign popcount31_x8ez_core_149 = input_a[18] ^ input_a[24];
  assign popcount31_x8ez_core_150 = ~input_a[25];
  assign popcount31_x8ez_core_152 = input_a[0] & input_a[13];
  assign popcount31_x8ez_core_154 = input_a[15] | input_a[14];
  assign popcount31_x8ez_core_156 = ~input_a[29];
  assign popcount31_x8ez_core_157 = ~input_a[8];
  assign popcount31_x8ez_core_158 = input_a[4] & input_a[25];
  assign popcount31_x8ez_core_159 = input_a[15] & input_a[23];
  assign popcount31_x8ez_core_160 = ~(input_a[28] | input_a[6]);
  assign popcount31_x8ez_core_161 = ~input_a[19];
  assign popcount31_x8ez_core_165 = input_a[10] ^ input_a[9];
  assign popcount31_x8ez_core_166 = input_a[27] | input_a[10];
  assign popcount31_x8ez_core_167 = input_a[19] & input_a[16];
  assign popcount31_x8ez_core_169 = ~(input_a[1] ^ input_a[4]);
  assign popcount31_x8ez_core_170 = input_a[6] & input_a[29];
  assign popcount31_x8ez_core_171 = popcount31_x8ez_core_148 ^ popcount31_x8ez_core_166;
  assign popcount31_x8ez_core_172 = popcount31_x8ez_core_148 & popcount31_x8ez_core_166;
  assign popcount31_x8ez_core_173 = popcount31_x8ez_core_171 ^ popcount31_x8ez_core_170;
  assign popcount31_x8ez_core_174 = popcount31_x8ez_core_171 & popcount31_x8ez_core_170;
  assign popcount31_x8ez_core_175 = popcount31_x8ez_core_172 | popcount31_x8ez_core_174;
  assign popcount31_x8ez_core_177 = ~(input_a[15] ^ input_a[2]);
  assign popcount31_x8ez_core_179 = input_a[11] | input_a[25];
  assign popcount31_x8ez_core_182 = ~input_a[10];
  assign popcount31_x8ez_core_183 = popcount31_x8ez_core_139 ^ popcount31_x8ez_core_173;
  assign popcount31_x8ez_core_184 = popcount31_x8ez_core_139 & popcount31_x8ez_core_173;
  assign popcount31_x8ez_core_186 = ~input_a[9];
  assign popcount31_x8ez_core_188 = popcount31_x8ez_core_144 ^ popcount31_x8ez_core_175;
  assign popcount31_x8ez_core_189 = popcount31_x8ez_core_144 & popcount31_x8ez_core_175;
  assign popcount31_x8ez_core_190 = popcount31_x8ez_core_188 ^ popcount31_x8ez_core_184;
  assign popcount31_x8ez_core_191 = popcount31_x8ez_core_188 & popcount31_x8ez_core_184;
  assign popcount31_x8ez_core_192 = popcount31_x8ez_core_189 | popcount31_x8ez_core_191;
  assign popcount31_x8ez_core_194 = input_a[23] ^ input_a[0];
  assign popcount31_x8ez_core_195 = popcount31_x8ez_core_145 | popcount31_x8ez_core_192;
  assign popcount31_x8ez_core_196 = input_a[17] | input_a[3];
  assign popcount31_x8ez_core_197 = ~(input_a[20] | input_a[3]);
  assign popcount31_x8ez_core_198 = input_a[21] & input_a[26];
  assign popcount31_x8ez_core_199 = ~(input_a[1] ^ input_a[26]);
  assign popcount31_x8ez_core_200 = popcount31_x8ez_core_100 ^ popcount31_x8ez_core_183;
  assign popcount31_x8ez_core_201 = popcount31_x8ez_core_100 & popcount31_x8ez_core_183;
  assign popcount31_x8ez_core_203 = input_a[16] & input_a[27];
  assign popcount31_x8ez_core_205 = popcount31_x8ez_core_105 ^ popcount31_x8ez_core_190;
  assign popcount31_x8ez_core_206 = popcount31_x8ez_core_105 & popcount31_x8ez_core_190;
  assign popcount31_x8ez_core_207 = popcount31_x8ez_core_205 ^ popcount31_x8ez_core_201;
  assign popcount31_x8ez_core_208 = popcount31_x8ez_core_205 & popcount31_x8ez_core_201;
  assign popcount31_x8ez_core_209 = popcount31_x8ez_core_206 | popcount31_x8ez_core_208;
  assign popcount31_x8ez_core_210 = popcount31_x8ez_core_110 ^ popcount31_x8ez_core_195;
  assign popcount31_x8ez_core_211 = popcount31_x8ez_core_110 & popcount31_x8ez_core_195;
  assign popcount31_x8ez_core_212 = popcount31_x8ez_core_210 ^ popcount31_x8ez_core_209;
  assign popcount31_x8ez_core_213 = popcount31_x8ez_core_210 & popcount31_x8ez_core_209;
  assign popcount31_x8ez_core_214 = popcount31_x8ez_core_211 | popcount31_x8ez_core_213;
  assign popcount31_x8ez_core_219 = ~input_a[0];

  assign popcount31_x8ez_out[0] = input_a[8];
  assign popcount31_x8ez_out[1] = popcount31_x8ez_core_200;
  assign popcount31_x8ez_out[2] = popcount31_x8ez_core_207;
  assign popcount31_x8ez_out[3] = popcount31_x8ez_core_212;
  assign popcount31_x8ez_out[4] = popcount31_x8ez_core_214;
endmodule