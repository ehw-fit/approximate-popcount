// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.76724
// WCE=17.0
// EP=0.887622%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount28_iswk(input [27:0] input_a, output [4:0] popcount28_iswk_out);
  wire popcount28_iswk_core_030;
  wire popcount28_iswk_core_031;
  wire popcount28_iswk_core_032;
  wire popcount28_iswk_core_034;
  wire popcount28_iswk_core_036;
  wire popcount28_iswk_core_038;
  wire popcount28_iswk_core_039;
  wire popcount28_iswk_core_040;
  wire popcount28_iswk_core_041;
  wire popcount28_iswk_core_042;
  wire popcount28_iswk_core_043;
  wire popcount28_iswk_core_044;
  wire popcount28_iswk_core_045;
  wire popcount28_iswk_core_046;
  wire popcount28_iswk_core_047;
  wire popcount28_iswk_core_048;
  wire popcount28_iswk_core_049;
  wire popcount28_iswk_core_053;
  wire popcount28_iswk_core_057;
  wire popcount28_iswk_core_059;
  wire popcount28_iswk_core_063;
  wire popcount28_iswk_core_064;
  wire popcount28_iswk_core_065;
  wire popcount28_iswk_core_066;
  wire popcount28_iswk_core_067;
  wire popcount28_iswk_core_068;
  wire popcount28_iswk_core_069;
  wire popcount28_iswk_core_072;
  wire popcount28_iswk_core_074;
  wire popcount28_iswk_core_075;
  wire popcount28_iswk_core_076;
  wire popcount28_iswk_core_077;
  wire popcount28_iswk_core_078;
  wire popcount28_iswk_core_079;
  wire popcount28_iswk_core_080;
  wire popcount28_iswk_core_081;
  wire popcount28_iswk_core_082;
  wire popcount28_iswk_core_084;
  wire popcount28_iswk_core_086;
  wire popcount28_iswk_core_087;
  wire popcount28_iswk_core_088;
  wire popcount28_iswk_core_089;
  wire popcount28_iswk_core_091;
  wire popcount28_iswk_core_092;
  wire popcount28_iswk_core_093;
  wire popcount28_iswk_core_094;
  wire popcount28_iswk_core_095;
  wire popcount28_iswk_core_096;
  wire popcount28_iswk_core_097;
  wire popcount28_iswk_core_098;
  wire popcount28_iswk_core_099;
  wire popcount28_iswk_core_100;
  wire popcount28_iswk_core_101;
  wire popcount28_iswk_core_103;
  wire popcount28_iswk_core_107;
  wire popcount28_iswk_core_108;
  wire popcount28_iswk_core_109;
  wire popcount28_iswk_core_110_not;
  wire popcount28_iswk_core_114;
  wire popcount28_iswk_core_115;
  wire popcount28_iswk_core_116_not;
  wire popcount28_iswk_core_118;
  wire popcount28_iswk_core_119;
  wire popcount28_iswk_core_122;
  wire popcount28_iswk_core_123;
  wire popcount28_iswk_core_125;
  wire popcount28_iswk_core_126;
  wire popcount28_iswk_core_127;
  wire popcount28_iswk_core_128;
  wire popcount28_iswk_core_129;
  wire popcount28_iswk_core_130;
  wire popcount28_iswk_core_133;
  wire popcount28_iswk_core_134;
  wire popcount28_iswk_core_137;
  wire popcount28_iswk_core_139;
  wire popcount28_iswk_core_140;
  wire popcount28_iswk_core_142;
  wire popcount28_iswk_core_143;
  wire popcount28_iswk_core_146;
  wire popcount28_iswk_core_149;
  wire popcount28_iswk_core_150;
  wire popcount28_iswk_core_152;
  wire popcount28_iswk_core_153;
  wire popcount28_iswk_core_154;
  wire popcount28_iswk_core_155;
  wire popcount28_iswk_core_156;
  wire popcount28_iswk_core_157;
  wire popcount28_iswk_core_158;
  wire popcount28_iswk_core_160;
  wire popcount28_iswk_core_161;
  wire popcount28_iswk_core_163;
  wire popcount28_iswk_core_164;
  wire popcount28_iswk_core_167_not;
  wire popcount28_iswk_core_168;
  wire popcount28_iswk_core_169;
  wire popcount28_iswk_core_170;
  wire popcount28_iswk_core_171;
  wire popcount28_iswk_core_172;
  wire popcount28_iswk_core_173;
  wire popcount28_iswk_core_174;
  wire popcount28_iswk_core_176;
  wire popcount28_iswk_core_177;
  wire popcount28_iswk_core_179;
  wire popcount28_iswk_core_180_not;
  wire popcount28_iswk_core_181;
  wire popcount28_iswk_core_183;
  wire popcount28_iswk_core_184;
  wire popcount28_iswk_core_185_not;
  wire popcount28_iswk_core_189;
  wire popcount28_iswk_core_190;
  wire popcount28_iswk_core_192;
  wire popcount28_iswk_core_194;
  wire popcount28_iswk_core_195_not;
  wire popcount28_iswk_core_197;
  wire popcount28_iswk_core_198;
  wire popcount28_iswk_core_200;
  wire popcount28_iswk_core_201;

  assign popcount28_iswk_core_030 = ~input_a[24];
  assign popcount28_iswk_core_031 = ~(input_a[5] & input_a[23]);
  assign popcount28_iswk_core_032 = ~(input_a[26] ^ input_a[2]);
  assign popcount28_iswk_core_034 = ~(input_a[14] ^ input_a[20]);
  assign popcount28_iswk_core_036 = ~(input_a[24] & input_a[0]);
  assign popcount28_iswk_core_038 = ~(input_a[26] ^ input_a[18]);
  assign popcount28_iswk_core_039 = ~(input_a[16] & input_a[2]);
  assign popcount28_iswk_core_040 = input_a[1] ^ input_a[10];
  assign popcount28_iswk_core_041 = ~(input_a[19] & input_a[4]);
  assign popcount28_iswk_core_042 = ~(input_a[25] & input_a[7]);
  assign popcount28_iswk_core_043 = ~(input_a[14] | input_a[25]);
  assign popcount28_iswk_core_044 = input_a[24] | input_a[0];
  assign popcount28_iswk_core_045 = ~(input_a[13] | input_a[26]);
  assign popcount28_iswk_core_046 = ~(input_a[15] ^ input_a[8]);
  assign popcount28_iswk_core_047 = ~(input_a[13] & input_a[17]);
  assign popcount28_iswk_core_048 = ~(input_a[1] | input_a[4]);
  assign popcount28_iswk_core_049 = ~(input_a[20] ^ input_a[3]);
  assign popcount28_iswk_core_053 = ~input_a[22];
  assign popcount28_iswk_core_057 = input_a[1] & input_a[2];
  assign popcount28_iswk_core_059 = input_a[11] | input_a[26];
  assign popcount28_iswk_core_063 = input_a[27] ^ input_a[23];
  assign popcount28_iswk_core_064 = ~input_a[5];
  assign popcount28_iswk_core_065 = input_a[27] ^ input_a[9];
  assign popcount28_iswk_core_066 = input_a[10] & input_a[19];
  assign popcount28_iswk_core_067 = ~(input_a[20] ^ input_a[14]);
  assign popcount28_iswk_core_068 = input_a[19] | input_a[1];
  assign popcount28_iswk_core_069 = input_a[22] ^ input_a[21];
  assign popcount28_iswk_core_072 = ~input_a[24];
  assign popcount28_iswk_core_074 = ~(input_a[0] & input_a[26]);
  assign popcount28_iswk_core_075 = ~input_a[2];
  assign popcount28_iswk_core_076 = input_a[14] | input_a[22];
  assign popcount28_iswk_core_077 = ~input_a[23];
  assign popcount28_iswk_core_078 = ~input_a[21];
  assign popcount28_iswk_core_079 = input_a[12] & input_a[25];
  assign popcount28_iswk_core_080 = ~(input_a[1] ^ input_a[7]);
  assign popcount28_iswk_core_081 = input_a[27] ^ input_a[14];
  assign popcount28_iswk_core_082 = ~input_a[20];
  assign popcount28_iswk_core_084 = ~input_a[17];
  assign popcount28_iswk_core_086 = ~(input_a[15] & input_a[19]);
  assign popcount28_iswk_core_087 = ~(input_a[20] ^ input_a[19]);
  assign popcount28_iswk_core_088 = ~(input_a[18] ^ input_a[21]);
  assign popcount28_iswk_core_089 = ~(input_a[10] | input_a[0]);
  assign popcount28_iswk_core_091 = ~input_a[19];
  assign popcount28_iswk_core_092 = ~(input_a[7] | input_a[6]);
  assign popcount28_iswk_core_093 = input_a[24] | input_a[0];
  assign popcount28_iswk_core_094 = ~input_a[12];
  assign popcount28_iswk_core_095 = input_a[22] & input_a[21];
  assign popcount28_iswk_core_096 = input_a[23] & input_a[14];
  assign popcount28_iswk_core_097 = ~(input_a[26] | input_a[16]);
  assign popcount28_iswk_core_098 = ~(input_a[22] | input_a[10]);
  assign popcount28_iswk_core_099 = input_a[3] ^ input_a[15];
  assign popcount28_iswk_core_100 = input_a[3] ^ input_a[4];
  assign popcount28_iswk_core_101 = input_a[7] & input_a[11];
  assign popcount28_iswk_core_103 = ~input_a[19];
  assign popcount28_iswk_core_107 = ~input_a[18];
  assign popcount28_iswk_core_108 = ~input_a[25];
  assign popcount28_iswk_core_109 = input_a[23] ^ input_a[12];
  assign popcount28_iswk_core_110_not = ~input_a[20];
  assign popcount28_iswk_core_114 = ~(input_a[7] & input_a[0]);
  assign popcount28_iswk_core_115 = input_a[18] & input_a[16];
  assign popcount28_iswk_core_116_not = ~input_a[5];
  assign popcount28_iswk_core_118 = input_a[6] & input_a[0];
  assign popcount28_iswk_core_119 = ~(input_a[14] & input_a[15]);
  assign popcount28_iswk_core_122 = ~(input_a[24] | input_a[5]);
  assign popcount28_iswk_core_123 = ~(input_a[22] ^ input_a[15]);
  assign popcount28_iswk_core_125 = ~(input_a[27] | input_a[11]);
  assign popcount28_iswk_core_126 = input_a[0] & input_a[10];
  assign popcount28_iswk_core_127 = ~(input_a[23] | input_a[14]);
  assign popcount28_iswk_core_128 = ~input_a[5];
  assign popcount28_iswk_core_129 = ~(input_a[23] & input_a[9]);
  assign popcount28_iswk_core_130 = input_a[25] | input_a[10];
  assign popcount28_iswk_core_133 = ~(input_a[9] ^ input_a[10]);
  assign popcount28_iswk_core_134 = input_a[19] & input_a[3];
  assign popcount28_iswk_core_137 = ~input_a[16];
  assign popcount28_iswk_core_139 = input_a[27] & input_a[20];
  assign popcount28_iswk_core_140 = ~(input_a[19] ^ input_a[26]);
  assign popcount28_iswk_core_142 = ~input_a[7];
  assign popcount28_iswk_core_143 = input_a[20] ^ input_a[13];
  assign popcount28_iswk_core_146 = ~(input_a[0] ^ input_a[12]);
  assign popcount28_iswk_core_149 = ~(input_a[4] | input_a[2]);
  assign popcount28_iswk_core_150 = ~input_a[19];
  assign popcount28_iswk_core_152 = ~(input_a[5] | input_a[17]);
  assign popcount28_iswk_core_153 = input_a[3] | input_a[9];
  assign popcount28_iswk_core_154 = ~(input_a[22] ^ input_a[1]);
  assign popcount28_iswk_core_155 = input_a[14] & input_a[0];
  assign popcount28_iswk_core_156 = input_a[3] ^ input_a[22];
  assign popcount28_iswk_core_157 = input_a[11] | input_a[9];
  assign popcount28_iswk_core_158 = ~input_a[21];
  assign popcount28_iswk_core_160 = ~input_a[15];
  assign popcount28_iswk_core_161 = input_a[3] & input_a[17];
  assign popcount28_iswk_core_163 = ~input_a[1];
  assign popcount28_iswk_core_164 = input_a[26] & input_a[18];
  assign popcount28_iswk_core_167_not = ~input_a[17];
  assign popcount28_iswk_core_168 = ~(input_a[9] | input_a[17]);
  assign popcount28_iswk_core_169 = input_a[4] | input_a[5];
  assign popcount28_iswk_core_170 = input_a[20] | input_a[7];
  assign popcount28_iswk_core_171 = ~(input_a[16] | input_a[7]);
  assign popcount28_iswk_core_172 = ~(input_a[19] | input_a[3]);
  assign popcount28_iswk_core_173 = ~(input_a[9] | input_a[22]);
  assign popcount28_iswk_core_174 = input_a[21] | input_a[20];
  assign popcount28_iswk_core_176 = ~(input_a[17] & input_a[8]);
  assign popcount28_iswk_core_177 = ~(input_a[23] | input_a[2]);
  assign popcount28_iswk_core_179 = ~(input_a[11] & input_a[14]);
  assign popcount28_iswk_core_180_not = ~input_a[11];
  assign popcount28_iswk_core_181 = ~(input_a[24] & input_a[7]);
  assign popcount28_iswk_core_183 = ~input_a[21];
  assign popcount28_iswk_core_184 = input_a[14] | input_a[9];
  assign popcount28_iswk_core_185_not = ~input_a[6];
  assign popcount28_iswk_core_189 = ~(input_a[12] ^ input_a[23]);
  assign popcount28_iswk_core_190 = ~(input_a[12] | input_a[9]);
  assign popcount28_iswk_core_192 = ~(input_a[10] & input_a[17]);
  assign popcount28_iswk_core_194 = ~input_a[18];
  assign popcount28_iswk_core_195_not = ~input_a[10];
  assign popcount28_iswk_core_197 = input_a[2] ^ input_a[13];
  assign popcount28_iswk_core_198 = ~(input_a[9] ^ input_a[21]);
  assign popcount28_iswk_core_200 = ~(input_a[10] | input_a[13]);
  assign popcount28_iswk_core_201 = input_a[19] ^ input_a[18];

  assign popcount28_iswk_out[0] = input_a[10];
  assign popcount28_iswk_out[1] = input_a[10];
  assign popcount28_iswk_out[2] = popcount28_iswk_core_194;
  assign popcount28_iswk_out[3] = popcount28_iswk_core_194;
  assign popcount28_iswk_out[4] = input_a[18];
endmodule