// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.25652
// WCE=13.0
// EP=0.863617%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_yqcn(input [24:0] input_a, output [4:0] popcount25_yqcn_out);
  wire popcount25_yqcn_core_030;
  wire popcount25_yqcn_core_032;
  wire popcount25_yqcn_core_033;
  wire popcount25_yqcn_core_034;
  wire popcount25_yqcn_core_035;
  wire popcount25_yqcn_core_036;
  wire popcount25_yqcn_core_037;
  wire popcount25_yqcn_core_039;
  wire popcount25_yqcn_core_041;
  wire popcount25_yqcn_core_044;
  wire popcount25_yqcn_core_046;
  wire popcount25_yqcn_core_049;
  wire popcount25_yqcn_core_050;
  wire popcount25_yqcn_core_052;
  wire popcount25_yqcn_core_053;
  wire popcount25_yqcn_core_054;
  wire popcount25_yqcn_core_055;
  wire popcount25_yqcn_core_056;
  wire popcount25_yqcn_core_058;
  wire popcount25_yqcn_core_059;
  wire popcount25_yqcn_core_062;
  wire popcount25_yqcn_core_064_not;
  wire popcount25_yqcn_core_066;
  wire popcount25_yqcn_core_068;
  wire popcount25_yqcn_core_069;
  wire popcount25_yqcn_core_070;
  wire popcount25_yqcn_core_072;
  wire popcount25_yqcn_core_073;
  wire popcount25_yqcn_core_074;
  wire popcount25_yqcn_core_075;
  wire popcount25_yqcn_core_076;
  wire popcount25_yqcn_core_077;
  wire popcount25_yqcn_core_079;
  wire popcount25_yqcn_core_081_not;
  wire popcount25_yqcn_core_083;
  wire popcount25_yqcn_core_084;
  wire popcount25_yqcn_core_086;
  wire popcount25_yqcn_core_088;
  wire popcount25_yqcn_core_089_not;
  wire popcount25_yqcn_core_090;
  wire popcount25_yqcn_core_091;
  wire popcount25_yqcn_core_092;
  wire popcount25_yqcn_core_093;
  wire popcount25_yqcn_core_096;
  wire popcount25_yqcn_core_097;
  wire popcount25_yqcn_core_102;
  wire popcount25_yqcn_core_103;
  wire popcount25_yqcn_core_104;
  wire popcount25_yqcn_core_105;
  wire popcount25_yqcn_core_107;
  wire popcount25_yqcn_core_109;
  wire popcount25_yqcn_core_110;
  wire popcount25_yqcn_core_111;
  wire popcount25_yqcn_core_113;
  wire popcount25_yqcn_core_114;
  wire popcount25_yqcn_core_115;
  wire popcount25_yqcn_core_117;
  wire popcount25_yqcn_core_118;
  wire popcount25_yqcn_core_121;
  wire popcount25_yqcn_core_123;
  wire popcount25_yqcn_core_124;
  wire popcount25_yqcn_core_125;
  wire popcount25_yqcn_core_126;
  wire popcount25_yqcn_core_129;
  wire popcount25_yqcn_core_131;
  wire popcount25_yqcn_core_133;
  wire popcount25_yqcn_core_134;
  wire popcount25_yqcn_core_135;
  wire popcount25_yqcn_core_138;
  wire popcount25_yqcn_core_140;
  wire popcount25_yqcn_core_141_not;
  wire popcount25_yqcn_core_142;
  wire popcount25_yqcn_core_143;
  wire popcount25_yqcn_core_144;
  wire popcount25_yqcn_core_146;
  wire popcount25_yqcn_core_147;
  wire popcount25_yqcn_core_148;
  wire popcount25_yqcn_core_149;
  wire popcount25_yqcn_core_150;
  wire popcount25_yqcn_core_152;
  wire popcount25_yqcn_core_155;
  wire popcount25_yqcn_core_156;
  wire popcount25_yqcn_core_157;
  wire popcount25_yqcn_core_159;
  wire popcount25_yqcn_core_160;
  wire popcount25_yqcn_core_163;
  wire popcount25_yqcn_core_165;
  wire popcount25_yqcn_core_167;
  wire popcount25_yqcn_core_169;
  wire popcount25_yqcn_core_171;
  wire popcount25_yqcn_core_173;
  wire popcount25_yqcn_core_175;
  wire popcount25_yqcn_core_178;
  wire popcount25_yqcn_core_180;
  wire popcount25_yqcn_core_181;
  wire popcount25_yqcn_core_182;

  assign popcount25_yqcn_core_030 = ~(input_a[9] & input_a[1]);
  assign popcount25_yqcn_core_032 = input_a[2] ^ input_a[1];
  assign popcount25_yqcn_core_033 = input_a[20] ^ input_a[6];
  assign popcount25_yqcn_core_034 = input_a[2] & input_a[15];
  assign popcount25_yqcn_core_035 = input_a[13] & input_a[11];
  assign popcount25_yqcn_core_036 = ~input_a[12];
  assign popcount25_yqcn_core_037 = input_a[18] & input_a[12];
  assign popcount25_yqcn_core_039 = ~(input_a[14] | input_a[23]);
  assign popcount25_yqcn_core_041 = input_a[16] ^ input_a[13];
  assign popcount25_yqcn_core_044 = input_a[10] | input_a[18];
  assign popcount25_yqcn_core_046 = input_a[5] | input_a[4];
  assign popcount25_yqcn_core_049 = ~input_a[16];
  assign popcount25_yqcn_core_050 = ~(input_a[12] ^ input_a[3]);
  assign popcount25_yqcn_core_052 = ~(input_a[20] & input_a[15]);
  assign popcount25_yqcn_core_053 = input_a[16] | input_a[19];
  assign popcount25_yqcn_core_054 = ~(input_a[1] | input_a[13]);
  assign popcount25_yqcn_core_055 = ~input_a[5];
  assign popcount25_yqcn_core_056 = ~(input_a[17] | input_a[3]);
  assign popcount25_yqcn_core_058 = input_a[14] ^ input_a[15];
  assign popcount25_yqcn_core_059 = ~(input_a[16] ^ input_a[7]);
  assign popcount25_yqcn_core_062 = ~input_a[3];
  assign popcount25_yqcn_core_064_not = ~input_a[0];
  assign popcount25_yqcn_core_066 = input_a[11] | input_a[11];
  assign popcount25_yqcn_core_068 = input_a[1] | input_a[7];
  assign popcount25_yqcn_core_069 = input_a[17] ^ input_a[18];
  assign popcount25_yqcn_core_070 = ~(input_a[11] | input_a[11]);
  assign popcount25_yqcn_core_072 = ~(input_a[24] & input_a[22]);
  assign popcount25_yqcn_core_073 = input_a[5] & input_a[1];
  assign popcount25_yqcn_core_074 = input_a[2] | input_a[13];
  assign popcount25_yqcn_core_075 = input_a[20] | input_a[1];
  assign popcount25_yqcn_core_076 = ~(input_a[1] ^ input_a[6]);
  assign popcount25_yqcn_core_077 = ~input_a[12];
  assign popcount25_yqcn_core_079 = input_a[16] ^ input_a[9];
  assign popcount25_yqcn_core_081_not = ~input_a[1];
  assign popcount25_yqcn_core_083 = input_a[13] ^ input_a[16];
  assign popcount25_yqcn_core_084 = ~(input_a[6] | input_a[16]);
  assign popcount25_yqcn_core_086 = input_a[17] & input_a[8];
  assign popcount25_yqcn_core_088 = ~input_a[8];
  assign popcount25_yqcn_core_089_not = ~input_a[13];
  assign popcount25_yqcn_core_090 = ~(input_a[8] | input_a[22]);
  assign popcount25_yqcn_core_091 = ~(input_a[4] & input_a[15]);
  assign popcount25_yqcn_core_092 = input_a[16] ^ input_a[8];
  assign popcount25_yqcn_core_093 = input_a[7] & input_a[19];
  assign popcount25_yqcn_core_096 = ~(input_a[24] & input_a[7]);
  assign popcount25_yqcn_core_097 = input_a[13] | input_a[21];
  assign popcount25_yqcn_core_102 = input_a[10] ^ input_a[14];
  assign popcount25_yqcn_core_103 = ~(input_a[6] ^ input_a[5]);
  assign popcount25_yqcn_core_104 = input_a[6] & input_a[1];
  assign popcount25_yqcn_core_105 = ~(input_a[13] ^ input_a[5]);
  assign popcount25_yqcn_core_107 = input_a[14] ^ input_a[18];
  assign popcount25_yqcn_core_109 = ~(input_a[13] ^ input_a[13]);
  assign popcount25_yqcn_core_110 = ~(input_a[5] & input_a[14]);
  assign popcount25_yqcn_core_111 = ~(input_a[3] ^ input_a[12]);
  assign popcount25_yqcn_core_113 = input_a[20] | input_a[16];
  assign popcount25_yqcn_core_114 = ~(input_a[18] & input_a[10]);
  assign popcount25_yqcn_core_115 = ~(input_a[18] & input_a[20]);
  assign popcount25_yqcn_core_117 = input_a[10] ^ input_a[15];
  assign popcount25_yqcn_core_118 = ~input_a[4];
  assign popcount25_yqcn_core_121 = ~(input_a[0] ^ input_a[17]);
  assign popcount25_yqcn_core_123 = ~(input_a[4] ^ input_a[18]);
  assign popcount25_yqcn_core_124 = ~(input_a[8] | input_a[10]);
  assign popcount25_yqcn_core_125 = ~(input_a[0] & input_a[2]);
  assign popcount25_yqcn_core_126 = ~input_a[20];
  assign popcount25_yqcn_core_129 = ~(input_a[7] | input_a[7]);
  assign popcount25_yqcn_core_131 = input_a[11] | input_a[8];
  assign popcount25_yqcn_core_133 = input_a[5] ^ input_a[2];
  assign popcount25_yqcn_core_134 = ~input_a[15];
  assign popcount25_yqcn_core_135 = ~(input_a[16] | input_a[0]);
  assign popcount25_yqcn_core_138 = ~(input_a[21] ^ input_a[19]);
  assign popcount25_yqcn_core_140 = ~(input_a[18] & input_a[3]);
  assign popcount25_yqcn_core_141_not = ~input_a[19];
  assign popcount25_yqcn_core_142 = input_a[22] ^ input_a[23];
  assign popcount25_yqcn_core_143 = input_a[23] | input_a[24];
  assign popcount25_yqcn_core_144 = ~(input_a[13] & input_a[5]);
  assign popcount25_yqcn_core_146 = ~input_a[11];
  assign popcount25_yqcn_core_147 = ~(input_a[9] & input_a[8]);
  assign popcount25_yqcn_core_148 = ~(input_a[12] & input_a[24]);
  assign popcount25_yqcn_core_149 = ~input_a[24];
  assign popcount25_yqcn_core_150 = ~(input_a[22] & input_a[4]);
  assign popcount25_yqcn_core_152 = input_a[13] | input_a[4];
  assign popcount25_yqcn_core_155 = input_a[0] | input_a[0];
  assign popcount25_yqcn_core_156 = ~(input_a[22] & input_a[19]);
  assign popcount25_yqcn_core_157 = ~(input_a[1] ^ input_a[8]);
  assign popcount25_yqcn_core_159 = input_a[12] & input_a[13];
  assign popcount25_yqcn_core_160 = ~(input_a[23] ^ input_a[16]);
  assign popcount25_yqcn_core_163 = ~input_a[19];
  assign popcount25_yqcn_core_165 = ~(input_a[6] | input_a[22]);
  assign popcount25_yqcn_core_167 = input_a[9] | input_a[16];
  assign popcount25_yqcn_core_169 = ~(input_a[23] ^ input_a[6]);
  assign popcount25_yqcn_core_171 = ~(input_a[4] & input_a[2]);
  assign popcount25_yqcn_core_173 = input_a[15] & input_a[20];
  assign popcount25_yqcn_core_175 = ~(input_a[15] | input_a[11]);
  assign popcount25_yqcn_core_178 = input_a[0] ^ input_a[23];
  assign popcount25_yqcn_core_180 = ~(input_a[7] & input_a[19]);
  assign popcount25_yqcn_core_181 = ~(input_a[6] & input_a[10]);
  assign popcount25_yqcn_core_182 = input_a[0] & input_a[16];

  assign popcount25_yqcn_out[0] = input_a[15];
  assign popcount25_yqcn_out[1] = 1'b1;
  assign popcount25_yqcn_out[2] = input_a[6];
  assign popcount25_yqcn_out[3] = 1'b1;
  assign popcount25_yqcn_out[4] = 1'b0;
endmodule