// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.78423
// WCE=38.0
// EP=0.913752%
// Printed PDK parameters:
//  Area=78422932.0
//  Delay=80385632.0
//  Power=3688400.0

module popcount39_gdnl(input [38:0] input_a, output [5:0] popcount39_gdnl_out);
  wire popcount39_gdnl_core_042;
  wire popcount39_gdnl_core_046;
  wire popcount39_gdnl_core_047;
  wire popcount39_gdnl_core_048;
  wire popcount39_gdnl_core_049;
  wire popcount39_gdnl_core_050;
  wire popcount39_gdnl_core_051;
  wire popcount39_gdnl_core_052;
  wire popcount39_gdnl_core_053;
  wire popcount39_gdnl_core_054;
  wire popcount39_gdnl_core_056;
  wire popcount39_gdnl_core_058_not;
  wire popcount39_gdnl_core_060;
  wire popcount39_gdnl_core_061;
  wire popcount39_gdnl_core_062;
  wire popcount39_gdnl_core_063;
  wire popcount39_gdnl_core_064;
  wire popcount39_gdnl_core_065;
  wire popcount39_gdnl_core_066;
  wire popcount39_gdnl_core_067;
  wire popcount39_gdnl_core_068;
  wire popcount39_gdnl_core_070;
  wire popcount39_gdnl_core_072;
  wire popcount39_gdnl_core_076;
  wire popcount39_gdnl_core_077;
  wire popcount39_gdnl_core_083;
  wire popcount39_gdnl_core_084;
  wire popcount39_gdnl_core_085;
  wire popcount39_gdnl_core_086;
  wire popcount39_gdnl_core_089;
  wire popcount39_gdnl_core_090;
  wire popcount39_gdnl_core_091;
  wire popcount39_gdnl_core_092;
  wire popcount39_gdnl_core_093;
  wire popcount39_gdnl_core_094;
  wire popcount39_gdnl_core_095;
  wire popcount39_gdnl_core_096;
  wire popcount39_gdnl_core_097;
  wire popcount39_gdnl_core_098;
  wire popcount39_gdnl_core_099;
  wire popcount39_gdnl_core_100;
  wire popcount39_gdnl_core_101;
  wire popcount39_gdnl_core_102;
  wire popcount39_gdnl_core_103;
  wire popcount39_gdnl_core_104;
  wire popcount39_gdnl_core_105;
  wire popcount39_gdnl_core_106;
  wire popcount39_gdnl_core_107;
  wire popcount39_gdnl_core_108;
  wire popcount39_gdnl_core_109;
  wire popcount39_gdnl_core_110;
  wire popcount39_gdnl_core_111;
  wire popcount39_gdnl_core_112;
  wire popcount39_gdnl_core_113;
  wire popcount39_gdnl_core_114;
  wire popcount39_gdnl_core_115;
  wire popcount39_gdnl_core_116;
  wire popcount39_gdnl_core_117;
  wire popcount39_gdnl_core_119;
  wire popcount39_gdnl_core_124;
  wire popcount39_gdnl_core_125;
  wire popcount39_gdnl_core_129;
  wire popcount39_gdnl_core_131;
  wire popcount39_gdnl_core_132;
  wire popcount39_gdnl_core_134_not;
  wire popcount39_gdnl_core_135_not;
  wire popcount39_gdnl_core_138;
  wire popcount39_gdnl_core_139;
  wire popcount39_gdnl_core_141;
  wire popcount39_gdnl_core_142;
  wire popcount39_gdnl_core_146;
  wire popcount39_gdnl_core_147;
  wire popcount39_gdnl_core_148;
  wire popcount39_gdnl_core_149;
  wire popcount39_gdnl_core_150;
  wire popcount39_gdnl_core_152;
  wire popcount39_gdnl_core_153;
  wire popcount39_gdnl_core_154;
  wire popcount39_gdnl_core_155;
  wire popcount39_gdnl_core_157;
  wire popcount39_gdnl_core_164;
  wire popcount39_gdnl_core_165;
  wire popcount39_gdnl_core_168;
  wire popcount39_gdnl_core_169;
  wire popcount39_gdnl_core_173;
  wire popcount39_gdnl_core_174;
  wire popcount39_gdnl_core_175;
  wire popcount39_gdnl_core_176;
  wire popcount39_gdnl_core_177;
  wire popcount39_gdnl_core_178;
  wire popcount39_gdnl_core_179;
  wire popcount39_gdnl_core_180;
  wire popcount39_gdnl_core_181;
  wire popcount39_gdnl_core_183;
  wire popcount39_gdnl_core_184;
  wire popcount39_gdnl_core_187;
  wire popcount39_gdnl_core_188;
  wire popcount39_gdnl_core_189;
  wire popcount39_gdnl_core_190;
  wire popcount39_gdnl_core_191;
  wire popcount39_gdnl_core_194;
  wire popcount39_gdnl_core_195;
  wire popcount39_gdnl_core_197;
  wire popcount39_gdnl_core_198;
  wire popcount39_gdnl_core_199;
  wire popcount39_gdnl_core_200;
  wire popcount39_gdnl_core_201;
  wire popcount39_gdnl_core_204;
  wire popcount39_gdnl_core_205;
  wire popcount39_gdnl_core_207;
  wire popcount39_gdnl_core_208;
  wire popcount39_gdnl_core_209;
  wire popcount39_gdnl_core_210;
  wire popcount39_gdnl_core_211;
  wire popcount39_gdnl_core_215;
  wire popcount39_gdnl_core_216;
  wire popcount39_gdnl_core_217;
  wire popcount39_gdnl_core_218;
  wire popcount39_gdnl_core_220;
  wire popcount39_gdnl_core_221;
  wire popcount39_gdnl_core_224;
  wire popcount39_gdnl_core_225;
  wire popcount39_gdnl_core_226;
  wire popcount39_gdnl_core_229;
  wire popcount39_gdnl_core_230_not;
  wire popcount39_gdnl_core_233;
  wire popcount39_gdnl_core_234;
  wire popcount39_gdnl_core_235;
  wire popcount39_gdnl_core_237;
  wire popcount39_gdnl_core_238;
  wire popcount39_gdnl_core_241_not;
  wire popcount39_gdnl_core_243;
  wire popcount39_gdnl_core_244;
  wire popcount39_gdnl_core_245;
  wire popcount39_gdnl_core_246;
  wire popcount39_gdnl_core_247;
  wire popcount39_gdnl_core_248;
  wire popcount39_gdnl_core_249;
  wire popcount39_gdnl_core_250;
  wire popcount39_gdnl_core_251;
  wire popcount39_gdnl_core_252;
  wire popcount39_gdnl_core_259;
  wire popcount39_gdnl_core_260;
  wire popcount39_gdnl_core_261;
  wire popcount39_gdnl_core_262;
  wire popcount39_gdnl_core_263;
  wire popcount39_gdnl_core_264;
  wire popcount39_gdnl_core_265;
  wire popcount39_gdnl_core_266;
  wire popcount39_gdnl_core_267;
  wire popcount39_gdnl_core_268;
  wire popcount39_gdnl_core_269;
  wire popcount39_gdnl_core_270;
  wire popcount39_gdnl_core_271;
  wire popcount39_gdnl_core_272;
  wire popcount39_gdnl_core_273;
  wire popcount39_gdnl_core_274;
  wire popcount39_gdnl_core_280_not;
  wire popcount39_gdnl_core_282;
  wire popcount39_gdnl_core_283;
  wire popcount39_gdnl_core_284;
  wire popcount39_gdnl_core_285;
  wire popcount39_gdnl_core_286;
  wire popcount39_gdnl_core_287;
  wire popcount39_gdnl_core_288;
  wire popcount39_gdnl_core_289;
  wire popcount39_gdnl_core_290;
  wire popcount39_gdnl_core_291;
  wire popcount39_gdnl_core_292;
  wire popcount39_gdnl_core_293;
  wire popcount39_gdnl_core_294;
  wire popcount39_gdnl_core_295;
  wire popcount39_gdnl_core_296;
  wire popcount39_gdnl_core_297;
  wire popcount39_gdnl_core_298;
  wire popcount39_gdnl_core_299;
  wire popcount39_gdnl_core_303;
  wire popcount39_gdnl_core_304;
  wire popcount39_gdnl_core_305;
  wire popcount39_gdnl_core_306;

  assign popcount39_gdnl_core_042 = ~input_a[27];
  assign popcount39_gdnl_core_046 = input_a[18] & input_a[24];
  assign popcount39_gdnl_core_047 = input_a[23] ^ input_a[2];
  assign popcount39_gdnl_core_048 = popcount39_gdnl_core_042 & input_a[2];
  assign popcount39_gdnl_core_049 = input_a[4] ^ input_a[13];
  assign popcount39_gdnl_core_050 = input_a[25] & popcount39_gdnl_core_046;
  assign popcount39_gdnl_core_051 = popcount39_gdnl_core_048 | popcount39_gdnl_core_050;
  assign popcount39_gdnl_core_052 = input_a[4] ^ input_a[5];
  assign popcount39_gdnl_core_053 = input_a[4] & input_a[5];
  assign popcount39_gdnl_core_054 = input_a[14] ^ input_a[19];
  assign popcount39_gdnl_core_056 = input_a[15] ^ popcount39_gdnl_core_054;
  assign popcount39_gdnl_core_058_not = ~input_a[7];
  assign popcount39_gdnl_core_060 = popcount39_gdnl_core_052 ^ input_a[28];
  assign popcount39_gdnl_core_061 = popcount39_gdnl_core_052 & input_a[17];
  assign popcount39_gdnl_core_062 = popcount39_gdnl_core_053 ^ popcount39_gdnl_core_058_not;
  assign popcount39_gdnl_core_063 = popcount39_gdnl_core_053 & popcount39_gdnl_core_058_not;
  assign popcount39_gdnl_core_064 = popcount39_gdnl_core_062 ^ input_a[25];
  assign popcount39_gdnl_core_065 = popcount39_gdnl_core_062 & popcount39_gdnl_core_061;
  assign popcount39_gdnl_core_066 = popcount39_gdnl_core_063 | popcount39_gdnl_core_065;
  assign popcount39_gdnl_core_067 = input_a[7] ^ popcount39_gdnl_core_066;
  assign popcount39_gdnl_core_068 = input_a[7] & popcount39_gdnl_core_066;
  assign popcount39_gdnl_core_070 = input_a[0] & input_a[31];
  assign popcount39_gdnl_core_072 = popcount39_gdnl_core_049 & input_a[35];
  assign popcount39_gdnl_core_076 = popcount39_gdnl_core_051 | input_a[32];
  assign popcount39_gdnl_core_077 = popcount39_gdnl_core_051 & popcount39_gdnl_core_067;
  assign popcount39_gdnl_core_083 = input_a[9] ^ input_a[10];
  assign popcount39_gdnl_core_084 = input_a[9] & input_a[10];
  assign popcount39_gdnl_core_085 = input_a[12] ^ input_a[13];
  assign popcount39_gdnl_core_086 = input_a[12] & input_a[23];
  assign popcount39_gdnl_core_089 = ~(popcount39_gdnl_core_086 & input_a[11]);
  assign popcount39_gdnl_core_090 = popcount39_gdnl_core_086 & input_a[11];
  assign popcount39_gdnl_core_091 = input_a[29] ^ input_a[36];
  assign popcount39_gdnl_core_092 = popcount39_gdnl_core_083 & input_a[30];
  assign popcount39_gdnl_core_093 = popcount39_gdnl_core_084 ^ popcount39_gdnl_core_089;
  assign popcount39_gdnl_core_094 = popcount39_gdnl_core_084 & popcount39_gdnl_core_089;
  assign popcount39_gdnl_core_095 = popcount39_gdnl_core_093 ^ input_a[16];
  assign popcount39_gdnl_core_096 = popcount39_gdnl_core_093 & popcount39_gdnl_core_092;
  assign popcount39_gdnl_core_097 = popcount39_gdnl_core_094 | popcount39_gdnl_core_096;
  assign popcount39_gdnl_core_098 = popcount39_gdnl_core_090 ^ popcount39_gdnl_core_097;
  assign popcount39_gdnl_core_099 = popcount39_gdnl_core_090 & popcount39_gdnl_core_097;
  assign popcount39_gdnl_core_100 = input_a[19] | input_a[4];
  assign popcount39_gdnl_core_101 = input_a[14] & input_a[15];
  assign popcount39_gdnl_core_102 = input_a[17] ^ input_a[18];
  assign popcount39_gdnl_core_103 = input_a[17] & input_a[18];
  assign popcount39_gdnl_core_104 = input_a[19] ^ popcount39_gdnl_core_102;
  assign popcount39_gdnl_core_105 = input_a[16] & popcount39_gdnl_core_102;
  assign popcount39_gdnl_core_106 = popcount39_gdnl_core_103 ^ popcount39_gdnl_core_105;
  assign popcount39_gdnl_core_107 = popcount39_gdnl_core_103 & popcount39_gdnl_core_105;
  assign popcount39_gdnl_core_108 = popcount39_gdnl_core_100 ^ popcount39_gdnl_core_104;
  assign popcount39_gdnl_core_109 = popcount39_gdnl_core_100 & popcount39_gdnl_core_104;
  assign popcount39_gdnl_core_110 = input_a[12] | popcount39_gdnl_core_106;
  assign popcount39_gdnl_core_111 = popcount39_gdnl_core_101 & popcount39_gdnl_core_106;
  assign popcount39_gdnl_core_112 = input_a[27] ^ popcount39_gdnl_core_109;
  assign popcount39_gdnl_core_113 = input_a[3] & popcount39_gdnl_core_109;
  assign popcount39_gdnl_core_114 = popcount39_gdnl_core_111 | popcount39_gdnl_core_113;
  assign popcount39_gdnl_core_115 = popcount39_gdnl_core_107 ^ popcount39_gdnl_core_114;
  assign popcount39_gdnl_core_116 = popcount39_gdnl_core_107 & popcount39_gdnl_core_114;
  assign popcount39_gdnl_core_117 = popcount39_gdnl_core_091 ^ popcount39_gdnl_core_108;
  assign popcount39_gdnl_core_119 = ~(input_a[4] & input_a[7]);
  assign popcount39_gdnl_core_124 = popcount39_gdnl_core_098 ^ popcount39_gdnl_core_115;
  assign popcount39_gdnl_core_125 = popcount39_gdnl_core_098 & popcount39_gdnl_core_115;
  assign popcount39_gdnl_core_129 = popcount39_gdnl_core_099 ^ popcount39_gdnl_core_116;
  assign popcount39_gdnl_core_131 = popcount39_gdnl_core_129 ^ popcount39_gdnl_core_125;
  assign popcount39_gdnl_core_132 = popcount39_gdnl_core_129 & popcount39_gdnl_core_125;
  assign popcount39_gdnl_core_134_not = ~popcount39_gdnl_core_117;
  assign popcount39_gdnl_core_135_not = ~popcount39_gdnl_core_117;
  assign popcount39_gdnl_core_138 = ~input_a[3];
  assign popcount39_gdnl_core_139 = input_a[13] & input_a[37];
  assign popcount39_gdnl_core_141 = popcount39_gdnl_core_076 ^ popcount39_gdnl_core_124;
  assign popcount39_gdnl_core_142 = popcount39_gdnl_core_076 & popcount39_gdnl_core_124;
  assign popcount39_gdnl_core_146 = popcount39_gdnl_core_068 ^ popcount39_gdnl_core_131;
  assign popcount39_gdnl_core_147 = popcount39_gdnl_core_068 & input_a[11];
  assign popcount39_gdnl_core_148 = popcount39_gdnl_core_146 | popcount39_gdnl_core_142;
  assign popcount39_gdnl_core_149 = popcount39_gdnl_core_146 & popcount39_gdnl_core_142;
  assign popcount39_gdnl_core_150 = popcount39_gdnl_core_147 | popcount39_gdnl_core_149;
  assign popcount39_gdnl_core_152 = input_a[27] & popcount39_gdnl_core_132;
  assign popcount39_gdnl_core_153 = popcount39_gdnl_core_132 ^ popcount39_gdnl_core_150;
  assign popcount39_gdnl_core_154 = popcount39_gdnl_core_132 & popcount39_gdnl_core_150;
  assign popcount39_gdnl_core_155 = popcount39_gdnl_core_152 | popcount39_gdnl_core_154;
  assign popcount39_gdnl_core_157 = input_a[19] & input_a[20];
  assign popcount39_gdnl_core_164 = input_a[19] ^ input_a[21];
  assign popcount39_gdnl_core_165 = input_a[36] & input_a[21];
  assign popcount39_gdnl_core_168 = popcount39_gdnl_core_157 ^ popcount39_gdnl_core_165;
  assign popcount39_gdnl_core_169 = popcount39_gdnl_core_157 & popcount39_gdnl_core_165;
  assign popcount39_gdnl_core_173 = input_a[24] ^ input_a[25];
  assign popcount39_gdnl_core_174 = input_a[24] & input_a[22];
  assign popcount39_gdnl_core_175 = input_a[35] ^ input_a[21];
  assign popcount39_gdnl_core_176 = input_a[27] & input_a[28];
  assign popcount39_gdnl_core_177 = input_a[32] ^ popcount39_gdnl_core_175;
  assign popcount39_gdnl_core_178 = input_a[26] & popcount39_gdnl_core_175;
  assign popcount39_gdnl_core_179 = popcount39_gdnl_core_176 ^ popcount39_gdnl_core_178;
  assign popcount39_gdnl_core_180 = popcount39_gdnl_core_176 & popcount39_gdnl_core_178;
  assign popcount39_gdnl_core_181 = popcount39_gdnl_core_173 ^ popcount39_gdnl_core_177;
  assign popcount39_gdnl_core_183 = popcount39_gdnl_core_174 ^ popcount39_gdnl_core_179;
  assign popcount39_gdnl_core_184 = popcount39_gdnl_core_174 & input_a[0];
  assign popcount39_gdnl_core_187 = popcount39_gdnl_core_184 | popcount39_gdnl_core_183;
  assign popcount39_gdnl_core_188 = popcount39_gdnl_core_180 ^ popcount39_gdnl_core_187;
  assign popcount39_gdnl_core_189 = popcount39_gdnl_core_180 & popcount39_gdnl_core_187;
  assign popcount39_gdnl_core_190 = popcount39_gdnl_core_164 ^ popcount39_gdnl_core_181;
  assign popcount39_gdnl_core_191 = popcount39_gdnl_core_164 & popcount39_gdnl_core_181;
  assign popcount39_gdnl_core_194 = popcount39_gdnl_core_168 ^ popcount39_gdnl_core_191;
  assign popcount39_gdnl_core_195 = popcount39_gdnl_core_168 & popcount39_gdnl_core_191;
  assign popcount39_gdnl_core_197 = popcount39_gdnl_core_169 ^ popcount39_gdnl_core_188;
  assign popcount39_gdnl_core_198 = popcount39_gdnl_core_169 & popcount39_gdnl_core_188;
  assign popcount39_gdnl_core_199 = popcount39_gdnl_core_197 ^ popcount39_gdnl_core_195;
  assign popcount39_gdnl_core_200 = popcount39_gdnl_core_197 & popcount39_gdnl_core_195;
  assign popcount39_gdnl_core_201 = popcount39_gdnl_core_198 | popcount39_gdnl_core_200;
  assign popcount39_gdnl_core_204 = popcount39_gdnl_core_189 ^ popcount39_gdnl_core_201;
  assign popcount39_gdnl_core_205 = input_a[11] & popcount39_gdnl_core_201;
  assign popcount39_gdnl_core_207 = input_a[29] ^ input_a[30];
  assign popcount39_gdnl_core_208 = input_a[29] & input_a[30];
  assign popcount39_gdnl_core_209 = input_a[32] ^ input_a[33];
  assign popcount39_gdnl_core_210 = input_a[14] & input_a[33];
  assign popcount39_gdnl_core_211 = ~(input_a[31] | input_a[29]);
  assign popcount39_gdnl_core_215 = popcount39_gdnl_core_207 ^ popcount39_gdnl_core_211;
  assign popcount39_gdnl_core_216 = input_a[26] & popcount39_gdnl_core_211;
  assign popcount39_gdnl_core_217 = input_a[23] ^ popcount39_gdnl_core_210;
  assign popcount39_gdnl_core_218 = popcount39_gdnl_core_208 & popcount39_gdnl_core_210;
  assign popcount39_gdnl_core_220 = ~(popcount39_gdnl_core_217 | input_a[34]);
  assign popcount39_gdnl_core_221 = ~(popcount39_gdnl_core_218 & input_a[9]);
  assign popcount39_gdnl_core_224 = input_a[34] ^ input_a[35];
  assign popcount39_gdnl_core_225 = input_a[34] & input_a[37];
  assign popcount39_gdnl_core_226 = input_a[37] ^ input_a[38];
  assign popcount39_gdnl_core_229 = input_a[36] & popcount39_gdnl_core_226;
  assign popcount39_gdnl_core_230_not = ~popcount39_gdnl_core_229;
  assign popcount39_gdnl_core_233 = popcount39_gdnl_core_224 & input_a[12];
  assign popcount39_gdnl_core_234 = popcount39_gdnl_core_225 ^ popcount39_gdnl_core_230_not;
  assign popcount39_gdnl_core_235 = popcount39_gdnl_core_225 & popcount39_gdnl_core_230_not;
  assign popcount39_gdnl_core_237 = input_a[7] & popcount39_gdnl_core_233;
  assign popcount39_gdnl_core_238 = popcount39_gdnl_core_235 | popcount39_gdnl_core_237;
  assign popcount39_gdnl_core_241_not = ~popcount39_gdnl_core_215;
  assign popcount39_gdnl_core_243 = popcount39_gdnl_core_217 ^ popcount39_gdnl_core_234;
  assign popcount39_gdnl_core_244 = popcount39_gdnl_core_217 & popcount39_gdnl_core_234;
  assign popcount39_gdnl_core_245 = popcount39_gdnl_core_243 ^ popcount39_gdnl_core_215;
  assign popcount39_gdnl_core_246 = popcount39_gdnl_core_243 & popcount39_gdnl_core_215;
  assign popcount39_gdnl_core_247 = popcount39_gdnl_core_244 | popcount39_gdnl_core_246;
  assign popcount39_gdnl_core_248 = popcount39_gdnl_core_221 ^ popcount39_gdnl_core_238;
  assign popcount39_gdnl_core_249 = popcount39_gdnl_core_221 & popcount39_gdnl_core_238;
  assign popcount39_gdnl_core_250 = popcount39_gdnl_core_248 ^ popcount39_gdnl_core_247;
  assign popcount39_gdnl_core_251 = popcount39_gdnl_core_248 & popcount39_gdnl_core_247;
  assign popcount39_gdnl_core_252 = popcount39_gdnl_core_249 | popcount39_gdnl_core_251;
  assign popcount39_gdnl_core_259 = popcount39_gdnl_core_190 & popcount39_gdnl_core_241_not;
  assign popcount39_gdnl_core_260 = popcount39_gdnl_core_194 ^ popcount39_gdnl_core_245;
  assign popcount39_gdnl_core_261 = popcount39_gdnl_core_194 & popcount39_gdnl_core_245;
  assign popcount39_gdnl_core_262 = popcount39_gdnl_core_260 ^ popcount39_gdnl_core_259;
  assign popcount39_gdnl_core_263 = popcount39_gdnl_core_260 & popcount39_gdnl_core_259;
  assign popcount39_gdnl_core_264 = popcount39_gdnl_core_261 | popcount39_gdnl_core_263;
  assign popcount39_gdnl_core_265 = popcount39_gdnl_core_199 ^ popcount39_gdnl_core_250;
  assign popcount39_gdnl_core_266 = popcount39_gdnl_core_199 & popcount39_gdnl_core_250;
  assign popcount39_gdnl_core_267 = popcount39_gdnl_core_265 ^ popcount39_gdnl_core_264;
  assign popcount39_gdnl_core_268 = popcount39_gdnl_core_265 & popcount39_gdnl_core_264;
  assign popcount39_gdnl_core_269 = popcount39_gdnl_core_266 | popcount39_gdnl_core_268;
  assign popcount39_gdnl_core_270 = popcount39_gdnl_core_204 ^ popcount39_gdnl_core_252;
  assign popcount39_gdnl_core_271 = popcount39_gdnl_core_204 & popcount39_gdnl_core_252;
  assign popcount39_gdnl_core_272 = popcount39_gdnl_core_270 ^ popcount39_gdnl_core_269;
  assign popcount39_gdnl_core_273 = popcount39_gdnl_core_270 & popcount39_gdnl_core_269;
  assign popcount39_gdnl_core_274 = popcount39_gdnl_core_271 | popcount39_gdnl_core_273;
  assign popcount39_gdnl_core_280_not = ~popcount39_gdnl_core_134_not;
  assign popcount39_gdnl_core_282 = popcount39_gdnl_core_138 ^ popcount39_gdnl_core_262;
  assign popcount39_gdnl_core_283 = popcount39_gdnl_core_138 & popcount39_gdnl_core_262;
  assign popcount39_gdnl_core_284 = popcount39_gdnl_core_282 ^ input_a[12];
  assign popcount39_gdnl_core_285 = popcount39_gdnl_core_282 & popcount39_gdnl_core_134_not;
  assign popcount39_gdnl_core_286 = popcount39_gdnl_core_283 | popcount39_gdnl_core_285;
  assign popcount39_gdnl_core_287 = popcount39_gdnl_core_141 ^ popcount39_gdnl_core_267;
  assign popcount39_gdnl_core_288 = popcount39_gdnl_core_141 & popcount39_gdnl_core_267;
  assign popcount39_gdnl_core_289 = popcount39_gdnl_core_287 ^ popcount39_gdnl_core_286;
  assign popcount39_gdnl_core_290 = popcount39_gdnl_core_287 & popcount39_gdnl_core_286;
  assign popcount39_gdnl_core_291 = popcount39_gdnl_core_288 | popcount39_gdnl_core_290;
  assign popcount39_gdnl_core_292 = popcount39_gdnl_core_148 ^ popcount39_gdnl_core_272;
  assign popcount39_gdnl_core_293 = popcount39_gdnl_core_148 & popcount39_gdnl_core_272;
  assign popcount39_gdnl_core_294 = popcount39_gdnl_core_292 ^ popcount39_gdnl_core_291;
  assign popcount39_gdnl_core_295 = popcount39_gdnl_core_292 & popcount39_gdnl_core_291;
  assign popcount39_gdnl_core_296 = popcount39_gdnl_core_293 | popcount39_gdnl_core_295;
  assign popcount39_gdnl_core_297 = popcount39_gdnl_core_153 ^ popcount39_gdnl_core_274;
  assign popcount39_gdnl_core_298 = popcount39_gdnl_core_153 & popcount39_gdnl_core_274;
  assign popcount39_gdnl_core_299 = popcount39_gdnl_core_297 ^ popcount39_gdnl_core_296;
  assign popcount39_gdnl_core_303 = popcount39_gdnl_core_155 & input_a[7];
  assign popcount39_gdnl_core_304 = popcount39_gdnl_core_155 ^ popcount39_gdnl_core_298;
  assign popcount39_gdnl_core_305 = popcount39_gdnl_core_155 & input_a[18];
  assign popcount39_gdnl_core_306 = ~(input_a[21] | popcount39_gdnl_core_305);

  assign popcount39_gdnl_out[0] = popcount39_gdnl_core_280_not;
  assign popcount39_gdnl_out[1] = popcount39_gdnl_core_153;
  assign popcount39_gdnl_out[2] = popcount39_gdnl_core_289;
  assign popcount39_gdnl_out[3] = popcount39_gdnl_core_294;
  assign popcount39_gdnl_out[4] = popcount39_gdnl_core_299;
  assign popcount39_gdnl_out[5] = popcount39_gdnl_core_304;
endmodule