// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.44973
// WCE=9.0
// EP=0.785622%
// Printed PDK parameters:
//  Area=38166873.0
//  Delay=65419536.0
//  Power=2207600.0

module popcount29_1nbj(input [28:0] input_a, output [4:0] popcount29_1nbj_out);
  wire popcount29_1nbj_core_031_not;
  wire popcount29_1nbj_core_032;
  wire popcount29_1nbj_core_033;
  wire popcount29_1nbj_core_034;
  wire popcount29_1nbj_core_035;
  wire popcount29_1nbj_core_036;
  wire popcount29_1nbj_core_038;
  wire popcount29_1nbj_core_042;
  wire popcount29_1nbj_core_044;
  wire popcount29_1nbj_core_046;
  wire popcount29_1nbj_core_047;
  wire popcount29_1nbj_core_048;
  wire popcount29_1nbj_core_049;
  wire popcount29_1nbj_core_050;
  wire popcount29_1nbj_core_051;
  wire popcount29_1nbj_core_053;
  wire popcount29_1nbj_core_057;
  wire popcount29_1nbj_core_059;
  wire popcount29_1nbj_core_061;
  wire popcount29_1nbj_core_066;
  wire popcount29_1nbj_core_067;
  wire popcount29_1nbj_core_068;
  wire popcount29_1nbj_core_069_not;
  wire popcount29_1nbj_core_070_not;
  wire popcount29_1nbj_core_072;
  wire popcount29_1nbj_core_073;
  wire popcount29_1nbj_core_074;
  wire popcount29_1nbj_core_075;
  wire popcount29_1nbj_core_076;
  wire popcount29_1nbj_core_077;
  wire popcount29_1nbj_core_079;
  wire popcount29_1nbj_core_080;
  wire popcount29_1nbj_core_082;
  wire popcount29_1nbj_core_088;
  wire popcount29_1nbj_core_089;
  wire popcount29_1nbj_core_090;
  wire popcount29_1nbj_core_091;
  wire popcount29_1nbj_core_093;
  wire popcount29_1nbj_core_095;
  wire popcount29_1nbj_core_096;
  wire popcount29_1nbj_core_098;
  wire popcount29_1nbj_core_099;
  wire popcount29_1nbj_core_100;
  wire popcount29_1nbj_core_102;
  wire popcount29_1nbj_core_106;
  wire popcount29_1nbj_core_109;
  wire popcount29_1nbj_core_110;
  wire popcount29_1nbj_core_111;
  wire popcount29_1nbj_core_112;
  wire popcount29_1nbj_core_113;
  wire popcount29_1nbj_core_114;
  wire popcount29_1nbj_core_115;
  wire popcount29_1nbj_core_117;
  wire popcount29_1nbj_core_118;
  wire popcount29_1nbj_core_120;
  wire popcount29_1nbj_core_121;
  wire popcount29_1nbj_core_124;
  wire popcount29_1nbj_core_125;
  wire popcount29_1nbj_core_126;
  wire popcount29_1nbj_core_127;
  wire popcount29_1nbj_core_128;
  wire popcount29_1nbj_core_129;
  wire popcount29_1nbj_core_131;
  wire popcount29_1nbj_core_133;
  wire popcount29_1nbj_core_134;
  wire popcount29_1nbj_core_136;
  wire popcount29_1nbj_core_137;
  wire popcount29_1nbj_core_138;
  wire popcount29_1nbj_core_139;
  wire popcount29_1nbj_core_141;
  wire popcount29_1nbj_core_142;
  wire popcount29_1nbj_core_146;
  wire popcount29_1nbj_core_147;
  wire popcount29_1nbj_core_149;
  wire popcount29_1nbj_core_151;
  wire popcount29_1nbj_core_152;
  wire popcount29_1nbj_core_153;
  wire popcount29_1nbj_core_158;
  wire popcount29_1nbj_core_159;
  wire popcount29_1nbj_core_160;
  wire popcount29_1nbj_core_161;
  wire popcount29_1nbj_core_162;
  wire popcount29_1nbj_core_163;
  wire popcount29_1nbj_core_164;
  wire popcount29_1nbj_core_166;
  wire popcount29_1nbj_core_170;
  wire popcount29_1nbj_core_171;
  wire popcount29_1nbj_core_172;
  wire popcount29_1nbj_core_173;
  wire popcount29_1nbj_core_174;
  wire popcount29_1nbj_core_175;
  wire popcount29_1nbj_core_176;
  wire popcount29_1nbj_core_177;
  wire popcount29_1nbj_core_178;
  wire popcount29_1nbj_core_179;
  wire popcount29_1nbj_core_180;
  wire popcount29_1nbj_core_182_not;
  wire popcount29_1nbj_core_186;
  wire popcount29_1nbj_core_187;
  wire popcount29_1nbj_core_188;
  wire popcount29_1nbj_core_189;
  wire popcount29_1nbj_core_190;
  wire popcount29_1nbj_core_191;
  wire popcount29_1nbj_core_192;
  wire popcount29_1nbj_core_193;
  wire popcount29_1nbj_core_194;
  wire popcount29_1nbj_core_195;
  wire popcount29_1nbj_core_196;
  wire popcount29_1nbj_core_197;
  wire popcount29_1nbj_core_198;
  wire popcount29_1nbj_core_199;
  wire popcount29_1nbj_core_200;
  wire popcount29_1nbj_core_201;
  wire popcount29_1nbj_core_202;
  wire popcount29_1nbj_core_205;
  wire popcount29_1nbj_core_206;
  wire popcount29_1nbj_core_207;

  assign popcount29_1nbj_core_031_not = ~input_a[9];
  assign popcount29_1nbj_core_032 = input_a[24] & input_a[23];
  assign popcount29_1nbj_core_033 = input_a[28] & input_a[28];
  assign popcount29_1nbj_core_034 = input_a[28] & input_a[14];
  assign popcount29_1nbj_core_035 = popcount29_1nbj_core_032 ^ input_a[0];
  assign popcount29_1nbj_core_036 = popcount29_1nbj_core_032 & input_a[0];
  assign popcount29_1nbj_core_038 = input_a[4] & input_a[28];
  assign popcount29_1nbj_core_042 = input_a[8] & input_a[23];
  assign popcount29_1nbj_core_044 = ~(input_a[23] ^ input_a[4]);
  assign popcount29_1nbj_core_046 = ~(input_a[8] | input_a[15]);
  assign popcount29_1nbj_core_047 = ~(input_a[13] | input_a[24]);
  assign popcount29_1nbj_core_048 = input_a[14] & input_a[27];
  assign popcount29_1nbj_core_049 = input_a[5] & input_a[12];
  assign popcount29_1nbj_core_050 = popcount29_1nbj_core_035 ^ popcount29_1nbj_core_038;
  assign popcount29_1nbj_core_051 = popcount29_1nbj_core_035 & popcount29_1nbj_core_038;
  assign popcount29_1nbj_core_053 = ~(input_a[20] & input_a[26]);
  assign popcount29_1nbj_core_057 = popcount29_1nbj_core_036 | popcount29_1nbj_core_051;
  assign popcount29_1nbj_core_059 = input_a[10] & input_a[3];
  assign popcount29_1nbj_core_061 = input_a[21] | input_a[27];
  assign popcount29_1nbj_core_066 = ~(input_a[6] ^ input_a[16]);
  assign popcount29_1nbj_core_067 = ~(input_a[9] | input_a[15]);
  assign popcount29_1nbj_core_068 = ~(input_a[27] | input_a[3]);
  assign popcount29_1nbj_core_069_not = ~input_a[13];
  assign popcount29_1nbj_core_070_not = ~input_a[19];
  assign popcount29_1nbj_core_072 = ~(input_a[17] & input_a[10]);
  assign popcount29_1nbj_core_073 = ~(input_a[26] | input_a[28]);
  assign popcount29_1nbj_core_074 = input_a[12] | input_a[11];
  assign popcount29_1nbj_core_075 = ~input_a[10];
  assign popcount29_1nbj_core_076 = ~(input_a[12] | input_a[6]);
  assign popcount29_1nbj_core_077 = ~input_a[19];
  assign popcount29_1nbj_core_079 = ~(input_a[18] & input_a[13]);
  assign popcount29_1nbj_core_080 = input_a[18] & input_a[13];
  assign popcount29_1nbj_core_082 = input_a[9] & input_a[26];
  assign popcount29_1nbj_core_088 = ~(input_a[3] | input_a[13]);
  assign popcount29_1nbj_core_089 = ~(input_a[7] & input_a[9]);
  assign popcount29_1nbj_core_090 = input_a[15] ^ input_a[17];
  assign popcount29_1nbj_core_091 = popcount29_1nbj_core_050 ^ popcount29_1nbj_core_079;
  assign popcount29_1nbj_core_093 = ~popcount29_1nbj_core_091;
  assign popcount29_1nbj_core_095 = popcount29_1nbj_core_050 | popcount29_1nbj_core_091;
  assign popcount29_1nbj_core_096 = popcount29_1nbj_core_057 ^ popcount29_1nbj_core_080;
  assign popcount29_1nbj_core_098 = popcount29_1nbj_core_096 ^ popcount29_1nbj_core_095;
  assign popcount29_1nbj_core_099 = popcount29_1nbj_core_096 & popcount29_1nbj_core_095;
  assign popcount29_1nbj_core_100 = popcount29_1nbj_core_057 | popcount29_1nbj_core_099;
  assign popcount29_1nbj_core_102 = input_a[8] | input_a[9];
  assign popcount29_1nbj_core_106 = ~(input_a[23] & input_a[1]);
  assign popcount29_1nbj_core_109 = ~(input_a[4] & input_a[13]);
  assign popcount29_1nbj_core_110 = input_a[20] | input_a[16];
  assign popcount29_1nbj_core_111 = input_a[26] | input_a[1];
  assign popcount29_1nbj_core_112 = ~input_a[27];
  assign popcount29_1nbj_core_113 = ~(input_a[1] & input_a[16]);
  assign popcount29_1nbj_core_114 = input_a[18] | input_a[2];
  assign popcount29_1nbj_core_115 = input_a[19] & input_a[16];
  assign popcount29_1nbj_core_117 = input_a[21] | input_a[1];
  assign popcount29_1nbj_core_118 = input_a[8] | popcount29_1nbj_core_115;
  assign popcount29_1nbj_core_120 = popcount29_1nbj_core_118 | input_a[21];
  assign popcount29_1nbj_core_121 = ~input_a[14];
  assign popcount29_1nbj_core_124 = input_a[5] & input_a[17];
  assign popcount29_1nbj_core_125 = ~(popcount29_1nbj_core_110 & popcount29_1nbj_core_120);
  assign popcount29_1nbj_core_126 = popcount29_1nbj_core_110 & popcount29_1nbj_core_120;
  assign popcount29_1nbj_core_127 = popcount29_1nbj_core_125 ^ popcount29_1nbj_core_124;
  assign popcount29_1nbj_core_128 = popcount29_1nbj_core_125 & popcount29_1nbj_core_124;
  assign popcount29_1nbj_core_129 = popcount29_1nbj_core_126 | popcount29_1nbj_core_128;
  assign popcount29_1nbj_core_131 = input_a[5] | input_a[16];
  assign popcount29_1nbj_core_133 = input_a[26] ^ input_a[19];
  assign popcount29_1nbj_core_134 = ~(input_a[5] & input_a[4]);
  assign popcount29_1nbj_core_136 = input_a[6] & input_a[1];
  assign popcount29_1nbj_core_137 = ~(input_a[21] | input_a[18]);
  assign popcount29_1nbj_core_138 = input_a[15] & input_a[11];
  assign popcount29_1nbj_core_139 = ~input_a[26];
  assign popcount29_1nbj_core_141 = popcount29_1nbj_core_136 ^ popcount29_1nbj_core_138;
  assign popcount29_1nbj_core_142 = popcount29_1nbj_core_136 & popcount29_1nbj_core_138;
  assign popcount29_1nbj_core_146 = ~(input_a[6] | input_a[0]);
  assign popcount29_1nbj_core_147 = input_a[10] & input_a[7];
  assign popcount29_1nbj_core_149 = input_a[22] & input_a[12];
  assign popcount29_1nbj_core_151 = input_a[25] & input_a[8];
  assign popcount29_1nbj_core_152 = popcount29_1nbj_core_147 ^ popcount29_1nbj_core_149;
  assign popcount29_1nbj_core_153 = popcount29_1nbj_core_147 & popcount29_1nbj_core_149;
  assign popcount29_1nbj_core_158 = input_a[14] & input_a[25];
  assign popcount29_1nbj_core_159 = popcount29_1nbj_core_141 ^ popcount29_1nbj_core_152;
  assign popcount29_1nbj_core_160 = popcount29_1nbj_core_141 & popcount29_1nbj_core_152;
  assign popcount29_1nbj_core_161 = popcount29_1nbj_core_159 ^ popcount29_1nbj_core_158;
  assign popcount29_1nbj_core_162 = popcount29_1nbj_core_159 & popcount29_1nbj_core_158;
  assign popcount29_1nbj_core_163 = popcount29_1nbj_core_160 | popcount29_1nbj_core_162;
  assign popcount29_1nbj_core_164 = popcount29_1nbj_core_142 | popcount29_1nbj_core_153;
  assign popcount29_1nbj_core_166 = popcount29_1nbj_core_164 | popcount29_1nbj_core_163;
  assign popcount29_1nbj_core_170 = input_a[26] & input_a[9];
  assign popcount29_1nbj_core_171 = popcount29_1nbj_core_127 ^ popcount29_1nbj_core_161;
  assign popcount29_1nbj_core_172 = popcount29_1nbj_core_127 & popcount29_1nbj_core_161;
  assign popcount29_1nbj_core_173 = popcount29_1nbj_core_171 ^ popcount29_1nbj_core_170;
  assign popcount29_1nbj_core_174 = popcount29_1nbj_core_171 & popcount29_1nbj_core_170;
  assign popcount29_1nbj_core_175 = popcount29_1nbj_core_172 | popcount29_1nbj_core_174;
  assign popcount29_1nbj_core_176 = popcount29_1nbj_core_129 ^ popcount29_1nbj_core_166;
  assign popcount29_1nbj_core_177 = popcount29_1nbj_core_129 & popcount29_1nbj_core_166;
  assign popcount29_1nbj_core_178 = popcount29_1nbj_core_176 ^ popcount29_1nbj_core_175;
  assign popcount29_1nbj_core_179 = popcount29_1nbj_core_176 & popcount29_1nbj_core_175;
  assign popcount29_1nbj_core_180 = popcount29_1nbj_core_177 | popcount29_1nbj_core_179;
  assign popcount29_1nbj_core_182_not = ~input_a[6];
  assign popcount29_1nbj_core_186 = ~(input_a[0] & input_a[13]);
  assign popcount29_1nbj_core_187 = input_a[3] & input_a[27];
  assign popcount29_1nbj_core_188 = popcount29_1nbj_core_093 ^ popcount29_1nbj_core_173;
  assign popcount29_1nbj_core_189 = popcount29_1nbj_core_093 & popcount29_1nbj_core_173;
  assign popcount29_1nbj_core_190 = popcount29_1nbj_core_188 ^ popcount29_1nbj_core_187;
  assign popcount29_1nbj_core_191 = popcount29_1nbj_core_188 & popcount29_1nbj_core_187;
  assign popcount29_1nbj_core_192 = popcount29_1nbj_core_189 | popcount29_1nbj_core_191;
  assign popcount29_1nbj_core_193 = popcount29_1nbj_core_098 ^ popcount29_1nbj_core_178;
  assign popcount29_1nbj_core_194 = popcount29_1nbj_core_098 & popcount29_1nbj_core_178;
  assign popcount29_1nbj_core_195 = popcount29_1nbj_core_193 ^ popcount29_1nbj_core_192;
  assign popcount29_1nbj_core_196 = popcount29_1nbj_core_193 & popcount29_1nbj_core_192;
  assign popcount29_1nbj_core_197 = popcount29_1nbj_core_194 | popcount29_1nbj_core_196;
  assign popcount29_1nbj_core_198 = popcount29_1nbj_core_100 ^ popcount29_1nbj_core_180;
  assign popcount29_1nbj_core_199 = popcount29_1nbj_core_100 & popcount29_1nbj_core_180;
  assign popcount29_1nbj_core_200 = popcount29_1nbj_core_198 ^ popcount29_1nbj_core_197;
  assign popcount29_1nbj_core_201 = popcount29_1nbj_core_198 & popcount29_1nbj_core_197;
  assign popcount29_1nbj_core_202 = popcount29_1nbj_core_199 | popcount29_1nbj_core_201;
  assign popcount29_1nbj_core_205 = input_a[8] | input_a[22];
  assign popcount29_1nbj_core_206 = input_a[24] & input_a[21];
  assign popcount29_1nbj_core_207 = ~(input_a[18] | input_a[0]);

  assign popcount29_1nbj_out[0] = popcount29_1nbj_core_200;
  assign popcount29_1nbj_out[1] = popcount29_1nbj_core_190;
  assign popcount29_1nbj_out[2] = popcount29_1nbj_core_195;
  assign popcount29_1nbj_out[3] = popcount29_1nbj_core_200;
  assign popcount29_1nbj_out[4] = popcount29_1nbj_core_202;
endmodule