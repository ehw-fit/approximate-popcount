// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.54028
// WCE=10.0
// EP=0.798672%
// Printed PDK parameters:
//  Area=37770884.0
//  Delay=61958700.0
//  Power=1636100.0

module popcount31_193u(input [30:0] input_a, output [4:0] popcount31_193u_out);
  wire popcount31_193u_core_033;
  wire popcount31_193u_core_034;
  wire popcount31_193u_core_035;
  wire popcount31_193u_core_036;
  wire popcount31_193u_core_037;
  wire popcount31_193u_core_039;
  wire popcount31_193u_core_040;
  wire popcount31_193u_core_042;
  wire popcount31_193u_core_045;
  wire popcount31_193u_core_047;
  wire popcount31_193u_core_048;
  wire popcount31_193u_core_052;
  wire popcount31_193u_core_053;
  wire popcount31_193u_core_055;
  wire popcount31_193u_core_058;
  wire popcount31_193u_core_059;
  wire popcount31_193u_core_061;
  wire popcount31_193u_core_062;
  wire popcount31_193u_core_063;
  wire popcount31_193u_core_064;
  wire popcount31_193u_core_065;
  wire popcount31_193u_core_066;
  wire popcount31_193u_core_067;
  wire popcount31_193u_core_068;
  wire popcount31_193u_core_069;
  wire popcount31_193u_core_071;
  wire popcount31_193u_core_072;
  wire popcount31_193u_core_073;
  wire popcount31_193u_core_074;
  wire popcount31_193u_core_075;
  wire popcount31_193u_core_076;
  wire popcount31_193u_core_082;
  wire popcount31_193u_core_083;
  wire popcount31_193u_core_084;
  wire popcount31_193u_core_086;
  wire popcount31_193u_core_087;
  wire popcount31_193u_core_088;
  wire popcount31_193u_core_091;
  wire popcount31_193u_core_093;
  wire popcount31_193u_core_094;
  wire popcount31_193u_core_096;
  wire popcount31_193u_core_097;
  wire popcount31_193u_core_098;
  wire popcount31_193u_core_099;
  wire popcount31_193u_core_100;
  wire popcount31_193u_core_101;
  wire popcount31_193u_core_102;
  wire popcount31_193u_core_103;
  wire popcount31_193u_core_105;
  wire popcount31_193u_core_106;
  wire popcount31_193u_core_107;
  wire popcount31_193u_core_111;
  wire popcount31_193u_core_112;
  wire popcount31_193u_core_115;
  wire popcount31_193u_core_116;
  wire popcount31_193u_core_117;
  wire popcount31_193u_core_119;
  wire popcount31_193u_core_120;
  wire popcount31_193u_core_122;
  wire popcount31_193u_core_123;
  wire popcount31_193u_core_124;
  wire popcount31_193u_core_128;
  wire popcount31_193u_core_130;
  wire popcount31_193u_core_131;
  wire popcount31_193u_core_132;
  wire popcount31_193u_core_136;
  wire popcount31_193u_core_137;
  wire popcount31_193u_core_138;
  wire popcount31_193u_core_139;
  wire popcount31_193u_core_140;
  wire popcount31_193u_core_141;
  wire popcount31_193u_core_143;
  wire popcount31_193u_core_146;
  wire popcount31_193u_core_147;
  wire popcount31_193u_core_148;
  wire popcount31_193u_core_149;
  wire popcount31_193u_core_150;
  wire popcount31_193u_core_152;
  wire popcount31_193u_core_153;
  wire popcount31_193u_core_154;
  wire popcount31_193u_core_155;
  wire popcount31_193u_core_156;
  wire popcount31_193u_core_158;
  wire popcount31_193u_core_161;
  wire popcount31_193u_core_162;
  wire popcount31_193u_core_163_not;
  wire popcount31_193u_core_165;
  wire popcount31_193u_core_168;
  wire popcount31_193u_core_169;
  wire popcount31_193u_core_170;
  wire popcount31_193u_core_171;
  wire popcount31_193u_core_172;
  wire popcount31_193u_core_177_not;
  wire popcount31_193u_core_178;
  wire popcount31_193u_core_179;
  wire popcount31_193u_core_181;
  wire popcount31_193u_core_183;
  wire popcount31_193u_core_184;
  wire popcount31_193u_core_186;
  wire popcount31_193u_core_188;
  wire popcount31_193u_core_189;
  wire popcount31_193u_core_190;
  wire popcount31_193u_core_191;
  wire popcount31_193u_core_192;
  wire popcount31_193u_core_196;
  wire popcount31_193u_core_197;
  wire popcount31_193u_core_198_not;
  wire popcount31_193u_core_200;
  wire popcount31_193u_core_201;
  wire popcount31_193u_core_202;
  wire popcount31_193u_core_203;
  wire popcount31_193u_core_204;
  wire popcount31_193u_core_205;
  wire popcount31_193u_core_206;
  wire popcount31_193u_core_207;
  wire popcount31_193u_core_208;
  wire popcount31_193u_core_209;
  wire popcount31_193u_core_210;
  wire popcount31_193u_core_211;
  wire popcount31_193u_core_212;
  wire popcount31_193u_core_213;
  wire popcount31_193u_core_214;
  wire popcount31_193u_core_215;
  wire popcount31_193u_core_216;
  wire popcount31_193u_core_217;
  wire popcount31_193u_core_218_not;
  wire popcount31_193u_core_219;

  assign popcount31_193u_core_033 = ~(input_a[21] | input_a[15]);
  assign popcount31_193u_core_034 = input_a[28] & input_a[3];
  assign popcount31_193u_core_035 = ~(input_a[20] | input_a[24]);
  assign popcount31_193u_core_036 = input_a[26] & input_a[23];
  assign popcount31_193u_core_037 = input_a[16] | popcount31_193u_core_036;
  assign popcount31_193u_core_039 = input_a[16] & input_a[29];
  assign popcount31_193u_core_040 = input_a[15] & input_a[20];
  assign popcount31_193u_core_042 = input_a[7] & input_a[2];
  assign popcount31_193u_core_045 = popcount31_193u_core_040 | popcount31_193u_core_042;
  assign popcount31_193u_core_047 = popcount31_193u_core_045 ^ input_a[5];
  assign popcount31_193u_core_048 = popcount31_193u_core_045 & input_a[5];
  assign popcount31_193u_core_052 = popcount31_193u_core_037 ^ popcount31_193u_core_047;
  assign popcount31_193u_core_053 = popcount31_193u_core_037 & popcount31_193u_core_047;
  assign popcount31_193u_core_055 = input_a[27] ^ input_a[18];
  assign popcount31_193u_core_058 = input_a[30] | input_a[7];
  assign popcount31_193u_core_059 = popcount31_193u_core_048 | popcount31_193u_core_053;
  assign popcount31_193u_core_061 = ~(input_a[1] & input_a[5]);
  assign popcount31_193u_core_062 = ~(input_a[4] & input_a[28]);
  assign popcount31_193u_core_063 = ~(input_a[24] & input_a[27]);
  assign popcount31_193u_core_064 = ~(input_a[16] | input_a[28]);
  assign popcount31_193u_core_065 = ~input_a[1];
  assign popcount31_193u_core_066 = ~popcount31_193u_core_062;
  assign popcount31_193u_core_067 = ~(input_a[19] & input_a[9]);
  assign popcount31_193u_core_068 = ~(input_a[1] & input_a[19]);
  assign popcount31_193u_core_069 = ~input_a[12];
  assign popcount31_193u_core_071 = input_a[14] & input_a[1];
  assign popcount31_193u_core_072 = ~(input_a[18] ^ input_a[25]);
  assign popcount31_193u_core_073 = ~(input_a[30] ^ input_a[25]);
  assign popcount31_193u_core_074 = input_a[2] | input_a[22];
  assign popcount31_193u_core_075 = input_a[3] ^ input_a[29];
  assign popcount31_193u_core_076 = ~input_a[8];
  assign popcount31_193u_core_082 = input_a[22] | input_a[11];
  assign popcount31_193u_core_083 = ~(input_a[17] ^ input_a[21]);
  assign popcount31_193u_core_084 = ~input_a[4];
  assign popcount31_193u_core_086 = ~popcount31_193u_core_068;
  assign popcount31_193u_core_087 = ~input_a[24];
  assign popcount31_193u_core_088 = popcount31_193u_core_086 | popcount31_193u_core_066;
  assign popcount31_193u_core_091 = ~(input_a[22] | input_a[23]);
  assign popcount31_193u_core_093 = ~(input_a[8] ^ input_a[12]);
  assign popcount31_193u_core_094 = ~(input_a[18] | input_a[9]);
  assign popcount31_193u_core_096 = ~(input_a[5] ^ input_a[10]);
  assign popcount31_193u_core_097 = input_a[9] & input_a[17];
  assign popcount31_193u_core_098 = popcount31_193u_core_052 ^ popcount31_193u_core_088;
  assign popcount31_193u_core_099 = popcount31_193u_core_052 & popcount31_193u_core_088;
  assign popcount31_193u_core_100 = popcount31_193u_core_098 ^ popcount31_193u_core_097;
  assign popcount31_193u_core_101 = popcount31_193u_core_098 & popcount31_193u_core_097;
  assign popcount31_193u_core_102 = popcount31_193u_core_099 | popcount31_193u_core_101;
  assign popcount31_193u_core_103 = ~popcount31_193u_core_059;
  assign popcount31_193u_core_105 = popcount31_193u_core_103 ^ popcount31_193u_core_102;
  assign popcount31_193u_core_106 = popcount31_193u_core_103 & popcount31_193u_core_102;
  assign popcount31_193u_core_107 = popcount31_193u_core_059 | popcount31_193u_core_106;
  assign popcount31_193u_core_111 = input_a[12] | input_a[13];
  assign popcount31_193u_core_112 = ~(input_a[10] | input_a[5]);
  assign popcount31_193u_core_115 = ~(input_a[12] & input_a[21]);
  assign popcount31_193u_core_116 = ~input_a[14];
  assign popcount31_193u_core_117 = input_a[24] & input_a[16];
  assign popcount31_193u_core_119 = input_a[24] | input_a[0];
  assign popcount31_193u_core_120 = ~(input_a[25] ^ input_a[15]);
  assign popcount31_193u_core_122 = ~(input_a[18] ^ input_a[14]);
  assign popcount31_193u_core_123 = ~(input_a[8] & input_a[23]);
  assign popcount31_193u_core_124 = input_a[0] ^ input_a[2];
  assign popcount31_193u_core_128 = ~(input_a[11] | input_a[27]);
  assign popcount31_193u_core_130 = input_a[10] | input_a[17];
  assign popcount31_193u_core_131 = input_a[24] | input_a[22];
  assign popcount31_193u_core_132 = input_a[30] | input_a[11];
  assign popcount31_193u_core_136 = input_a[10] & input_a[27];
  assign popcount31_193u_core_137 = ~(popcount31_193u_core_119 & popcount31_193u_core_132);
  assign popcount31_193u_core_138 = popcount31_193u_core_119 & popcount31_193u_core_132;
  assign popcount31_193u_core_139 = popcount31_193u_core_137 ^ popcount31_193u_core_136;
  assign popcount31_193u_core_140 = input_a[27] & input_a[10];
  assign popcount31_193u_core_141 = popcount31_193u_core_138 | popcount31_193u_core_140;
  assign popcount31_193u_core_143 = input_a[5] & input_a[18];
  assign popcount31_193u_core_146 = ~(input_a[3] ^ input_a[0]);
  assign popcount31_193u_core_147 = ~(input_a[28] | input_a[28]);
  assign popcount31_193u_core_148 = input_a[8] & input_a[25];
  assign popcount31_193u_core_149 = ~(input_a[8] | input_a[27]);
  assign popcount31_193u_core_150 = input_a[3] & input_a[12];
  assign popcount31_193u_core_152 = input_a[21] & input_a[22];
  assign popcount31_193u_core_153 = popcount31_193u_core_148 ^ popcount31_193u_core_150;
  assign popcount31_193u_core_154 = popcount31_193u_core_148 & popcount31_193u_core_150;
  assign popcount31_193u_core_155 = popcount31_193u_core_153 | popcount31_193u_core_152;
  assign popcount31_193u_core_156 = input_a[10] & input_a[18];
  assign popcount31_193u_core_158 = ~input_a[2];
  assign popcount31_193u_core_161 = input_a[13] & input_a[18];
  assign popcount31_193u_core_162 = input_a[29] ^ input_a[26];
  assign popcount31_193u_core_163_not = ~input_a[7];
  assign popcount31_193u_core_165 = ~(input_a[28] | input_a[16]);
  assign popcount31_193u_core_168 = input_a[26] ^ input_a[21];
  assign popcount31_193u_core_169 = input_a[14] & input_a[15];
  assign popcount31_193u_core_170 = input_a[8] ^ input_a[29];
  assign popcount31_193u_core_171 = popcount31_193u_core_155 ^ popcount31_193u_core_161;
  assign popcount31_193u_core_172 = popcount31_193u_core_155 & popcount31_193u_core_161;
  assign popcount31_193u_core_177_not = ~input_a[14];
  assign popcount31_193u_core_178 = popcount31_193u_core_154 | popcount31_193u_core_172;
  assign popcount31_193u_core_179 = ~(input_a[26] | input_a[9]);
  assign popcount31_193u_core_181 = ~(input_a[19] & input_a[29]);
  assign popcount31_193u_core_183 = popcount31_193u_core_139 ^ popcount31_193u_core_171;
  assign popcount31_193u_core_184 = popcount31_193u_core_139 & popcount31_193u_core_171;
  assign popcount31_193u_core_186 = ~(input_a[29] & input_a[18]);
  assign popcount31_193u_core_188 = popcount31_193u_core_141 ^ popcount31_193u_core_178;
  assign popcount31_193u_core_189 = popcount31_193u_core_141 & popcount31_193u_core_178;
  assign popcount31_193u_core_190 = popcount31_193u_core_188 ^ popcount31_193u_core_184;
  assign popcount31_193u_core_191 = popcount31_193u_core_188 & popcount31_193u_core_184;
  assign popcount31_193u_core_192 = popcount31_193u_core_189 | popcount31_193u_core_191;
  assign popcount31_193u_core_196 = ~(input_a[12] | input_a[2]);
  assign popcount31_193u_core_197 = input_a[5] & input_a[3];
  assign popcount31_193u_core_198_not = ~input_a[6];
  assign popcount31_193u_core_200 = popcount31_193u_core_100 ^ popcount31_193u_core_183;
  assign popcount31_193u_core_201 = popcount31_193u_core_100 & popcount31_193u_core_183;
  assign popcount31_193u_core_202 = popcount31_193u_core_200 ^ input_a[14];
  assign popcount31_193u_core_203 = popcount31_193u_core_200 & input_a[14];
  assign popcount31_193u_core_204 = popcount31_193u_core_201 | popcount31_193u_core_203;
  assign popcount31_193u_core_205 = popcount31_193u_core_105 ^ popcount31_193u_core_190;
  assign popcount31_193u_core_206 = popcount31_193u_core_105 & popcount31_193u_core_190;
  assign popcount31_193u_core_207 = popcount31_193u_core_205 ^ popcount31_193u_core_204;
  assign popcount31_193u_core_208 = popcount31_193u_core_205 & popcount31_193u_core_204;
  assign popcount31_193u_core_209 = popcount31_193u_core_206 | popcount31_193u_core_208;
  assign popcount31_193u_core_210 = popcount31_193u_core_107 ^ popcount31_193u_core_192;
  assign popcount31_193u_core_211 = popcount31_193u_core_107 & popcount31_193u_core_192;
  assign popcount31_193u_core_212 = popcount31_193u_core_210 ^ popcount31_193u_core_209;
  assign popcount31_193u_core_213 = popcount31_193u_core_210 & popcount31_193u_core_209;
  assign popcount31_193u_core_214 = popcount31_193u_core_211 | popcount31_193u_core_213;
  assign popcount31_193u_core_215 = ~(input_a[27] ^ input_a[7]);
  assign popcount31_193u_core_216 = ~(input_a[21] ^ input_a[15]);
  assign popcount31_193u_core_217 = input_a[13] ^ input_a[11];
  assign popcount31_193u_core_218_not = ~input_a[13];
  assign popcount31_193u_core_219 = input_a[2] | input_a[29];

  assign popcount31_193u_out[0] = popcount31_193u_core_212;
  assign popcount31_193u_out[1] = popcount31_193u_core_202;
  assign popcount31_193u_out[2] = popcount31_193u_core_207;
  assign popcount31_193u_out[3] = popcount31_193u_core_212;
  assign popcount31_193u_out[4] = popcount31_193u_core_214;
endmodule