// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.8865
// WCE=14.0
// EP=0.834608%
// Printed PDK parameters:
//  Area=36776600.0
//  Delay=64881052.0
//  Power=1919000.0

module popcount38_wm2a(input [37:0] input_a, output [5:0] popcount38_wm2a_out);
  wire popcount38_wm2a_core_041;
  wire popcount38_wm2a_core_042;
  wire popcount38_wm2a_core_048;
  wire popcount38_wm2a_core_051_not;
  wire popcount38_wm2a_core_052;
  wire popcount38_wm2a_core_053;
  wire popcount38_wm2a_core_054;
  wire popcount38_wm2a_core_055;
  wire popcount38_wm2a_core_056;
  wire popcount38_wm2a_core_058;
  wire popcount38_wm2a_core_059;
  wire popcount38_wm2a_core_060;
  wire popcount38_wm2a_core_061;
  wire popcount38_wm2a_core_062;
  wire popcount38_wm2a_core_064;
  wire popcount38_wm2a_core_065;
  wire popcount38_wm2a_core_066;
  wire popcount38_wm2a_core_068;
  wire popcount38_wm2a_core_069;
  wire popcount38_wm2a_core_070;
  wire popcount38_wm2a_core_073;
  wire popcount38_wm2a_core_078;
  wire popcount38_wm2a_core_079;
  wire popcount38_wm2a_core_083;
  wire popcount38_wm2a_core_084;
  wire popcount38_wm2a_core_086;
  wire popcount38_wm2a_core_087;
  wire popcount38_wm2a_core_090;
  wire popcount38_wm2a_core_092;
  wire popcount38_wm2a_core_094;
  wire popcount38_wm2a_core_095;
  wire popcount38_wm2a_core_099;
  wire popcount38_wm2a_core_100;
  wire popcount38_wm2a_core_101;
  wire popcount38_wm2a_core_102;
  wire popcount38_wm2a_core_103;
  wire popcount38_wm2a_core_104;
  wire popcount38_wm2a_core_105;
  wire popcount38_wm2a_core_116;
  wire popcount38_wm2a_core_118;
  wire popcount38_wm2a_core_119;
  wire popcount38_wm2a_core_121;
  wire popcount38_wm2a_core_122;
  wire popcount38_wm2a_core_123;
  wire popcount38_wm2a_core_124;
  wire popcount38_wm2a_core_126;
  wire popcount38_wm2a_core_127;
  wire popcount38_wm2a_core_131;
  wire popcount38_wm2a_core_132;
  wire popcount38_wm2a_core_134;
  wire popcount38_wm2a_core_135;
  wire popcount38_wm2a_core_137;
  wire popcount38_wm2a_core_139;
  wire popcount38_wm2a_core_140;
  wire popcount38_wm2a_core_142;
  wire popcount38_wm2a_core_143;
  wire popcount38_wm2a_core_144;
  wire popcount38_wm2a_core_146;
  wire popcount38_wm2a_core_150;
  wire popcount38_wm2a_core_151;
  wire popcount38_wm2a_core_152;
  wire popcount38_wm2a_core_153;
  wire popcount38_wm2a_core_156;
  wire popcount38_wm2a_core_157;
  wire popcount38_wm2a_core_160;
  wire popcount38_wm2a_core_161;
  wire popcount38_wm2a_core_162;
  wire popcount38_wm2a_core_163;
  wire popcount38_wm2a_core_164;
  wire popcount38_wm2a_core_165;
  wire popcount38_wm2a_core_166;
  wire popcount38_wm2a_core_167;
  wire popcount38_wm2a_core_168;
  wire popcount38_wm2a_core_170;
  wire popcount38_wm2a_core_171;
  wire popcount38_wm2a_core_173;
  wire popcount38_wm2a_core_175;
  wire popcount38_wm2a_core_176;
  wire popcount38_wm2a_core_177;
  wire popcount38_wm2a_core_183;
  wire popcount38_wm2a_core_184;
  wire popcount38_wm2a_core_185;
  wire popcount38_wm2a_core_186;
  wire popcount38_wm2a_core_188;
  wire popcount38_wm2a_core_192;
  wire popcount38_wm2a_core_193;
  wire popcount38_wm2a_core_194;
  wire popcount38_wm2a_core_196;
  wire popcount38_wm2a_core_198;
  wire popcount38_wm2a_core_199;
  wire popcount38_wm2a_core_200;
  wire popcount38_wm2a_core_201;
  wire popcount38_wm2a_core_202;
  wire popcount38_wm2a_core_203;
  wire popcount38_wm2a_core_205;
  wire popcount38_wm2a_core_206;
  wire popcount38_wm2a_core_207;
  wire popcount38_wm2a_core_211;
  wire popcount38_wm2a_core_213;
  wire popcount38_wm2a_core_214;
  wire popcount38_wm2a_core_215;
  wire popcount38_wm2a_core_216;
  wire popcount38_wm2a_core_218;
  wire popcount38_wm2a_core_219;
  wire popcount38_wm2a_core_220;
  wire popcount38_wm2a_core_222;
  wire popcount38_wm2a_core_223;
  wire popcount38_wm2a_core_224;
  wire popcount38_wm2a_core_225;
  wire popcount38_wm2a_core_226;
  wire popcount38_wm2a_core_227;
  wire popcount38_wm2a_core_228;
  wire popcount38_wm2a_core_230;
  wire popcount38_wm2a_core_231;
  wire popcount38_wm2a_core_232;
  wire popcount38_wm2a_core_233_not;
  wire popcount38_wm2a_core_235;
  wire popcount38_wm2a_core_236;
  wire popcount38_wm2a_core_237;
  wire popcount38_wm2a_core_240;
  wire popcount38_wm2a_core_241;
  wire popcount38_wm2a_core_246;
  wire popcount38_wm2a_core_247;
  wire popcount38_wm2a_core_249;
  wire popcount38_wm2a_core_250;
  wire popcount38_wm2a_core_251;
  wire popcount38_wm2a_core_253;
  wire popcount38_wm2a_core_255;
  wire popcount38_wm2a_core_256;
  wire popcount38_wm2a_core_257;
  wire popcount38_wm2a_core_258;
  wire popcount38_wm2a_core_259;
  wire popcount38_wm2a_core_261;
  wire popcount38_wm2a_core_262;
  wire popcount38_wm2a_core_263;
  wire popcount38_wm2a_core_264;
  wire popcount38_wm2a_core_265;
  wire popcount38_wm2a_core_266;
  wire popcount38_wm2a_core_267;
  wire popcount38_wm2a_core_268;
  wire popcount38_wm2a_core_269;
  wire popcount38_wm2a_core_270;
  wire popcount38_wm2a_core_272;
  wire popcount38_wm2a_core_273;
  wire popcount38_wm2a_core_274;
  wire popcount38_wm2a_core_275;
  wire popcount38_wm2a_core_276;
  wire popcount38_wm2a_core_277;
  wire popcount38_wm2a_core_278;
  wire popcount38_wm2a_core_279;
  wire popcount38_wm2a_core_280;
  wire popcount38_wm2a_core_281;
  wire popcount38_wm2a_core_282_not;
  wire popcount38_wm2a_core_284;
  wire popcount38_wm2a_core_285;
  wire popcount38_wm2a_core_286;
  wire popcount38_wm2a_core_288;
  wire popcount38_wm2a_core_290;
  wire popcount38_wm2a_core_291;
  wire popcount38_wm2a_core_293;
  wire popcount38_wm2a_core_294;
  wire popcount38_wm2a_core_296;

  assign popcount38_wm2a_core_041 = ~(input_a[13] ^ input_a[18]);
  assign popcount38_wm2a_core_042 = ~(input_a[23] & input_a[25]);
  assign popcount38_wm2a_core_048 = input_a[11] | input_a[26];
  assign popcount38_wm2a_core_051_not = ~input_a[26];
  assign popcount38_wm2a_core_052 = input_a[5] & input_a[35];
  assign popcount38_wm2a_core_053 = input_a[7] & input_a[31];
  assign popcount38_wm2a_core_054 = input_a[2] & input_a[9];
  assign popcount38_wm2a_core_055 = input_a[30] ^ input_a[0];
  assign popcount38_wm2a_core_056 = input_a[9] & input_a[0];
  assign popcount38_wm2a_core_058 = ~input_a[22];
  assign popcount38_wm2a_core_059 = input_a[26] ^ input_a[2];
  assign popcount38_wm2a_core_060 = ~(input_a[24] & input_a[33]);
  assign popcount38_wm2a_core_061 = popcount38_wm2a_core_052 | popcount38_wm2a_core_054;
  assign popcount38_wm2a_core_062 = input_a[14] & input_a[6];
  assign popcount38_wm2a_core_064 = input_a[23] ^ input_a[6];
  assign popcount38_wm2a_core_065 = input_a[35] | input_a[25];
  assign popcount38_wm2a_core_066 = input_a[18] ^ input_a[0];
  assign popcount38_wm2a_core_068 = input_a[9] & input_a[17];
  assign popcount38_wm2a_core_069 = ~(input_a[20] ^ input_a[34]);
  assign popcount38_wm2a_core_070 = ~(popcount38_wm2a_core_048 & popcount38_wm2a_core_061);
  assign popcount38_wm2a_core_073 = ~popcount38_wm2a_core_070;
  assign popcount38_wm2a_core_078 = input_a[20] | input_a[34];
  assign popcount38_wm2a_core_079 = ~(input_a[16] & input_a[37]);
  assign popcount38_wm2a_core_083 = ~(input_a[11] | input_a[9]);
  assign popcount38_wm2a_core_084 = ~(input_a[19] ^ input_a[35]);
  assign popcount38_wm2a_core_086 = ~(input_a[20] & input_a[27]);
  assign popcount38_wm2a_core_087 = input_a[34] & input_a[8];
  assign popcount38_wm2a_core_090 = input_a[14] ^ input_a[28];
  assign popcount38_wm2a_core_092 = input_a[32] & input_a[31];
  assign popcount38_wm2a_core_094 = ~(popcount38_wm2a_core_092 & input_a[18]);
  assign popcount38_wm2a_core_095 = popcount38_wm2a_core_092 & input_a[18];
  assign popcount38_wm2a_core_099 = ~(input_a[14] & input_a[15]);
  assign popcount38_wm2a_core_100 = input_a[14] & input_a[15];
  assign popcount38_wm2a_core_101 = input_a[31] ^ input_a[21];
  assign popcount38_wm2a_core_102 = ~(input_a[34] ^ input_a[14]);
  assign popcount38_wm2a_core_103 = ~(input_a[23] & input_a[23]);
  assign popcount38_wm2a_core_104 = ~(input_a[26] ^ input_a[35]);
  assign popcount38_wm2a_core_105 = ~(input_a[14] ^ input_a[9]);
  assign popcount38_wm2a_core_116 = ~input_a[7];
  assign popcount38_wm2a_core_118 = popcount38_wm2a_core_094 ^ popcount38_wm2a_core_099;
  assign popcount38_wm2a_core_119 = ~(input_a[13] ^ input_a[11]);
  assign popcount38_wm2a_core_121 = ~input_a[28];
  assign popcount38_wm2a_core_122 = ~(input_a[7] ^ input_a[6]);
  assign popcount38_wm2a_core_123 = ~(popcount38_wm2a_core_095 & popcount38_wm2a_core_100);
  assign popcount38_wm2a_core_124 = ~(input_a[10] & input_a[20]);
  assign popcount38_wm2a_core_126 = ~(input_a[17] & input_a[32]);
  assign popcount38_wm2a_core_127 = input_a[20] ^ input_a[36];
  assign popcount38_wm2a_core_131 = input_a[21] & input_a[19];
  assign popcount38_wm2a_core_132 = input_a[15] ^ input_a[11];
  assign popcount38_wm2a_core_134 = ~(input_a[31] ^ input_a[5]);
  assign popcount38_wm2a_core_135 = popcount38_wm2a_core_070 ^ popcount38_wm2a_core_118;
  assign popcount38_wm2a_core_137 = ~popcount38_wm2a_core_135;
  assign popcount38_wm2a_core_139 = popcount38_wm2a_core_070 | popcount38_wm2a_core_135;
  assign popcount38_wm2a_core_140 = popcount38_wm2a_core_073 ^ popcount38_wm2a_core_123;
  assign popcount38_wm2a_core_142 = popcount38_wm2a_core_140 ^ popcount38_wm2a_core_139;
  assign popcount38_wm2a_core_143 = ~(input_a[10] ^ input_a[21]);
  assign popcount38_wm2a_core_144 = ~input_a[27];
  assign popcount38_wm2a_core_146 = input_a[9] ^ input_a[14];
  assign popcount38_wm2a_core_150 = input_a[29] & input_a[34];
  assign popcount38_wm2a_core_151 = ~(input_a[18] | input_a[13]);
  assign popcount38_wm2a_core_152 = ~(input_a[5] | input_a[23]);
  assign popcount38_wm2a_core_153 = ~(input_a[27] ^ input_a[0]);
  assign popcount38_wm2a_core_156 = input_a[1] & input_a[12];
  assign popcount38_wm2a_core_157 = ~input_a[0];
  assign popcount38_wm2a_core_160 = input_a[19] & input_a[16];
  assign popcount38_wm2a_core_161 = popcount38_wm2a_core_156 ^ input_a[21];
  assign popcount38_wm2a_core_162 = popcount38_wm2a_core_156 & input_a[21];
  assign popcount38_wm2a_core_163 = popcount38_wm2a_core_161 ^ popcount38_wm2a_core_160;
  assign popcount38_wm2a_core_164 = popcount38_wm2a_core_161 & popcount38_wm2a_core_160;
  assign popcount38_wm2a_core_165 = popcount38_wm2a_core_162 | popcount38_wm2a_core_164;
  assign popcount38_wm2a_core_166 = ~(input_a[7] & input_a[5]);
  assign popcount38_wm2a_core_167 = input_a[4] & input_a[23];
  assign popcount38_wm2a_core_168 = ~input_a[3];
  assign popcount38_wm2a_core_170 = ~(input_a[7] ^ input_a[9]);
  assign popcount38_wm2a_core_171 = input_a[25] & input_a[28];
  assign popcount38_wm2a_core_173 = ~(input_a[23] ^ input_a[33]);
  assign popcount38_wm2a_core_175 = ~(input_a[20] & input_a[6]);
  assign popcount38_wm2a_core_176 = popcount38_wm2a_core_167 | popcount38_wm2a_core_171;
  assign popcount38_wm2a_core_177 = ~input_a[13];
  assign popcount38_wm2a_core_183 = input_a[30] | input_a[37];
  assign popcount38_wm2a_core_184 = ~(input_a[26] | input_a[10]);
  assign popcount38_wm2a_core_185 = popcount38_wm2a_core_163 ^ popcount38_wm2a_core_176;
  assign popcount38_wm2a_core_186 = popcount38_wm2a_core_163 & popcount38_wm2a_core_176;
  assign popcount38_wm2a_core_188 = ~(input_a[36] | input_a[32]);
  assign popcount38_wm2a_core_192 = popcount38_wm2a_core_165 | popcount38_wm2a_core_186;
  assign popcount38_wm2a_core_193 = input_a[27] ^ input_a[2];
  assign popcount38_wm2a_core_194 = ~(input_a[1] | input_a[35]);
  assign popcount38_wm2a_core_196 = ~input_a[23];
  assign popcount38_wm2a_core_198 = input_a[6] ^ input_a[6];
  assign popcount38_wm2a_core_199 = ~(input_a[1] ^ input_a[7]);
  assign popcount38_wm2a_core_200 = ~(input_a[7] ^ input_a[12]);
  assign popcount38_wm2a_core_201 = ~(input_a[8] ^ input_a[24]);
  assign popcount38_wm2a_core_202 = ~(input_a[28] ^ input_a[0]);
  assign popcount38_wm2a_core_203 = ~(input_a[36] & input_a[30]);
  assign popcount38_wm2a_core_205 = input_a[34] & input_a[33];
  assign popcount38_wm2a_core_206 = ~(input_a[13] ^ input_a[13]);
  assign popcount38_wm2a_core_207 = ~(input_a[33] ^ input_a[28]);
  assign popcount38_wm2a_core_211 = ~(input_a[17] ^ input_a[35]);
  assign popcount38_wm2a_core_213 = input_a[35] | input_a[23];
  assign popcount38_wm2a_core_214 = ~(input_a[13] & input_a[15]);
  assign popcount38_wm2a_core_215 = input_a[10] & input_a[29];
  assign popcount38_wm2a_core_216 = input_a[26] | input_a[17];
  assign popcount38_wm2a_core_218 = ~input_a[7];
  assign popcount38_wm2a_core_219 = input_a[31] ^ input_a[12];
  assign popcount38_wm2a_core_220 = input_a[13] | input_a[22];
  assign popcount38_wm2a_core_222 = ~(input_a[29] & input_a[33]);
  assign popcount38_wm2a_core_223 = input_a[27] & input_a[33];
  assign popcount38_wm2a_core_224 = popcount38_wm2a_core_215 ^ popcount38_wm2a_core_220;
  assign popcount38_wm2a_core_225 = popcount38_wm2a_core_215 & popcount38_wm2a_core_220;
  assign popcount38_wm2a_core_226 = popcount38_wm2a_core_224 ^ popcount38_wm2a_core_223;
  assign popcount38_wm2a_core_227 = popcount38_wm2a_core_224 & popcount38_wm2a_core_223;
  assign popcount38_wm2a_core_228 = popcount38_wm2a_core_225 | popcount38_wm2a_core_227;
  assign popcount38_wm2a_core_230 = input_a[2] | input_a[0];
  assign popcount38_wm2a_core_231 = input_a[7] & input_a[15];
  assign popcount38_wm2a_core_232 = input_a[36] & input_a[0];
  assign popcount38_wm2a_core_233_not = ~popcount38_wm2a_core_226;
  assign popcount38_wm2a_core_235 = popcount38_wm2a_core_233_not ^ popcount38_wm2a_core_232;
  assign popcount38_wm2a_core_236 = input_a[0] & input_a[36];
  assign popcount38_wm2a_core_237 = popcount38_wm2a_core_226 | popcount38_wm2a_core_236;
  assign popcount38_wm2a_core_240 = popcount38_wm2a_core_228 ^ popcount38_wm2a_core_237;
  assign popcount38_wm2a_core_241 = popcount38_wm2a_core_228 & popcount38_wm2a_core_237;
  assign popcount38_wm2a_core_246 = input_a[1] ^ input_a[34];
  assign popcount38_wm2a_core_247 = input_a[25] ^ input_a[28];
  assign popcount38_wm2a_core_249 = ~(input_a[25] | input_a[18]);
  assign popcount38_wm2a_core_250 = popcount38_wm2a_core_185 ^ popcount38_wm2a_core_235;
  assign popcount38_wm2a_core_251 = popcount38_wm2a_core_185 & popcount38_wm2a_core_235;
  assign popcount38_wm2a_core_253 = ~input_a[18];
  assign popcount38_wm2a_core_255 = popcount38_wm2a_core_192 ^ popcount38_wm2a_core_240;
  assign popcount38_wm2a_core_256 = popcount38_wm2a_core_192 & popcount38_wm2a_core_240;
  assign popcount38_wm2a_core_257 = popcount38_wm2a_core_255 ^ popcount38_wm2a_core_251;
  assign popcount38_wm2a_core_258 = popcount38_wm2a_core_255 & popcount38_wm2a_core_251;
  assign popcount38_wm2a_core_259 = popcount38_wm2a_core_256 | popcount38_wm2a_core_258;
  assign popcount38_wm2a_core_261 = input_a[7] & input_a[26];
  assign popcount38_wm2a_core_262 = popcount38_wm2a_core_241 | popcount38_wm2a_core_259;
  assign popcount38_wm2a_core_263 = ~(input_a[10] & input_a[30]);
  assign popcount38_wm2a_core_264 = input_a[6] ^ input_a[11];
  assign popcount38_wm2a_core_265 = input_a[2] & input_a[0];
  assign popcount38_wm2a_core_266 = input_a[9] ^ input_a[24];
  assign popcount38_wm2a_core_267 = ~input_a[29];
  assign popcount38_wm2a_core_268 = input_a[28] & input_a[14];
  assign popcount38_wm2a_core_269 = input_a[29] | input_a[9];
  assign popcount38_wm2a_core_270 = input_a[33] | input_a[3];
  assign popcount38_wm2a_core_272 = popcount38_wm2a_core_137 ^ popcount38_wm2a_core_250;
  assign popcount38_wm2a_core_273 = popcount38_wm2a_core_137 & popcount38_wm2a_core_250;
  assign popcount38_wm2a_core_274 = popcount38_wm2a_core_272 ^ popcount38_wm2a_core_183;
  assign popcount38_wm2a_core_275 = popcount38_wm2a_core_272 & popcount38_wm2a_core_183;
  assign popcount38_wm2a_core_276 = popcount38_wm2a_core_273 | popcount38_wm2a_core_275;
  assign popcount38_wm2a_core_277 = popcount38_wm2a_core_142 ^ popcount38_wm2a_core_257;
  assign popcount38_wm2a_core_278 = popcount38_wm2a_core_142 & popcount38_wm2a_core_257;
  assign popcount38_wm2a_core_279 = popcount38_wm2a_core_277 ^ popcount38_wm2a_core_276;
  assign popcount38_wm2a_core_280 = popcount38_wm2a_core_277 & popcount38_wm2a_core_276;
  assign popcount38_wm2a_core_281 = popcount38_wm2a_core_278 | popcount38_wm2a_core_280;
  assign popcount38_wm2a_core_282_not = ~popcount38_wm2a_core_262;
  assign popcount38_wm2a_core_284 = popcount38_wm2a_core_282_not ^ popcount38_wm2a_core_281;
  assign popcount38_wm2a_core_285 = popcount38_wm2a_core_282_not & popcount38_wm2a_core_281;
  assign popcount38_wm2a_core_286 = popcount38_wm2a_core_262 | popcount38_wm2a_core_285;
  assign popcount38_wm2a_core_288 = ~(input_a[27] ^ input_a[10]);
  assign popcount38_wm2a_core_290 = ~(input_a[25] ^ input_a[21]);
  assign popcount38_wm2a_core_291 = input_a[32] | input_a[23];
  assign popcount38_wm2a_core_293 = ~(input_a[22] | input_a[7]);
  assign popcount38_wm2a_core_294 = ~(input_a[9] ^ input_a[5]);
  assign popcount38_wm2a_core_296 = input_a[21] | input_a[9];

  assign popcount38_wm2a_out[0] = popcount38_wm2a_core_087;
  assign popcount38_wm2a_out[1] = popcount38_wm2a_core_274;
  assign popcount38_wm2a_out[2] = popcount38_wm2a_core_279;
  assign popcount38_wm2a_out[3] = popcount38_wm2a_core_284;
  assign popcount38_wm2a_out[4] = popcount38_wm2a_core_286;
  assign popcount38_wm2a_out[5] = 1'b0;
endmodule