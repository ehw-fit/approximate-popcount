// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.05623
// WCE=14.0
// EP=0.963036%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_rr23(input [20:0] input_a, output [4:0] popcount21_rr23_out);
  wire popcount21_rr23_core_023;
  wire popcount21_rr23_core_025;
  wire popcount21_rr23_core_026;
  wire popcount21_rr23_core_027;
  wire popcount21_rr23_core_028;
  wire popcount21_rr23_core_029;
  wire popcount21_rr23_core_031_not;
  wire popcount21_rr23_core_033;
  wire popcount21_rr23_core_034;
  wire popcount21_rr23_core_036;
  wire popcount21_rr23_core_037;
  wire popcount21_rr23_core_041;
  wire popcount21_rr23_core_043;
  wire popcount21_rr23_core_044;
  wire popcount21_rr23_core_046;
  wire popcount21_rr23_core_047;
  wire popcount21_rr23_core_048;
  wire popcount21_rr23_core_051;
  wire popcount21_rr23_core_053;
  wire popcount21_rr23_core_055;
  wire popcount21_rr23_core_056;
  wire popcount21_rr23_core_057;
  wire popcount21_rr23_core_058;
  wire popcount21_rr23_core_059;
  wire popcount21_rr23_core_060;
  wire popcount21_rr23_core_062;
  wire popcount21_rr23_core_063;
  wire popcount21_rr23_core_065_not;
  wire popcount21_rr23_core_067;
  wire popcount21_rr23_core_068;
  wire popcount21_rr23_core_069;
  wire popcount21_rr23_core_070;
  wire popcount21_rr23_core_071;
  wire popcount21_rr23_core_072;
  wire popcount21_rr23_core_074;
  wire popcount21_rr23_core_075;
  wire popcount21_rr23_core_076;
  wire popcount21_rr23_core_078;
  wire popcount21_rr23_core_079;
  wire popcount21_rr23_core_080;
  wire popcount21_rr23_core_083;
  wire popcount21_rr23_core_084;
  wire popcount21_rr23_core_085;
  wire popcount21_rr23_core_088;
  wire popcount21_rr23_core_090;
  wire popcount21_rr23_core_091;
  wire popcount21_rr23_core_092;
  wire popcount21_rr23_core_093;
  wire popcount21_rr23_core_094;
  wire popcount21_rr23_core_095;
  wire popcount21_rr23_core_097;
  wire popcount21_rr23_core_102;
  wire popcount21_rr23_core_103;
  wire popcount21_rr23_core_104;
  wire popcount21_rr23_core_105;
  wire popcount21_rr23_core_106;
  wire popcount21_rr23_core_108;
  wire popcount21_rr23_core_109;
  wire popcount21_rr23_core_111;
  wire popcount21_rr23_core_112;
  wire popcount21_rr23_core_113;
  wire popcount21_rr23_core_114;
  wire popcount21_rr23_core_116;
  wire popcount21_rr23_core_118;
  wire popcount21_rr23_core_119;
  wire popcount21_rr23_core_121;
  wire popcount21_rr23_core_123_not;
  wire popcount21_rr23_core_125;
  wire popcount21_rr23_core_127;
  wire popcount21_rr23_core_128_not;
  wire popcount21_rr23_core_129;
  wire popcount21_rr23_core_130;
  wire popcount21_rr23_core_131;
  wire popcount21_rr23_core_132;
  wire popcount21_rr23_core_134;
  wire popcount21_rr23_core_136;
  wire popcount21_rr23_core_137;
  wire popcount21_rr23_core_139;
  wire popcount21_rr23_core_142;
  wire popcount21_rr23_core_144;
  wire popcount21_rr23_core_146;
  wire popcount21_rr23_core_148;
  wire popcount21_rr23_core_149;
  wire popcount21_rr23_core_150;
  wire popcount21_rr23_core_151;
  wire popcount21_rr23_core_152;

  assign popcount21_rr23_core_023 = ~(input_a[18] & input_a[7]);
  assign popcount21_rr23_core_025 = ~input_a[16];
  assign popcount21_rr23_core_026 = input_a[13] | input_a[7];
  assign popcount21_rr23_core_027 = ~(input_a[9] ^ input_a[9]);
  assign popcount21_rr23_core_028 = ~(input_a[13] | input_a[15]);
  assign popcount21_rr23_core_029 = input_a[18] | input_a[4];
  assign popcount21_rr23_core_031_not = ~input_a[14];
  assign popcount21_rr23_core_033 = input_a[15] ^ input_a[2];
  assign popcount21_rr23_core_034 = ~(input_a[12] ^ input_a[5]);
  assign popcount21_rr23_core_036 = input_a[5] & input_a[14];
  assign popcount21_rr23_core_037 = ~input_a[9];
  assign popcount21_rr23_core_041 = ~(input_a[12] | input_a[6]);
  assign popcount21_rr23_core_043 = input_a[17] | input_a[14];
  assign popcount21_rr23_core_044 = input_a[8] & input_a[7];
  assign popcount21_rr23_core_046 = ~(input_a[17] ^ input_a[3]);
  assign popcount21_rr23_core_047 = input_a[16] | input_a[18];
  assign popcount21_rr23_core_048 = input_a[7] | input_a[4];
  assign popcount21_rr23_core_051 = ~(input_a[2] & input_a[2]);
  assign popcount21_rr23_core_053 = ~(input_a[2] & input_a[4]);
  assign popcount21_rr23_core_055 = input_a[11] | input_a[15];
  assign popcount21_rr23_core_056 = input_a[11] | input_a[10];
  assign popcount21_rr23_core_057 = input_a[9] & input_a[6];
  assign popcount21_rr23_core_058 = input_a[8] ^ input_a[19];
  assign popcount21_rr23_core_059 = input_a[12] | input_a[11];
  assign popcount21_rr23_core_060 = ~(input_a[17] ^ input_a[2]);
  assign popcount21_rr23_core_062 = ~(input_a[8] | input_a[5]);
  assign popcount21_rr23_core_063 = input_a[2] & input_a[14];
  assign popcount21_rr23_core_065_not = ~input_a[7];
  assign popcount21_rr23_core_067 = ~(input_a[11] ^ input_a[8]);
  assign popcount21_rr23_core_068 = ~(input_a[19] ^ input_a[6]);
  assign popcount21_rr23_core_069 = ~(input_a[1] | input_a[12]);
  assign popcount21_rr23_core_070 = input_a[12] & input_a[7];
  assign popcount21_rr23_core_071 = input_a[17] ^ input_a[7];
  assign popcount21_rr23_core_072 = ~(input_a[4] | input_a[14]);
  assign popcount21_rr23_core_074 = ~(input_a[1] & input_a[1]);
  assign popcount21_rr23_core_075 = input_a[19] & input_a[16];
  assign popcount21_rr23_core_076 = ~input_a[0];
  assign popcount21_rr23_core_078 = ~(input_a[10] & input_a[12]);
  assign popcount21_rr23_core_079 = input_a[5] | input_a[4];
  assign popcount21_rr23_core_080 = ~input_a[5];
  assign popcount21_rr23_core_083 = ~(input_a[18] & input_a[15]);
  assign popcount21_rr23_core_084 = ~(input_a[1] & input_a[17]);
  assign popcount21_rr23_core_085 = input_a[17] | input_a[11];
  assign popcount21_rr23_core_088 = ~(input_a[1] & input_a[17]);
  assign popcount21_rr23_core_090 = input_a[7] | input_a[3];
  assign popcount21_rr23_core_091 = input_a[11] ^ input_a[2];
  assign popcount21_rr23_core_092 = ~input_a[3];
  assign popcount21_rr23_core_093 = ~(input_a[7] & input_a[18]);
  assign popcount21_rr23_core_094 = input_a[11] ^ input_a[3];
  assign popcount21_rr23_core_095 = ~(input_a[12] ^ input_a[19]);
  assign popcount21_rr23_core_097 = input_a[10] ^ input_a[9];
  assign popcount21_rr23_core_102 = input_a[17] | input_a[10];
  assign popcount21_rr23_core_103 = input_a[3] | input_a[1];
  assign popcount21_rr23_core_104 = input_a[6] & input_a[4];
  assign popcount21_rr23_core_105 = ~input_a[3];
  assign popcount21_rr23_core_106 = input_a[11] & input_a[0];
  assign popcount21_rr23_core_108 = ~input_a[15];
  assign popcount21_rr23_core_109 = ~(input_a[11] | input_a[19]);
  assign popcount21_rr23_core_111 = input_a[5] & input_a[17];
  assign popcount21_rr23_core_112 = ~(input_a[19] & input_a[10]);
  assign popcount21_rr23_core_113 = input_a[9] ^ input_a[12];
  assign popcount21_rr23_core_114 = ~(input_a[13] & input_a[15]);
  assign popcount21_rr23_core_116 = ~(input_a[17] | input_a[5]);
  assign popcount21_rr23_core_118 = ~input_a[11];
  assign popcount21_rr23_core_119 = input_a[7] ^ input_a[19];
  assign popcount21_rr23_core_121 = input_a[10] | input_a[20];
  assign popcount21_rr23_core_123_not = ~input_a[2];
  assign popcount21_rr23_core_125 = ~(input_a[12] | input_a[18]);
  assign popcount21_rr23_core_127 = ~(input_a[7] ^ input_a[11]);
  assign popcount21_rr23_core_128_not = ~input_a[10];
  assign popcount21_rr23_core_129 = ~input_a[16];
  assign popcount21_rr23_core_130 = ~(input_a[8] & input_a[4]);
  assign popcount21_rr23_core_131 = ~(input_a[16] | input_a[18]);
  assign popcount21_rr23_core_132 = input_a[3] | input_a[1];
  assign popcount21_rr23_core_134 = input_a[8] ^ input_a[15];
  assign popcount21_rr23_core_136 = input_a[20] | input_a[20];
  assign popcount21_rr23_core_137 = ~(input_a[4] & input_a[5]);
  assign popcount21_rr23_core_139 = ~(input_a[0] | input_a[17]);
  assign popcount21_rr23_core_142 = ~(input_a[15] & input_a[16]);
  assign popcount21_rr23_core_144 = ~(input_a[12] ^ input_a[15]);
  assign popcount21_rr23_core_146 = ~(input_a[5] ^ input_a[17]);
  assign popcount21_rr23_core_148 = ~input_a[10];
  assign popcount21_rr23_core_149 = input_a[7] & input_a[12];
  assign popcount21_rr23_core_150 = input_a[20] ^ input_a[19];
  assign popcount21_rr23_core_151 = ~(input_a[4] | input_a[16]);
  assign popcount21_rr23_core_152 = input_a[18] ^ input_a[4];

  assign popcount21_rr23_out[0] = input_a[18];
  assign popcount21_rr23_out[1] = 1'b1;
  assign popcount21_rr23_out[2] = 1'b1;
  assign popcount21_rr23_out[3] = 1'b0;
  assign popcount21_rr23_out[4] = 1'b0;
endmodule