// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.40814
// WCE=5.0
// EP=0.787842%
// Printed PDK parameters:
//  Area=41955420.0
//  Delay=57655176.0
//  Power=1703600.0

module popcount21_6w8j(input [20:0] input_a, output [4:0] popcount21_6w8j_out);
  wire popcount21_6w8j_core_023;
  wire popcount21_6w8j_core_024;
  wire popcount21_6w8j_core_025;
  wire popcount21_6w8j_core_026;
  wire popcount21_6w8j_core_027;
  wire popcount21_6w8j_core_028;
  wire popcount21_6w8j_core_029;
  wire popcount21_6w8j_core_031;
  wire popcount21_6w8j_core_032;
  wire popcount21_6w8j_core_033;
  wire popcount21_6w8j_core_034;
  wire popcount21_6w8j_core_035;
  wire popcount21_6w8j_core_036;
  wire popcount21_6w8j_core_037;
  wire popcount21_6w8j_core_039_not;
  wire popcount21_6w8j_core_040;
  wire popcount21_6w8j_core_041;
  wire popcount21_6w8j_core_042;
  wire popcount21_6w8j_core_043;
  wire popcount21_6w8j_core_044;
  wire popcount21_6w8j_core_045;
  wire popcount21_6w8j_core_046;
  wire popcount21_6w8j_core_049;
  wire popcount21_6w8j_core_050;
  wire popcount21_6w8j_core_051;
  wire popcount21_6w8j_core_052;
  wire popcount21_6w8j_core_053;
  wire popcount21_6w8j_core_054;
  wire popcount21_6w8j_core_058;
  wire popcount21_6w8j_core_059;
  wire popcount21_6w8j_core_060;
  wire popcount21_6w8j_core_062;
  wire popcount21_6w8j_core_064;
  wire popcount21_6w8j_core_065;
  wire popcount21_6w8j_core_066;
  wire popcount21_6w8j_core_067;
  wire popcount21_6w8j_core_073;
  wire popcount21_6w8j_core_074;
  wire popcount21_6w8j_core_075;
  wire popcount21_6w8j_core_077;
  wire popcount21_6w8j_core_078;
  wire popcount21_6w8j_core_079;
  wire popcount21_6w8j_core_080;
  wire popcount21_6w8j_core_081;
  wire popcount21_6w8j_core_082;
  wire popcount21_6w8j_core_083;
  wire popcount21_6w8j_core_084;
  wire popcount21_6w8j_core_085;
  wire popcount21_6w8j_core_086;
  wire popcount21_6w8j_core_087;
  wire popcount21_6w8j_core_088;
  wire popcount21_6w8j_core_089;
  wire popcount21_6w8j_core_090;
  wire popcount21_6w8j_core_092;
  wire popcount21_6w8j_core_093;
  wire popcount21_6w8j_core_097;
  wire popcount21_6w8j_core_099;
  wire popcount21_6w8j_core_100;
  wire popcount21_6w8j_core_101;
  wire popcount21_6w8j_core_103;
  wire popcount21_6w8j_core_104;
  wire popcount21_6w8j_core_105;
  wire popcount21_6w8j_core_106;
  wire popcount21_6w8j_core_107;
  wire popcount21_6w8j_core_108;
  wire popcount21_6w8j_core_109;
  wire popcount21_6w8j_core_111;
  wire popcount21_6w8j_core_113;
  wire popcount21_6w8j_core_114;
  wire popcount21_6w8j_core_116;
  wire popcount21_6w8j_core_117;
  wire popcount21_6w8j_core_118;
  wire popcount21_6w8j_core_119;
  wire popcount21_6w8j_core_120;
  wire popcount21_6w8j_core_121;
  wire popcount21_6w8j_core_122;
  wire popcount21_6w8j_core_123;
  wire popcount21_6w8j_core_124;
  wire popcount21_6w8j_core_125;
  wire popcount21_6w8j_core_126;
  wire popcount21_6w8j_core_128;
  wire popcount21_6w8j_core_130;
  wire popcount21_6w8j_core_134_not;
  wire popcount21_6w8j_core_136;
  wire popcount21_6w8j_core_139;
  wire popcount21_6w8j_core_140;
  wire popcount21_6w8j_core_141;
  wire popcount21_6w8j_core_142;
  wire popcount21_6w8j_core_143;
  wire popcount21_6w8j_core_144;
  wire popcount21_6w8j_core_145;
  wire popcount21_6w8j_core_146;
  wire popcount21_6w8j_core_147;
  wire popcount21_6w8j_core_148;
  wire popcount21_6w8j_core_149;
  wire popcount21_6w8j_core_150;
  wire popcount21_6w8j_core_152;

  assign popcount21_6w8j_core_023 = input_a[0] ^ input_a[1];
  assign popcount21_6w8j_core_024 = input_a[0] & input_a[1];
  assign popcount21_6w8j_core_025 = input_a[3] ^ input_a[4];
  assign popcount21_6w8j_core_026 = input_a[3] & input_a[4];
  assign popcount21_6w8j_core_027 = input_a[2] ^ popcount21_6w8j_core_025;
  assign popcount21_6w8j_core_028 = input_a[2] & popcount21_6w8j_core_025;
  assign popcount21_6w8j_core_029 = popcount21_6w8j_core_026 | popcount21_6w8j_core_028;
  assign popcount21_6w8j_core_031 = ~input_a[2];
  assign popcount21_6w8j_core_032 = popcount21_6w8j_core_023 & popcount21_6w8j_core_027;
  assign popcount21_6w8j_core_033 = popcount21_6w8j_core_024 ^ popcount21_6w8j_core_029;
  assign popcount21_6w8j_core_034 = popcount21_6w8j_core_024 & popcount21_6w8j_core_029;
  assign popcount21_6w8j_core_035 = popcount21_6w8j_core_033 ^ popcount21_6w8j_core_032;
  assign popcount21_6w8j_core_036 = popcount21_6w8j_core_033 & popcount21_6w8j_core_032;
  assign popcount21_6w8j_core_037 = popcount21_6w8j_core_034 | popcount21_6w8j_core_036;
  assign popcount21_6w8j_core_039_not = ~input_a[6];
  assign popcount21_6w8j_core_040 = input_a[11] & input_a[15];
  assign popcount21_6w8j_core_041 = input_a[5] & input_a[6];
  assign popcount21_6w8j_core_042 = input_a[8] | input_a[9];
  assign popcount21_6w8j_core_043 = input_a[8] & input_a[9];
  assign popcount21_6w8j_core_044 = input_a[18] & input_a[20];
  assign popcount21_6w8j_core_045 = input_a[7] & popcount21_6w8j_core_042;
  assign popcount21_6w8j_core_046 = popcount21_6w8j_core_043 | popcount21_6w8j_core_045;
  assign popcount21_6w8j_core_049 = input_a[19] & input_a[15];
  assign popcount21_6w8j_core_050 = popcount21_6w8j_core_041 | popcount21_6w8j_core_046;
  assign popcount21_6w8j_core_051 = popcount21_6w8j_core_041 & popcount21_6w8j_core_046;
  assign popcount21_6w8j_core_052 = popcount21_6w8j_core_050 | popcount21_6w8j_core_049;
  assign popcount21_6w8j_core_053 = popcount21_6w8j_core_050 & popcount21_6w8j_core_049;
  assign popcount21_6w8j_core_054 = popcount21_6w8j_core_051 | popcount21_6w8j_core_053;
  assign popcount21_6w8j_core_058 = ~(input_a[7] | input_a[19]);
  assign popcount21_6w8j_core_059 = input_a[14] ^ input_a[6];
  assign popcount21_6w8j_core_060 = popcount21_6w8j_core_035 & popcount21_6w8j_core_052;
  assign popcount21_6w8j_core_062 = input_a[3] ^ input_a[6];
  assign popcount21_6w8j_core_064 = popcount21_6w8j_core_037 ^ popcount21_6w8j_core_054;
  assign popcount21_6w8j_core_065 = popcount21_6w8j_core_037 & popcount21_6w8j_core_054;
  assign popcount21_6w8j_core_066 = popcount21_6w8j_core_064 | popcount21_6w8j_core_060;
  assign popcount21_6w8j_core_067 = ~(input_a[15] ^ input_a[2]);
  assign popcount21_6w8j_core_073 = ~(input_a[20] ^ input_a[9]);
  assign popcount21_6w8j_core_074 = input_a[10] ^ input_a[11];
  assign popcount21_6w8j_core_075 = input_a[10] & input_a[11];
  assign popcount21_6w8j_core_077 = input_a[13] & input_a[14];
  assign popcount21_6w8j_core_078 = ~input_a[12];
  assign popcount21_6w8j_core_079 = input_a[14] ^ input_a[13];
  assign popcount21_6w8j_core_080 = popcount21_6w8j_core_077 ^ input_a[12];
  assign popcount21_6w8j_core_081 = popcount21_6w8j_core_077 & input_a[12];
  assign popcount21_6w8j_core_082 = popcount21_6w8j_core_074 ^ popcount21_6w8j_core_078;
  assign popcount21_6w8j_core_083 = popcount21_6w8j_core_074 & popcount21_6w8j_core_078;
  assign popcount21_6w8j_core_084 = popcount21_6w8j_core_075 ^ popcount21_6w8j_core_080;
  assign popcount21_6w8j_core_085 = popcount21_6w8j_core_075 & popcount21_6w8j_core_080;
  assign popcount21_6w8j_core_086 = popcount21_6w8j_core_084 ^ popcount21_6w8j_core_083;
  assign popcount21_6w8j_core_087 = popcount21_6w8j_core_084 & popcount21_6w8j_core_083;
  assign popcount21_6w8j_core_088 = popcount21_6w8j_core_085 | popcount21_6w8j_core_087;
  assign popcount21_6w8j_core_089 = popcount21_6w8j_core_081 | popcount21_6w8j_core_088;
  assign popcount21_6w8j_core_090 = ~(input_a[11] & input_a[12]);
  assign popcount21_6w8j_core_092 = ~input_a[7];
  assign popcount21_6w8j_core_093 = input_a[17] | input_a[16];
  assign popcount21_6w8j_core_097 = input_a[16] | input_a[20];
  assign popcount21_6w8j_core_099 = input_a[18] ^ popcount21_6w8j_core_097;
  assign popcount21_6w8j_core_100 = input_a[8] ^ input_a[6];
  assign popcount21_6w8j_core_101 = input_a[20] | input_a[16];
  assign popcount21_6w8j_core_103 = input_a[17] ^ popcount21_6w8j_core_099;
  assign popcount21_6w8j_core_104 = input_a[17] & popcount21_6w8j_core_099;
  assign popcount21_6w8j_core_105 = ~input_a[18];
  assign popcount21_6w8j_core_106 = input_a[18] & popcount21_6w8j_core_101;
  assign popcount21_6w8j_core_107 = popcount21_6w8j_core_105 ^ popcount21_6w8j_core_104;
  assign popcount21_6w8j_core_108 = popcount21_6w8j_core_105 & popcount21_6w8j_core_104;
  assign popcount21_6w8j_core_109 = popcount21_6w8j_core_106 | popcount21_6w8j_core_108;
  assign popcount21_6w8j_core_111 = ~(input_a[9] & input_a[17]);
  assign popcount21_6w8j_core_113 = ~input_a[9];
  assign popcount21_6w8j_core_114 = input_a[16] ^ input_a[14];
  assign popcount21_6w8j_core_116 = popcount21_6w8j_core_082 & popcount21_6w8j_core_103;
  assign popcount21_6w8j_core_117 = popcount21_6w8j_core_086 ^ popcount21_6w8j_core_107;
  assign popcount21_6w8j_core_118 = popcount21_6w8j_core_086 & popcount21_6w8j_core_107;
  assign popcount21_6w8j_core_119 = popcount21_6w8j_core_117 ^ popcount21_6w8j_core_116;
  assign popcount21_6w8j_core_120 = popcount21_6w8j_core_117 & popcount21_6w8j_core_116;
  assign popcount21_6w8j_core_121 = popcount21_6w8j_core_118 | popcount21_6w8j_core_120;
  assign popcount21_6w8j_core_122 = popcount21_6w8j_core_089 ^ popcount21_6w8j_core_109;
  assign popcount21_6w8j_core_123 = popcount21_6w8j_core_089 & popcount21_6w8j_core_109;
  assign popcount21_6w8j_core_124 = popcount21_6w8j_core_122 ^ popcount21_6w8j_core_121;
  assign popcount21_6w8j_core_125 = popcount21_6w8j_core_122 & popcount21_6w8j_core_121;
  assign popcount21_6w8j_core_126 = popcount21_6w8j_core_123 | popcount21_6w8j_core_125;
  assign popcount21_6w8j_core_128 = ~(input_a[19] | input_a[5]);
  assign popcount21_6w8j_core_130 = input_a[18] | input_a[0];
  assign popcount21_6w8j_core_134_not = ~popcount21_6w8j_core_119;
  assign popcount21_6w8j_core_136 = ~(input_a[1] | input_a[9]);
  assign popcount21_6w8j_core_139 = popcount21_6w8j_core_066 ^ popcount21_6w8j_core_124;
  assign popcount21_6w8j_core_140 = popcount21_6w8j_core_066 & popcount21_6w8j_core_124;
  assign popcount21_6w8j_core_141 = popcount21_6w8j_core_139 ^ popcount21_6w8j_core_119;
  assign popcount21_6w8j_core_142 = popcount21_6w8j_core_139 & popcount21_6w8j_core_119;
  assign popcount21_6w8j_core_143 = popcount21_6w8j_core_140 | popcount21_6w8j_core_142;
  assign popcount21_6w8j_core_144 = popcount21_6w8j_core_065 ^ popcount21_6w8j_core_126;
  assign popcount21_6w8j_core_145 = popcount21_6w8j_core_065 & popcount21_6w8j_core_126;
  assign popcount21_6w8j_core_146 = popcount21_6w8j_core_144 ^ popcount21_6w8j_core_143;
  assign popcount21_6w8j_core_147 = popcount21_6w8j_core_144 & popcount21_6w8j_core_143;
  assign popcount21_6w8j_core_148 = popcount21_6w8j_core_145 | popcount21_6w8j_core_147;
  assign popcount21_6w8j_core_149 = ~(input_a[19] ^ input_a[1]);
  assign popcount21_6w8j_core_150 = ~(input_a[20] & input_a[6]);
  assign popcount21_6w8j_core_152 = input_a[7] ^ input_a[7];

  assign popcount21_6w8j_out[0] = 1'b0;
  assign popcount21_6w8j_out[1] = popcount21_6w8j_core_134_not;
  assign popcount21_6w8j_out[2] = popcount21_6w8j_core_141;
  assign popcount21_6w8j_out[3] = popcount21_6w8j_core_146;
  assign popcount21_6w8j_out[4] = popcount21_6w8j_core_148;
endmodule