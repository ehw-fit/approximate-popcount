// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.61026
// WCE=8.0
// EP=0.808505%
// Printed PDK parameters:
//  Area=63639387.0
//  Delay=79895880.0
//  Power=3553900.0

module popcount38_j2g7(input [37:0] input_a, output [5:0] popcount38_j2g7_out);
  wire popcount38_j2g7_core_040;
  wire popcount38_j2g7_core_042;
  wire popcount38_j2g7_core_043;
  wire popcount38_j2g7_core_047;
  wire popcount38_j2g7_core_051;
  wire popcount38_j2g7_core_053;
  wire popcount38_j2g7_core_054;
  wire popcount38_j2g7_core_055;
  wire popcount38_j2g7_core_056;
  wire popcount38_j2g7_core_058;
  wire popcount38_j2g7_core_059;
  wire popcount38_j2g7_core_060;
  wire popcount38_j2g7_core_061;
  wire popcount38_j2g7_core_062;
  wire popcount38_j2g7_core_065;
  wire popcount38_j2g7_core_068;
  wire popcount38_j2g7_core_069;
  wire popcount38_j2g7_core_073;
  wire popcount38_j2g7_core_075;
  wire popcount38_j2g7_core_078;
  wire popcount38_j2g7_core_079;
  wire popcount38_j2g7_core_080_not;
  wire popcount38_j2g7_core_081;
  wire popcount38_j2g7_core_082;
  wire popcount38_j2g7_core_083;
  wire popcount38_j2g7_core_087;
  wire popcount38_j2g7_core_090;
  wire popcount38_j2g7_core_091;
  wire popcount38_j2g7_core_093;
  wire popcount38_j2g7_core_094;
  wire popcount38_j2g7_core_095;
  wire popcount38_j2g7_core_096;
  wire popcount38_j2g7_core_097;
  wire popcount38_j2g7_core_098;
  wire popcount38_j2g7_core_103;
  wire popcount38_j2g7_core_105;
  wire popcount38_j2g7_core_107;
  wire popcount38_j2g7_core_108;
  wire popcount38_j2g7_core_109;
  wire popcount38_j2g7_core_110;
  wire popcount38_j2g7_core_111;
  wire popcount38_j2g7_core_112;
  wire popcount38_j2g7_core_113;
  wire popcount38_j2g7_core_114;
  wire popcount38_j2g7_core_116;
  wire popcount38_j2g7_core_117;
  wire popcount38_j2g7_core_120;
  wire popcount38_j2g7_core_121;
  wire popcount38_j2g7_core_124;
  wire popcount38_j2g7_core_126;
  wire popcount38_j2g7_core_127;
  wire popcount38_j2g7_core_129;
  wire popcount38_j2g7_core_130;
  wire popcount38_j2g7_core_131;
  wire popcount38_j2g7_core_133;
  wire popcount38_j2g7_core_134;
  wire popcount38_j2g7_core_135;
  wire popcount38_j2g7_core_136;
  wire popcount38_j2g7_core_137;
  wire popcount38_j2g7_core_138;
  wire popcount38_j2g7_core_139;
  wire popcount38_j2g7_core_142;
  wire popcount38_j2g7_core_143;
  wire popcount38_j2g7_core_144;
  wire popcount38_j2g7_core_146;
  wire popcount38_j2g7_core_148;
  wire popcount38_j2g7_core_149;
  wire popcount38_j2g7_core_150;
  wire popcount38_j2g7_core_156;
  wire popcount38_j2g7_core_157;
  wire popcount38_j2g7_core_158;
  wire popcount38_j2g7_core_159;
  wire popcount38_j2g7_core_160;
  wire popcount38_j2g7_core_161;
  wire popcount38_j2g7_core_162;
  wire popcount38_j2g7_core_163;
  wire popcount38_j2g7_core_164;
  wire popcount38_j2g7_core_166;
  wire popcount38_j2g7_core_167;
  wire popcount38_j2g7_core_169;
  wire popcount38_j2g7_core_171;
  wire popcount38_j2g7_core_172;
  wire popcount38_j2g7_core_173;
  wire popcount38_j2g7_core_175;
  wire popcount38_j2g7_core_176;
  wire popcount38_j2g7_core_177;
  wire popcount38_j2g7_core_181;
  wire popcount38_j2g7_core_183;
  wire popcount38_j2g7_core_184;
  wire popcount38_j2g7_core_185;
  wire popcount38_j2g7_core_186;
  wire popcount38_j2g7_core_187;
  wire popcount38_j2g7_core_188;
  wire popcount38_j2g7_core_189;
  wire popcount38_j2g7_core_190;
  wire popcount38_j2g7_core_191;
  wire popcount38_j2g7_core_192;
  wire popcount38_j2g7_core_193;
  wire popcount38_j2g7_core_194;
  wire popcount38_j2g7_core_197;
  wire popcount38_j2g7_core_198;
  wire popcount38_j2g7_core_199_not;
  wire popcount38_j2g7_core_200;
  wire popcount38_j2g7_core_201_not;
  wire popcount38_j2g7_core_202;
  wire popcount38_j2g7_core_203;
  wire popcount38_j2g7_core_205;
  wire popcount38_j2g7_core_206;
  wire popcount38_j2g7_core_207;
  wire popcount38_j2g7_core_208;
  wire popcount38_j2g7_core_214;
  wire popcount38_j2g7_core_215;
  wire popcount38_j2g7_core_217;
  wire popcount38_j2g7_core_218;
  wire popcount38_j2g7_core_219;
  wire popcount38_j2g7_core_220;
  wire popcount38_j2g7_core_223;
  wire popcount38_j2g7_core_224;
  wire popcount38_j2g7_core_225;
  wire popcount38_j2g7_core_226;
  wire popcount38_j2g7_core_227;
  wire popcount38_j2g7_core_228;
  wire popcount38_j2g7_core_230;
  wire popcount38_j2g7_core_233;
  wire popcount38_j2g7_core_234;
  wire popcount38_j2g7_core_238;
  wire popcount38_j2g7_core_239;
  wire popcount38_j2g7_core_240;
  wire popcount38_j2g7_core_241;
  wire popcount38_j2g7_core_242;
  wire popcount38_j2g7_core_244;
  wire popcount38_j2g7_core_246;
  wire popcount38_j2g7_core_247;
  wire popcount38_j2g7_core_248;
  wire popcount38_j2g7_core_249;
  wire popcount38_j2g7_core_250;
  wire popcount38_j2g7_core_251;
  wire popcount38_j2g7_core_252;
  wire popcount38_j2g7_core_253;
  wire popcount38_j2g7_core_254;
  wire popcount38_j2g7_core_255;
  wire popcount38_j2g7_core_256;
  wire popcount38_j2g7_core_257;
  wire popcount38_j2g7_core_258;
  wire popcount38_j2g7_core_259;
  wire popcount38_j2g7_core_260;
  wire popcount38_j2g7_core_261;
  wire popcount38_j2g7_core_262;
  wire popcount38_j2g7_core_263;
  wire popcount38_j2g7_core_264;
  wire popcount38_j2g7_core_266;
  wire popcount38_j2g7_core_268;
  wire popcount38_j2g7_core_271;
  wire popcount38_j2g7_core_272;
  wire popcount38_j2g7_core_273;
  wire popcount38_j2g7_core_274;
  wire popcount38_j2g7_core_275;
  wire popcount38_j2g7_core_276;
  wire popcount38_j2g7_core_277;
  wire popcount38_j2g7_core_278;
  wire popcount38_j2g7_core_279;
  wire popcount38_j2g7_core_280;
  wire popcount38_j2g7_core_281;
  wire popcount38_j2g7_core_282_not;
  wire popcount38_j2g7_core_284;
  wire popcount38_j2g7_core_285;
  wire popcount38_j2g7_core_286;
  wire popcount38_j2g7_core_289;
  wire popcount38_j2g7_core_290;
  wire popcount38_j2g7_core_292;
  wire popcount38_j2g7_core_293;
  wire popcount38_j2g7_core_296;

  assign popcount38_j2g7_core_040 = input_a[15] | input_a[30];
  assign popcount38_j2g7_core_042 = input_a[22] & input_a[31];
  assign popcount38_j2g7_core_043 = input_a[27] & input_a[22];
  assign popcount38_j2g7_core_047 = ~(input_a[11] ^ input_a[18]);
  assign popcount38_j2g7_core_051 = ~(input_a[5] & input_a[7]);
  assign popcount38_j2g7_core_053 = ~(input_a[28] & input_a[9]);
  assign popcount38_j2g7_core_054 = ~(input_a[16] & input_a[27]);
  assign popcount38_j2g7_core_055 = ~input_a[23];
  assign popcount38_j2g7_core_056 = ~input_a[33];
  assign popcount38_j2g7_core_058 = ~(input_a[0] | input_a[4]);
  assign popcount38_j2g7_core_059 = ~(input_a[31] ^ input_a[7]);
  assign popcount38_j2g7_core_060 = ~input_a[37];
  assign popcount38_j2g7_core_061 = input_a[8] | input_a[18];
  assign popcount38_j2g7_core_062 = input_a[8] & input_a[3];
  assign popcount38_j2g7_core_065 = ~(input_a[6] & input_a[3]);
  assign popcount38_j2g7_core_068 = input_a[22] | input_a[33];
  assign popcount38_j2g7_core_069 = input_a[17] ^ input_a[6];
  assign popcount38_j2g7_core_073 = ~input_a[35];
  assign popcount38_j2g7_core_075 = input_a[30] | input_a[4];
  assign popcount38_j2g7_core_078 = ~(input_a[31] & input_a[11]);
  assign popcount38_j2g7_core_079 = input_a[15] | input_a[12];
  assign popcount38_j2g7_core_080_not = ~input_a[5];
  assign popcount38_j2g7_core_081 = input_a[16] | input_a[21];
  assign popcount38_j2g7_core_082 = input_a[9] ^ input_a[10];
  assign popcount38_j2g7_core_083 = input_a[9] & input_a[10];
  assign popcount38_j2g7_core_087 = input_a[15] ^ input_a[21];
  assign popcount38_j2g7_core_090 = popcount38_j2g7_core_082 ^ input_a[24];
  assign popcount38_j2g7_core_091 = popcount38_j2g7_core_082 & input_a[24];
  assign popcount38_j2g7_core_093 = input_a[33] & input_a[18];
  assign popcount38_j2g7_core_094 = popcount38_j2g7_core_083 | popcount38_j2g7_core_091;
  assign popcount38_j2g7_core_095 = input_a[27] | input_a[29];
  assign popcount38_j2g7_core_096 = ~(input_a[31] & input_a[16]);
  assign popcount38_j2g7_core_097 = input_a[33] ^ input_a[2];
  assign popcount38_j2g7_core_098 = ~input_a[28];
  assign popcount38_j2g7_core_103 = input_a[0] | input_a[17];
  assign popcount38_j2g7_core_105 = input_a[34] ^ input_a[5];
  assign popcount38_j2g7_core_107 = ~(input_a[32] ^ input_a[5]);
  assign popcount38_j2g7_core_108 = ~input_a[2];
  assign popcount38_j2g7_core_109 = input_a[20] ^ input_a[12];
  assign popcount38_j2g7_core_110 = ~(input_a[35] & input_a[35]);
  assign popcount38_j2g7_core_111 = input_a[2] ^ input_a[29];
  assign popcount38_j2g7_core_112 = ~input_a[15];
  assign popcount38_j2g7_core_113 = input_a[22] & input_a[9];
  assign popcount38_j2g7_core_114 = input_a[6] & input_a[2];
  assign popcount38_j2g7_core_116 = popcount38_j2g7_core_090 ^ input_a[3];
  assign popcount38_j2g7_core_117 = popcount38_j2g7_core_090 & input_a[3];
  assign popcount38_j2g7_core_120 = popcount38_j2g7_core_094 ^ popcount38_j2g7_core_117;
  assign popcount38_j2g7_core_121 = popcount38_j2g7_core_094 & popcount38_j2g7_core_117;
  assign popcount38_j2g7_core_124 = input_a[1] | input_a[24];
  assign popcount38_j2g7_core_126 = input_a[23] ^ input_a[22];
  assign popcount38_j2g7_core_127 = ~(input_a[27] & input_a[25]);
  assign popcount38_j2g7_core_129 = ~(input_a[1] | input_a[27]);
  assign popcount38_j2g7_core_130 = input_a[36] & input_a[20];
  assign popcount38_j2g7_core_131 = ~input_a[12];
  assign popcount38_j2g7_core_133 = input_a[12] ^ popcount38_j2g7_core_116;
  assign popcount38_j2g7_core_134 = input_a[12] & popcount38_j2g7_core_116;
  assign popcount38_j2g7_core_135 = popcount38_j2g7_core_043 ^ popcount38_j2g7_core_120;
  assign popcount38_j2g7_core_136 = popcount38_j2g7_core_043 & popcount38_j2g7_core_120;
  assign popcount38_j2g7_core_137 = popcount38_j2g7_core_135 ^ popcount38_j2g7_core_134;
  assign popcount38_j2g7_core_138 = popcount38_j2g7_core_135 & popcount38_j2g7_core_134;
  assign popcount38_j2g7_core_139 = popcount38_j2g7_core_136 | popcount38_j2g7_core_138;
  assign popcount38_j2g7_core_142 = popcount38_j2g7_core_121 | popcount38_j2g7_core_139;
  assign popcount38_j2g7_core_143 = input_a[34] & input_a[27];
  assign popcount38_j2g7_core_144 = input_a[18] ^ input_a[9];
  assign popcount38_j2g7_core_146 = input_a[28] & input_a[26];
  assign popcount38_j2g7_core_148 = ~(input_a[26] & input_a[7]);
  assign popcount38_j2g7_core_149 = input_a[15] ^ input_a[2];
  assign popcount38_j2g7_core_150 = ~(input_a[5] | input_a[17]);
  assign popcount38_j2g7_core_156 = input_a[19] & input_a[21];
  assign popcount38_j2g7_core_157 = ~input_a[36];
  assign popcount38_j2g7_core_158 = input_a[28] & input_a[15];
  assign popcount38_j2g7_core_159 = input_a[15] | input_a[12];
  assign popcount38_j2g7_core_160 = input_a[0] & input_a[8];
  assign popcount38_j2g7_core_161 = popcount38_j2g7_core_156 ^ popcount38_j2g7_core_158;
  assign popcount38_j2g7_core_162 = popcount38_j2g7_core_156 & popcount38_j2g7_core_158;
  assign popcount38_j2g7_core_163 = popcount38_j2g7_core_161 | popcount38_j2g7_core_160;
  assign popcount38_j2g7_core_164 = ~(input_a[16] ^ input_a[27]);
  assign popcount38_j2g7_core_166 = input_a[31] & input_a[2];
  assign popcount38_j2g7_core_167 = input_a[32] & input_a[30];
  assign popcount38_j2g7_core_169 = input_a[13] & input_a[2];
  assign popcount38_j2g7_core_171 = input_a[6] & input_a[34];
  assign popcount38_j2g7_core_172 = popcount38_j2g7_core_169 ^ popcount38_j2g7_core_171;
  assign popcount38_j2g7_core_173 = popcount38_j2g7_core_169 & popcount38_j2g7_core_171;
  assign popcount38_j2g7_core_175 = ~(input_a[9] | input_a[31]);
  assign popcount38_j2g7_core_176 = popcount38_j2g7_core_167 ^ popcount38_j2g7_core_172;
  assign popcount38_j2g7_core_177 = popcount38_j2g7_core_167 & popcount38_j2g7_core_172;
  assign popcount38_j2g7_core_181 = popcount38_j2g7_core_173 | popcount38_j2g7_core_177;
  assign popcount38_j2g7_core_183 = input_a[1] & input_a[14];
  assign popcount38_j2g7_core_184 = input_a[20] & input_a[26];
  assign popcount38_j2g7_core_185 = popcount38_j2g7_core_163 ^ popcount38_j2g7_core_176;
  assign popcount38_j2g7_core_186 = popcount38_j2g7_core_163 & popcount38_j2g7_core_176;
  assign popcount38_j2g7_core_187 = popcount38_j2g7_core_185 ^ popcount38_j2g7_core_184;
  assign popcount38_j2g7_core_188 = popcount38_j2g7_core_185 & popcount38_j2g7_core_184;
  assign popcount38_j2g7_core_189 = popcount38_j2g7_core_186 | popcount38_j2g7_core_188;
  assign popcount38_j2g7_core_190 = popcount38_j2g7_core_162 ^ popcount38_j2g7_core_181;
  assign popcount38_j2g7_core_191 = popcount38_j2g7_core_162 & popcount38_j2g7_core_181;
  assign popcount38_j2g7_core_192 = popcount38_j2g7_core_190 ^ popcount38_j2g7_core_189;
  assign popcount38_j2g7_core_193 = popcount38_j2g7_core_190 & popcount38_j2g7_core_189;
  assign popcount38_j2g7_core_194 = popcount38_j2g7_core_191 | popcount38_j2g7_core_193;
  assign popcount38_j2g7_core_197 = ~(input_a[28] | input_a[33]);
  assign popcount38_j2g7_core_198 = input_a[36] & input_a[7];
  assign popcount38_j2g7_core_199_not = ~input_a[20];
  assign popcount38_j2g7_core_200 = input_a[33] & input_a[25];
  assign popcount38_j2g7_core_201_not = ~input_a[6];
  assign popcount38_j2g7_core_202 = input_a[4] & input_a[1];
  assign popcount38_j2g7_core_203 = popcount38_j2g7_core_200 | popcount38_j2g7_core_202;
  assign popcount38_j2g7_core_205 = ~(input_a[1] & input_a[11]);
  assign popcount38_j2g7_core_206 = ~(input_a[29] & input_a[1]);
  assign popcount38_j2g7_core_207 = popcount38_j2g7_core_198 ^ popcount38_j2g7_core_203;
  assign popcount38_j2g7_core_208 = popcount38_j2g7_core_198 & popcount38_j2g7_core_203;
  assign popcount38_j2g7_core_214 = input_a[22] | input_a[8];
  assign popcount38_j2g7_core_215 = input_a[29] & input_a[35];
  assign popcount38_j2g7_core_217 = input_a[16] & input_a[31];
  assign popcount38_j2g7_core_218 = ~(input_a[30] & input_a[0]);
  assign popcount38_j2g7_core_219 = input_a[18] & input_a[5];
  assign popcount38_j2g7_core_220 = popcount38_j2g7_core_217 | popcount38_j2g7_core_219;
  assign popcount38_j2g7_core_223 = input_a[14] & input_a[23];
  assign popcount38_j2g7_core_224 = popcount38_j2g7_core_215 ^ popcount38_j2g7_core_220;
  assign popcount38_j2g7_core_225 = popcount38_j2g7_core_215 & popcount38_j2g7_core_220;
  assign popcount38_j2g7_core_226 = popcount38_j2g7_core_224 ^ popcount38_j2g7_core_223;
  assign popcount38_j2g7_core_227 = popcount38_j2g7_core_224 & popcount38_j2g7_core_223;
  assign popcount38_j2g7_core_228 = popcount38_j2g7_core_225 | popcount38_j2g7_core_227;
  assign popcount38_j2g7_core_230 = ~(input_a[10] | input_a[27]);
  assign popcount38_j2g7_core_233 = popcount38_j2g7_core_207 ^ popcount38_j2g7_core_226;
  assign popcount38_j2g7_core_234 = popcount38_j2g7_core_207 & popcount38_j2g7_core_226;
  assign popcount38_j2g7_core_238 = popcount38_j2g7_core_208 ^ popcount38_j2g7_core_228;
  assign popcount38_j2g7_core_239 = popcount38_j2g7_core_208 & popcount38_j2g7_core_228;
  assign popcount38_j2g7_core_240 = popcount38_j2g7_core_238 ^ popcount38_j2g7_core_234;
  assign popcount38_j2g7_core_241 = popcount38_j2g7_core_238 & popcount38_j2g7_core_234;
  assign popcount38_j2g7_core_242 = popcount38_j2g7_core_239 | popcount38_j2g7_core_241;
  assign popcount38_j2g7_core_244 = input_a[14] ^ input_a[19];
  assign popcount38_j2g7_core_246 = ~(input_a[33] & input_a[26]);
  assign popcount38_j2g7_core_247 = ~(input_a[4] ^ input_a[28]);
  assign popcount38_j2g7_core_248 = input_a[17] ^ input_a[11];
  assign popcount38_j2g7_core_249 = input_a[17] & input_a[11];
  assign popcount38_j2g7_core_250 = popcount38_j2g7_core_187 ^ popcount38_j2g7_core_233;
  assign popcount38_j2g7_core_251 = popcount38_j2g7_core_187 & popcount38_j2g7_core_233;
  assign popcount38_j2g7_core_252 = popcount38_j2g7_core_250 ^ popcount38_j2g7_core_249;
  assign popcount38_j2g7_core_253 = popcount38_j2g7_core_250 & popcount38_j2g7_core_249;
  assign popcount38_j2g7_core_254 = popcount38_j2g7_core_251 | popcount38_j2g7_core_253;
  assign popcount38_j2g7_core_255 = popcount38_j2g7_core_192 ^ popcount38_j2g7_core_240;
  assign popcount38_j2g7_core_256 = popcount38_j2g7_core_192 & popcount38_j2g7_core_240;
  assign popcount38_j2g7_core_257 = popcount38_j2g7_core_255 ^ popcount38_j2g7_core_254;
  assign popcount38_j2g7_core_258 = popcount38_j2g7_core_255 & popcount38_j2g7_core_254;
  assign popcount38_j2g7_core_259 = popcount38_j2g7_core_256 | popcount38_j2g7_core_258;
  assign popcount38_j2g7_core_260 = popcount38_j2g7_core_194 ^ popcount38_j2g7_core_242;
  assign popcount38_j2g7_core_261 = popcount38_j2g7_core_194 & popcount38_j2g7_core_242;
  assign popcount38_j2g7_core_262 = popcount38_j2g7_core_260 ^ popcount38_j2g7_core_259;
  assign popcount38_j2g7_core_263 = popcount38_j2g7_core_260 & popcount38_j2g7_core_259;
  assign popcount38_j2g7_core_264 = popcount38_j2g7_core_261 | popcount38_j2g7_core_263;
  assign popcount38_j2g7_core_266 = ~(input_a[36] & input_a[20]);
  assign popcount38_j2g7_core_268 = ~(input_a[34] | input_a[22]);
  assign popcount38_j2g7_core_271 = popcount38_j2g7_core_133 & popcount38_j2g7_core_248;
  assign popcount38_j2g7_core_272 = popcount38_j2g7_core_137 ^ popcount38_j2g7_core_252;
  assign popcount38_j2g7_core_273 = popcount38_j2g7_core_137 & popcount38_j2g7_core_252;
  assign popcount38_j2g7_core_274 = popcount38_j2g7_core_272 ^ popcount38_j2g7_core_271;
  assign popcount38_j2g7_core_275 = popcount38_j2g7_core_272 & popcount38_j2g7_core_271;
  assign popcount38_j2g7_core_276 = popcount38_j2g7_core_273 | popcount38_j2g7_core_275;
  assign popcount38_j2g7_core_277 = popcount38_j2g7_core_142 ^ popcount38_j2g7_core_257;
  assign popcount38_j2g7_core_278 = popcount38_j2g7_core_142 & popcount38_j2g7_core_257;
  assign popcount38_j2g7_core_279 = popcount38_j2g7_core_277 ^ popcount38_j2g7_core_276;
  assign popcount38_j2g7_core_280 = popcount38_j2g7_core_277 & popcount38_j2g7_core_276;
  assign popcount38_j2g7_core_281 = popcount38_j2g7_core_278 | popcount38_j2g7_core_280;
  assign popcount38_j2g7_core_282_not = ~popcount38_j2g7_core_262;
  assign popcount38_j2g7_core_284 = popcount38_j2g7_core_282_not ^ popcount38_j2g7_core_281;
  assign popcount38_j2g7_core_285 = popcount38_j2g7_core_282_not & popcount38_j2g7_core_281;
  assign popcount38_j2g7_core_286 = popcount38_j2g7_core_262 | popcount38_j2g7_core_285;
  assign popcount38_j2g7_core_289 = popcount38_j2g7_core_264 ^ popcount38_j2g7_core_286;
  assign popcount38_j2g7_core_290 = popcount38_j2g7_core_264 & popcount38_j2g7_core_286;
  assign popcount38_j2g7_core_292 = input_a[4] & input_a[26];
  assign popcount38_j2g7_core_293 = ~(input_a[13] | input_a[28]);
  assign popcount38_j2g7_core_296 = ~(input_a[26] | input_a[29]);

  assign popcount38_j2g7_out[0] = input_a[37];
  assign popcount38_j2g7_out[1] = popcount38_j2g7_core_274;
  assign popcount38_j2g7_out[2] = popcount38_j2g7_core_279;
  assign popcount38_j2g7_out[3] = popcount38_j2g7_core_284;
  assign popcount38_j2g7_out[4] = popcount38_j2g7_core_289;
  assign popcount38_j2g7_out[5] = popcount38_j2g7_core_290;
endmodule