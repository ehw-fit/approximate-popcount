// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.71472
// WCE=9.0
// EP=0.968254%
// Printed PDK parameters:
//  Area=22964282.0
//  Delay=45631804.0
//  Power=1201900.0

module popcount18_88r5(input [17:0] input_a, output [4:0] popcount18_88r5_out);
  wire popcount18_88r5_core_020;
  wire popcount18_88r5_core_021;
  wire popcount18_88r5_core_022;
  wire popcount18_88r5_core_023;
  wire popcount18_88r5_core_024;
  wire popcount18_88r5_core_025;
  wire popcount18_88r5_core_026;
  wire popcount18_88r5_core_027;
  wire popcount18_88r5_core_028;
  wire popcount18_88r5_core_031;
  wire popcount18_88r5_core_032;
  wire popcount18_88r5_core_033;
  wire popcount18_88r5_core_034;
  wire popcount18_88r5_core_035_not;
  wire popcount18_88r5_core_036;
  wire popcount18_88r5_core_037;
  wire popcount18_88r5_core_039;
  wire popcount18_88r5_core_041;
  wire popcount18_88r5_core_042;
  wire popcount18_88r5_core_044;
  wire popcount18_88r5_core_048;
  wire popcount18_88r5_core_049;
  wire popcount18_88r5_core_050;
  wire popcount18_88r5_core_051;
  wire popcount18_88r5_core_052;
  wire popcount18_88r5_core_053;
  wire popcount18_88r5_core_054;
  wire popcount18_88r5_core_055;
  wire popcount18_88r5_core_056;
  wire popcount18_88r5_core_057;
  wire popcount18_88r5_core_058;
  wire popcount18_88r5_core_059;
  wire popcount18_88r5_core_063;
  wire popcount18_88r5_core_064;
  wire popcount18_88r5_core_065;
  wire popcount18_88r5_core_066;
  wire popcount18_88r5_core_068;
  wire popcount18_88r5_core_069;
  wire popcount18_88r5_core_070;
  wire popcount18_88r5_core_071;
  wire popcount18_88r5_core_072;
  wire popcount18_88r5_core_073;
  wire popcount18_88r5_core_074;
  wire popcount18_88r5_core_075;
  wire popcount18_88r5_core_076;
  wire popcount18_88r5_core_081;
  wire popcount18_88r5_core_082;
  wire popcount18_88r5_core_083;
  wire popcount18_88r5_core_084;
  wire popcount18_88r5_core_085;
  wire popcount18_88r5_core_086;
  wire popcount18_88r5_core_087;
  wire popcount18_88r5_core_090;
  wire popcount18_88r5_core_094;
  wire popcount18_88r5_core_095;
  wire popcount18_88r5_core_099_not;
  wire popcount18_88r5_core_104;
  wire popcount18_88r5_core_106;
  wire popcount18_88r5_core_109;
  wire popcount18_88r5_core_111;
  wire popcount18_88r5_core_113;
  wire popcount18_88r5_core_114;
  wire popcount18_88r5_core_116;
  wire popcount18_88r5_core_117;
  wire popcount18_88r5_core_118;
  wire popcount18_88r5_core_119;
  wire popcount18_88r5_core_120;
  wire popcount18_88r5_core_122;
  wire popcount18_88r5_core_123;
  wire popcount18_88r5_core_124;
  wire popcount18_88r5_core_125;

  assign popcount18_88r5_core_020 = input_a[0] ^ input_a[1];
  assign popcount18_88r5_core_021 = input_a[0] & input_a[1];
  assign popcount18_88r5_core_022 = input_a[2] ^ input_a[3];
  assign popcount18_88r5_core_023 = input_a[2] & input_a[3];
  assign popcount18_88r5_core_024 = popcount18_88r5_core_020 ^ popcount18_88r5_core_022;
  assign popcount18_88r5_core_025 = popcount18_88r5_core_020 & popcount18_88r5_core_022;
  assign popcount18_88r5_core_026 = popcount18_88r5_core_021 ^ popcount18_88r5_core_023;
  assign popcount18_88r5_core_027 = popcount18_88r5_core_021 & popcount18_88r5_core_023;
  assign popcount18_88r5_core_028 = popcount18_88r5_core_026 | popcount18_88r5_core_025;
  assign popcount18_88r5_core_031 = ~(input_a[4] | input_a[4]);
  assign popcount18_88r5_core_032 = input_a[16] & input_a[8];
  assign popcount18_88r5_core_033 = ~(input_a[6] ^ input_a[2]);
  assign popcount18_88r5_core_034 = input_a[15] & input_a[5];
  assign popcount18_88r5_core_035_not = ~input_a[9];
  assign popcount18_88r5_core_036 = input_a[6] & input_a[17];
  assign popcount18_88r5_core_037 = popcount18_88r5_core_034 | popcount18_88r5_core_036;
  assign popcount18_88r5_core_039 = ~(input_a[14] & input_a[13]);
  assign popcount18_88r5_core_041 = popcount18_88r5_core_032 ^ popcount18_88r5_core_037;
  assign popcount18_88r5_core_042 = popcount18_88r5_core_032 & popcount18_88r5_core_037;
  assign popcount18_88r5_core_044 = ~input_a[15];
  assign popcount18_88r5_core_048 = input_a[7] & input_a[9];
  assign popcount18_88r5_core_049 = popcount18_88r5_core_024 & input_a[7];
  assign popcount18_88r5_core_050 = popcount18_88r5_core_028 ^ popcount18_88r5_core_041;
  assign popcount18_88r5_core_051 = popcount18_88r5_core_028 & popcount18_88r5_core_041;
  assign popcount18_88r5_core_052 = popcount18_88r5_core_050 ^ popcount18_88r5_core_049;
  assign popcount18_88r5_core_053 = popcount18_88r5_core_050 & popcount18_88r5_core_049;
  assign popcount18_88r5_core_054 = popcount18_88r5_core_051 | popcount18_88r5_core_053;
  assign popcount18_88r5_core_055 = popcount18_88r5_core_027 ^ popcount18_88r5_core_042;
  assign popcount18_88r5_core_056 = popcount18_88r5_core_027 & popcount18_88r5_core_042;
  assign popcount18_88r5_core_057 = popcount18_88r5_core_055 ^ popcount18_88r5_core_054;
  assign popcount18_88r5_core_058 = popcount18_88r5_core_055 & popcount18_88r5_core_054;
  assign popcount18_88r5_core_059 = popcount18_88r5_core_056 | popcount18_88r5_core_058;
  assign popcount18_88r5_core_063 = input_a[9] & input_a[10];
  assign popcount18_88r5_core_064 = input_a[11] ^ input_a[12];
  assign popcount18_88r5_core_065 = input_a[11] & input_a[12];
  assign popcount18_88r5_core_066 = ~(input_a[9] & input_a[10]);
  assign popcount18_88r5_core_068 = popcount18_88r5_core_063 ^ popcount18_88r5_core_065;
  assign popcount18_88r5_core_069 = popcount18_88r5_core_063 & input_a[11];
  assign popcount18_88r5_core_070 = popcount18_88r5_core_068 ^ popcount18_88r5_core_064;
  assign popcount18_88r5_core_071 = popcount18_88r5_core_068 & popcount18_88r5_core_064;
  assign popcount18_88r5_core_072 = popcount18_88r5_core_069 | popcount18_88r5_core_071;
  assign popcount18_88r5_core_073 = ~(input_a[3] ^ input_a[7]);
  assign popcount18_88r5_core_074 = input_a[17] | input_a[9];
  assign popcount18_88r5_core_075 = input_a[7] | input_a[8];
  assign popcount18_88r5_core_076 = ~(input_a[14] | input_a[3]);
  assign popcount18_88r5_core_081 = ~(input_a[3] | input_a[0]);
  assign popcount18_88r5_core_082 = ~input_a[10];
  assign popcount18_88r5_core_083 = input_a[8] ^ input_a[11];
  assign popcount18_88r5_core_084 = input_a[6] ^ input_a[5];
  assign popcount18_88r5_core_085 = input_a[2] ^ input_a[16];
  assign popcount18_88r5_core_086 = ~input_a[5];
  assign popcount18_88r5_core_087 = ~(input_a[6] | input_a[16]);
  assign popcount18_88r5_core_090 = input_a[12] & input_a[1];
  assign popcount18_88r5_core_094 = popcount18_88r5_core_070 | popcount18_88r5_core_066;
  assign popcount18_88r5_core_095 = ~input_a[3];
  assign popcount18_88r5_core_099_not = ~popcount18_88r5_core_070;
  assign popcount18_88r5_core_104 = input_a[3] | input_a[15];
  assign popcount18_88r5_core_106 = popcount18_88r5_core_052 ^ popcount18_88r5_core_094;
  assign popcount18_88r5_core_109 = input_a[2] & input_a[0];
  assign popcount18_88r5_core_111 = popcount18_88r5_core_057 ^ popcount18_88r5_core_099_not;
  assign popcount18_88r5_core_113 = popcount18_88r5_core_111 ^ popcount18_88r5_core_052;
  assign popcount18_88r5_core_114 = popcount18_88r5_core_111 & popcount18_88r5_core_052;
  assign popcount18_88r5_core_116 = popcount18_88r5_core_059 | popcount18_88r5_core_070;
  assign popcount18_88r5_core_117 = popcount18_88r5_core_059 & popcount18_88r5_core_070;
  assign popcount18_88r5_core_118 = ~(input_a[10] ^ input_a[6]);
  assign popcount18_88r5_core_119 = popcount18_88r5_core_116 & popcount18_88r5_core_114;
  assign popcount18_88r5_core_120 = popcount18_88r5_core_117 | popcount18_88r5_core_119;
  assign popcount18_88r5_core_122 = input_a[6] & input_a[7];
  assign popcount18_88r5_core_123 = input_a[10] & input_a[7];
  assign popcount18_88r5_core_124 = input_a[1] & input_a[1];
  assign popcount18_88r5_core_125 = input_a[1] | input_a[6];

  assign popcount18_88r5_out[0] = input_a[4];
  assign popcount18_88r5_out[1] = popcount18_88r5_core_106;
  assign popcount18_88r5_out[2] = popcount18_88r5_core_113;
  assign popcount18_88r5_out[3] = popcount18_88r5_core_072;
  assign popcount18_88r5_out[4] = popcount18_88r5_core_120;
endmodule