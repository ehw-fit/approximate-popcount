// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.52066
// WCE=16.0
// EP=0.876707%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_aqmn(input [27:0] input_a, output [4:0] popcount28_aqmn_out);
  wire popcount28_aqmn_core_030;
  wire popcount28_aqmn_core_032;
  wire popcount28_aqmn_core_033;
  wire popcount28_aqmn_core_034;
  wire popcount28_aqmn_core_035;
  wire popcount28_aqmn_core_036;
  wire popcount28_aqmn_core_037;
  wire popcount28_aqmn_core_038;
  wire popcount28_aqmn_core_039;
  wire popcount28_aqmn_core_040;
  wire popcount28_aqmn_core_041;
  wire popcount28_aqmn_core_042;
  wire popcount28_aqmn_core_043;
  wire popcount28_aqmn_core_044;
  wire popcount28_aqmn_core_045;
  wire popcount28_aqmn_core_046;
  wire popcount28_aqmn_core_048;
  wire popcount28_aqmn_core_050;
  wire popcount28_aqmn_core_051;
  wire popcount28_aqmn_core_052;
  wire popcount28_aqmn_core_054;
  wire popcount28_aqmn_core_057;
  wire popcount28_aqmn_core_058;
  wire popcount28_aqmn_core_060;
  wire popcount28_aqmn_core_061;
  wire popcount28_aqmn_core_063_not;
  wire popcount28_aqmn_core_065;
  wire popcount28_aqmn_core_066;
  wire popcount28_aqmn_core_067;
  wire popcount28_aqmn_core_068;
  wire popcount28_aqmn_core_070_not;
  wire popcount28_aqmn_core_071;
  wire popcount28_aqmn_core_072;
  wire popcount28_aqmn_core_073;
  wire popcount28_aqmn_core_074;
  wire popcount28_aqmn_core_076;
  wire popcount28_aqmn_core_078;
  wire popcount28_aqmn_core_079;
  wire popcount28_aqmn_core_080;
  wire popcount28_aqmn_core_082;
  wire popcount28_aqmn_core_083;
  wire popcount28_aqmn_core_084;
  wire popcount28_aqmn_core_085;
  wire popcount28_aqmn_core_086;
  wire popcount28_aqmn_core_087;
  wire popcount28_aqmn_core_088;
  wire popcount28_aqmn_core_089;
  wire popcount28_aqmn_core_090;
  wire popcount28_aqmn_core_092;
  wire popcount28_aqmn_core_093;
  wire popcount28_aqmn_core_094;
  wire popcount28_aqmn_core_095;
  wire popcount28_aqmn_core_096;
  wire popcount28_aqmn_core_098;
  wire popcount28_aqmn_core_099_not;
  wire popcount28_aqmn_core_100;
  wire popcount28_aqmn_core_101;
  wire popcount28_aqmn_core_102;
  wire popcount28_aqmn_core_103;
  wire popcount28_aqmn_core_104;
  wire popcount28_aqmn_core_105;
  wire popcount28_aqmn_core_108;
  wire popcount28_aqmn_core_110;
  wire popcount28_aqmn_core_111_not;
  wire popcount28_aqmn_core_112_not;
  wire popcount28_aqmn_core_113;
  wire popcount28_aqmn_core_115;
  wire popcount28_aqmn_core_116;
  wire popcount28_aqmn_core_117;
  wire popcount28_aqmn_core_120;
  wire popcount28_aqmn_core_122;
  wire popcount28_aqmn_core_125;
  wire popcount28_aqmn_core_127;
  wire popcount28_aqmn_core_128;
  wire popcount28_aqmn_core_131;
  wire popcount28_aqmn_core_132;
  wire popcount28_aqmn_core_133;
  wire popcount28_aqmn_core_134;
  wire popcount28_aqmn_core_136_not;
  wire popcount28_aqmn_core_140;
  wire popcount28_aqmn_core_141;
  wire popcount28_aqmn_core_142;
  wire popcount28_aqmn_core_145;
  wire popcount28_aqmn_core_146;
  wire popcount28_aqmn_core_147;
  wire popcount28_aqmn_core_148;
  wire popcount28_aqmn_core_149;
  wire popcount28_aqmn_core_150;
  wire popcount28_aqmn_core_151;
  wire popcount28_aqmn_core_153;
  wire popcount28_aqmn_core_154;
  wire popcount28_aqmn_core_155;
  wire popcount28_aqmn_core_156;
  wire popcount28_aqmn_core_158;
  wire popcount28_aqmn_core_160;
  wire popcount28_aqmn_core_162;
  wire popcount28_aqmn_core_163;
  wire popcount28_aqmn_core_164;
  wire popcount28_aqmn_core_165;
  wire popcount28_aqmn_core_166;
  wire popcount28_aqmn_core_167;
  wire popcount28_aqmn_core_170;
  wire popcount28_aqmn_core_171;
  wire popcount28_aqmn_core_172;
  wire popcount28_aqmn_core_173;
  wire popcount28_aqmn_core_174;
  wire popcount28_aqmn_core_175;
  wire popcount28_aqmn_core_176;
  wire popcount28_aqmn_core_177;
  wire popcount28_aqmn_core_179;
  wire popcount28_aqmn_core_180;
  wire popcount28_aqmn_core_182;
  wire popcount28_aqmn_core_183;
  wire popcount28_aqmn_core_184;
  wire popcount28_aqmn_core_186;
  wire popcount28_aqmn_core_187_not;
  wire popcount28_aqmn_core_188;
  wire popcount28_aqmn_core_189;
  wire popcount28_aqmn_core_192;
  wire popcount28_aqmn_core_193;
  wire popcount28_aqmn_core_194_not;
  wire popcount28_aqmn_core_197;
  wire popcount28_aqmn_core_198;
  wire popcount28_aqmn_core_199;
  wire popcount28_aqmn_core_200;
  wire popcount28_aqmn_core_201;

  assign popcount28_aqmn_core_030 = input_a[4] & input_a[13];
  assign popcount28_aqmn_core_032 = input_a[11] | input_a[23];
  assign popcount28_aqmn_core_033 = ~(input_a[7] | input_a[26]);
  assign popcount28_aqmn_core_034 = input_a[10] & input_a[15];
  assign popcount28_aqmn_core_035 = input_a[18] | input_a[1];
  assign popcount28_aqmn_core_036 = ~(input_a[14] ^ input_a[20]);
  assign popcount28_aqmn_core_037 = ~(input_a[11] | input_a[2]);
  assign popcount28_aqmn_core_038 = input_a[1] ^ input_a[3];
  assign popcount28_aqmn_core_039 = ~(input_a[0] & input_a[27]);
  assign popcount28_aqmn_core_040 = ~(input_a[19] ^ input_a[13]);
  assign popcount28_aqmn_core_041 = input_a[6] ^ input_a[13];
  assign popcount28_aqmn_core_042 = ~(input_a[23] | input_a[26]);
  assign popcount28_aqmn_core_043 = input_a[8] | input_a[0];
  assign popcount28_aqmn_core_044 = input_a[3] & input_a[15];
  assign popcount28_aqmn_core_045 = input_a[20] ^ input_a[16];
  assign popcount28_aqmn_core_046 = input_a[17] | input_a[7];
  assign popcount28_aqmn_core_048 = ~(input_a[4] & input_a[8]);
  assign popcount28_aqmn_core_050 = input_a[1] & input_a[18];
  assign popcount28_aqmn_core_051 = ~(input_a[5] ^ input_a[0]);
  assign popcount28_aqmn_core_052 = input_a[4] | input_a[19];
  assign popcount28_aqmn_core_054 = input_a[19] & input_a[16];
  assign popcount28_aqmn_core_057 = ~input_a[19];
  assign popcount28_aqmn_core_058 = input_a[13] & input_a[24];
  assign popcount28_aqmn_core_060 = input_a[26] ^ input_a[25];
  assign popcount28_aqmn_core_061 = ~(input_a[26] & input_a[2]);
  assign popcount28_aqmn_core_063_not = ~input_a[15];
  assign popcount28_aqmn_core_065 = ~input_a[4];
  assign popcount28_aqmn_core_066 = ~(input_a[20] | input_a[13]);
  assign popcount28_aqmn_core_067 = ~(input_a[10] ^ input_a[15]);
  assign popcount28_aqmn_core_068 = input_a[7] | input_a[20];
  assign popcount28_aqmn_core_070_not = ~input_a[26];
  assign popcount28_aqmn_core_071 = ~(input_a[11] ^ input_a[27]);
  assign popcount28_aqmn_core_072 = ~(input_a[15] | input_a[7]);
  assign popcount28_aqmn_core_073 = ~input_a[18];
  assign popcount28_aqmn_core_074 = input_a[9] & input_a[7];
  assign popcount28_aqmn_core_076 = ~(input_a[18] ^ input_a[0]);
  assign popcount28_aqmn_core_078 = ~(input_a[17] & input_a[5]);
  assign popcount28_aqmn_core_079 = ~input_a[25];
  assign popcount28_aqmn_core_080 = input_a[4] & input_a[26];
  assign popcount28_aqmn_core_082 = input_a[23] | input_a[6];
  assign popcount28_aqmn_core_083 = ~input_a[6];
  assign popcount28_aqmn_core_084 = ~(input_a[14] ^ input_a[7]);
  assign popcount28_aqmn_core_085 = ~input_a[2];
  assign popcount28_aqmn_core_086 = ~(input_a[18] | input_a[23]);
  assign popcount28_aqmn_core_087 = ~input_a[26];
  assign popcount28_aqmn_core_088 = ~(input_a[4] & input_a[5]);
  assign popcount28_aqmn_core_089 = ~input_a[8];
  assign popcount28_aqmn_core_090 = ~(input_a[10] & input_a[3]);
  assign popcount28_aqmn_core_092 = ~(input_a[18] & input_a[14]);
  assign popcount28_aqmn_core_093 = input_a[9] | input_a[17];
  assign popcount28_aqmn_core_094 = ~input_a[17];
  assign popcount28_aqmn_core_095 = ~(input_a[24] | input_a[5]);
  assign popcount28_aqmn_core_096 = ~(input_a[2] ^ input_a[15]);
  assign popcount28_aqmn_core_098 = ~input_a[1];
  assign popcount28_aqmn_core_099_not = ~input_a[8];
  assign popcount28_aqmn_core_100 = input_a[11] & input_a[7];
  assign popcount28_aqmn_core_101 = ~input_a[9];
  assign popcount28_aqmn_core_102 = ~input_a[19];
  assign popcount28_aqmn_core_103 = ~(input_a[11] & input_a[0]);
  assign popcount28_aqmn_core_104 = input_a[27] ^ input_a[5];
  assign popcount28_aqmn_core_105 = input_a[20] & input_a[10];
  assign popcount28_aqmn_core_108 = ~(input_a[13] & input_a[21]);
  assign popcount28_aqmn_core_110 = input_a[1] & input_a[19];
  assign popcount28_aqmn_core_111_not = ~input_a[9];
  assign popcount28_aqmn_core_112_not = ~input_a[11];
  assign popcount28_aqmn_core_113 = input_a[14] ^ input_a[3];
  assign popcount28_aqmn_core_115 = input_a[9] ^ input_a[2];
  assign popcount28_aqmn_core_116 = ~(input_a[26] ^ input_a[18]);
  assign popcount28_aqmn_core_117 = ~(input_a[27] & input_a[0]);
  assign popcount28_aqmn_core_120 = ~(input_a[2] & input_a[25]);
  assign popcount28_aqmn_core_122 = input_a[4] & input_a[4];
  assign popcount28_aqmn_core_125 = input_a[2] | input_a[18];
  assign popcount28_aqmn_core_127 = input_a[10] | input_a[16];
  assign popcount28_aqmn_core_128 = input_a[17] & input_a[1];
  assign popcount28_aqmn_core_131 = ~input_a[23];
  assign popcount28_aqmn_core_132 = ~input_a[6];
  assign popcount28_aqmn_core_133 = input_a[13] | input_a[3];
  assign popcount28_aqmn_core_134 = ~input_a[6];
  assign popcount28_aqmn_core_136_not = ~input_a[21];
  assign popcount28_aqmn_core_140 = input_a[0] & input_a[6];
  assign popcount28_aqmn_core_141 = ~(input_a[6] & input_a[23]);
  assign popcount28_aqmn_core_142 = input_a[17] ^ input_a[20];
  assign popcount28_aqmn_core_145 = ~(input_a[16] | input_a[20]);
  assign popcount28_aqmn_core_146 = input_a[20] & input_a[6];
  assign popcount28_aqmn_core_147 = ~input_a[24];
  assign popcount28_aqmn_core_148 = ~(input_a[13] ^ input_a[25]);
  assign popcount28_aqmn_core_149 = input_a[4] ^ input_a[3];
  assign popcount28_aqmn_core_150 = ~input_a[4];
  assign popcount28_aqmn_core_151 = input_a[14] & input_a[22];
  assign popcount28_aqmn_core_153 = input_a[17] & input_a[27];
  assign popcount28_aqmn_core_154 = ~(input_a[16] ^ input_a[1]);
  assign popcount28_aqmn_core_155 = ~input_a[13];
  assign popcount28_aqmn_core_156 = ~input_a[13];
  assign popcount28_aqmn_core_158 = input_a[10] & input_a[9];
  assign popcount28_aqmn_core_160 = input_a[24] ^ input_a[11];
  assign popcount28_aqmn_core_162 = ~(input_a[2] | input_a[24]);
  assign popcount28_aqmn_core_163 = ~(input_a[9] & input_a[23]);
  assign popcount28_aqmn_core_164 = ~(input_a[3] ^ input_a[15]);
  assign popcount28_aqmn_core_165 = ~(input_a[0] & input_a[10]);
  assign popcount28_aqmn_core_166 = ~input_a[7];
  assign popcount28_aqmn_core_167 = input_a[26] & input_a[27];
  assign popcount28_aqmn_core_170 = ~(input_a[22] | input_a[25]);
  assign popcount28_aqmn_core_171 = ~(input_a[5] & input_a[0]);
  assign popcount28_aqmn_core_172 = input_a[12] & input_a[3];
  assign popcount28_aqmn_core_173 = ~(input_a[17] & input_a[12]);
  assign popcount28_aqmn_core_174 = ~(input_a[13] & input_a[6]);
  assign popcount28_aqmn_core_175 = ~(input_a[16] & input_a[1]);
  assign popcount28_aqmn_core_176 = input_a[17] | input_a[23];
  assign popcount28_aqmn_core_177 = ~input_a[13];
  assign popcount28_aqmn_core_179 = input_a[25] ^ input_a[22];
  assign popcount28_aqmn_core_180 = ~(input_a[5] | input_a[25]);
  assign popcount28_aqmn_core_182 = ~(input_a[10] & input_a[15]);
  assign popcount28_aqmn_core_183 = input_a[12] | input_a[23];
  assign popcount28_aqmn_core_184 = ~(input_a[3] & input_a[25]);
  assign popcount28_aqmn_core_186 = ~(input_a[14] & input_a[0]);
  assign popcount28_aqmn_core_187_not = ~input_a[6];
  assign popcount28_aqmn_core_188 = ~input_a[4];
  assign popcount28_aqmn_core_189 = ~(input_a[8] | input_a[6]);
  assign popcount28_aqmn_core_192 = ~(input_a[0] & input_a[12]);
  assign popcount28_aqmn_core_193 = ~(input_a[9] | input_a[12]);
  assign popcount28_aqmn_core_194_not = ~input_a[16];
  assign popcount28_aqmn_core_197 = input_a[24] | input_a[10];
  assign popcount28_aqmn_core_198 = input_a[6] | input_a[14];
  assign popcount28_aqmn_core_199 = input_a[25] ^ input_a[16];
  assign popcount28_aqmn_core_200 = input_a[7] | input_a[5];
  assign popcount28_aqmn_core_201 = ~(input_a[6] | input_a[20]);

  assign popcount28_aqmn_out[0] = 1'b1;
  assign popcount28_aqmn_out[1] = 1'b1;
  assign popcount28_aqmn_out[2] = input_a[14];
  assign popcount28_aqmn_out[3] = 1'b1;
  assign popcount28_aqmn_out[4] = 1'b0;
endmodule