// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.39114
// WCE=15.0
// EP=0.87048%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount29_4kz0(input [28:0] input_a, output [4:0] popcount29_4kz0_out);
  wire popcount29_4kz0_core_032;
  wire popcount29_4kz0_core_033;
  wire popcount29_4kz0_core_038_not;
  wire popcount29_4kz0_core_040;
  wire popcount29_4kz0_core_041;
  wire popcount29_4kz0_core_042;
  wire popcount29_4kz0_core_044;
  wire popcount29_4kz0_core_045;
  wire popcount29_4kz0_core_047;
  wire popcount29_4kz0_core_048;
  wire popcount29_4kz0_core_049;
  wire popcount29_4kz0_core_050;
  wire popcount29_4kz0_core_051;
  wire popcount29_4kz0_core_052;
  wire popcount29_4kz0_core_053;
  wire popcount29_4kz0_core_054;
  wire popcount29_4kz0_core_057;
  wire popcount29_4kz0_core_058;
  wire popcount29_4kz0_core_062;
  wire popcount29_4kz0_core_063;
  wire popcount29_4kz0_core_064;
  wire popcount29_4kz0_core_066;
  wire popcount29_4kz0_core_067;
  wire popcount29_4kz0_core_068;
  wire popcount29_4kz0_core_069;
  wire popcount29_4kz0_core_070;
  wire popcount29_4kz0_core_071;
  wire popcount29_4kz0_core_072;
  wire popcount29_4kz0_core_074;
  wire popcount29_4kz0_core_075;
  wire popcount29_4kz0_core_077;
  wire popcount29_4kz0_core_078;
  wire popcount29_4kz0_core_079;
  wire popcount29_4kz0_core_081;
  wire popcount29_4kz0_core_083;
  wire popcount29_4kz0_core_084;
  wire popcount29_4kz0_core_085;
  wire popcount29_4kz0_core_086;
  wire popcount29_4kz0_core_088;
  wire popcount29_4kz0_core_089;
  wire popcount29_4kz0_core_090;
  wire popcount29_4kz0_core_091;
  wire popcount29_4kz0_core_092;
  wire popcount29_4kz0_core_093;
  wire popcount29_4kz0_core_096;
  wire popcount29_4kz0_core_100;
  wire popcount29_4kz0_core_101;
  wire popcount29_4kz0_core_103;
  wire popcount29_4kz0_core_105;
  wire popcount29_4kz0_core_106;
  wire popcount29_4kz0_core_107;
  wire popcount29_4kz0_core_108;
  wire popcount29_4kz0_core_110;
  wire popcount29_4kz0_core_111;
  wire popcount29_4kz0_core_112;
  wire popcount29_4kz0_core_113;
  wire popcount29_4kz0_core_114;
  wire popcount29_4kz0_core_115;
  wire popcount29_4kz0_core_116;
  wire popcount29_4kz0_core_117;
  wire popcount29_4kz0_core_118;
  wire popcount29_4kz0_core_119;
  wire popcount29_4kz0_core_120;
  wire popcount29_4kz0_core_122;
  wire popcount29_4kz0_core_124;
  wire popcount29_4kz0_core_125;
  wire popcount29_4kz0_core_126;
  wire popcount29_4kz0_core_127;
  wire popcount29_4kz0_core_129;
  wire popcount29_4kz0_core_132;
  wire popcount29_4kz0_core_133;
  wire popcount29_4kz0_core_134;
  wire popcount29_4kz0_core_135;
  wire popcount29_4kz0_core_136;
  wire popcount29_4kz0_core_137;
  wire popcount29_4kz0_core_138;
  wire popcount29_4kz0_core_140;
  wire popcount29_4kz0_core_141;
  wire popcount29_4kz0_core_143;
  wire popcount29_4kz0_core_144;
  wire popcount29_4kz0_core_145;
  wire popcount29_4kz0_core_146;
  wire popcount29_4kz0_core_147;
  wire popcount29_4kz0_core_148;
  wire popcount29_4kz0_core_149;
  wire popcount29_4kz0_core_150;
  wire popcount29_4kz0_core_152;
  wire popcount29_4kz0_core_154;
  wire popcount29_4kz0_core_157;
  wire popcount29_4kz0_core_158;
  wire popcount29_4kz0_core_159;
  wire popcount29_4kz0_core_162;
  wire popcount29_4kz0_core_163;
  wire popcount29_4kz0_core_164;
  wire popcount29_4kz0_core_166;
  wire popcount29_4kz0_core_167;
  wire popcount29_4kz0_core_169;
  wire popcount29_4kz0_core_171;
  wire popcount29_4kz0_core_176_not;
  wire popcount29_4kz0_core_177;
  wire popcount29_4kz0_core_179;
  wire popcount29_4kz0_core_180;
  wire popcount29_4kz0_core_181;
  wire popcount29_4kz0_core_182;
  wire popcount29_4kz0_core_183;
  wire popcount29_4kz0_core_184;
  wire popcount29_4kz0_core_186;
  wire popcount29_4kz0_core_188;
  wire popcount29_4kz0_core_189;
  wire popcount29_4kz0_core_190;
  wire popcount29_4kz0_core_191;
  wire popcount29_4kz0_core_192;
  wire popcount29_4kz0_core_193;
  wire popcount29_4kz0_core_194;
  wire popcount29_4kz0_core_198;
  wire popcount29_4kz0_core_199;
  wire popcount29_4kz0_core_200;
  wire popcount29_4kz0_core_201;
  wire popcount29_4kz0_core_202;
  wire popcount29_4kz0_core_205;
  wire popcount29_4kz0_core_206;
  wire popcount29_4kz0_core_207;

  assign popcount29_4kz0_core_032 = ~(input_a[4] & input_a[13]);
  assign popcount29_4kz0_core_033 = input_a[19] | input_a[28];
  assign popcount29_4kz0_core_038_not = ~input_a[14];
  assign popcount29_4kz0_core_040 = ~(input_a[19] ^ input_a[26]);
  assign popcount29_4kz0_core_041 = input_a[28] ^ input_a[17];
  assign popcount29_4kz0_core_042 = input_a[0] ^ input_a[9];
  assign popcount29_4kz0_core_044 = ~(input_a[3] & input_a[23]);
  assign popcount29_4kz0_core_045 = ~(input_a[7] & input_a[4]);
  assign popcount29_4kz0_core_047 = ~input_a[8];
  assign popcount29_4kz0_core_048 = ~input_a[26];
  assign popcount29_4kz0_core_049 = ~input_a[9];
  assign popcount29_4kz0_core_050 = input_a[13] | input_a[4];
  assign popcount29_4kz0_core_051 = input_a[16] ^ input_a[9];
  assign popcount29_4kz0_core_052 = input_a[5] | input_a[16];
  assign popcount29_4kz0_core_053 = ~(input_a[16] & input_a[23]);
  assign popcount29_4kz0_core_054 = ~(input_a[16] | input_a[25]);
  assign popcount29_4kz0_core_057 = ~input_a[19];
  assign popcount29_4kz0_core_058 = ~(input_a[13] | input_a[20]);
  assign popcount29_4kz0_core_062 = input_a[5] & input_a[22];
  assign popcount29_4kz0_core_063 = input_a[20] ^ input_a[17];
  assign popcount29_4kz0_core_064 = ~input_a[8];
  assign popcount29_4kz0_core_066 = input_a[8] ^ input_a[18];
  assign popcount29_4kz0_core_067 = ~(input_a[14] ^ input_a[28]);
  assign popcount29_4kz0_core_068 = ~(input_a[19] | input_a[7]);
  assign popcount29_4kz0_core_069 = ~input_a[24];
  assign popcount29_4kz0_core_070 = ~(input_a[16] ^ input_a[19]);
  assign popcount29_4kz0_core_071 = ~(input_a[18] & input_a[24]);
  assign popcount29_4kz0_core_072 = ~input_a[11];
  assign popcount29_4kz0_core_074 = ~input_a[27];
  assign popcount29_4kz0_core_075 = input_a[22] ^ input_a[14];
  assign popcount29_4kz0_core_077 = ~(input_a[9] | input_a[3]);
  assign popcount29_4kz0_core_078 = input_a[26] | input_a[1];
  assign popcount29_4kz0_core_079 = ~(input_a[6] | input_a[21]);
  assign popcount29_4kz0_core_081 = ~(input_a[20] ^ input_a[18]);
  assign popcount29_4kz0_core_083 = ~input_a[22];
  assign popcount29_4kz0_core_084 = ~(input_a[12] ^ input_a[19]);
  assign popcount29_4kz0_core_085 = input_a[4] | input_a[3];
  assign popcount29_4kz0_core_086 = ~(input_a[26] | input_a[8]);
  assign popcount29_4kz0_core_088 = input_a[13] & input_a[2];
  assign popcount29_4kz0_core_089 = ~(input_a[4] ^ input_a[2]);
  assign popcount29_4kz0_core_090 = ~(input_a[4] ^ input_a[0]);
  assign popcount29_4kz0_core_091 = ~input_a[8];
  assign popcount29_4kz0_core_092 = ~(input_a[2] & input_a[16]);
  assign popcount29_4kz0_core_093 = ~input_a[16];
  assign popcount29_4kz0_core_096 = ~input_a[2];
  assign popcount29_4kz0_core_100 = ~(input_a[11] & input_a[4]);
  assign popcount29_4kz0_core_101 = input_a[10] & input_a[4];
  assign popcount29_4kz0_core_103 = ~(input_a[17] | input_a[20]);
  assign popcount29_4kz0_core_105 = input_a[7] ^ input_a[6];
  assign popcount29_4kz0_core_106 = input_a[11] ^ input_a[20];
  assign popcount29_4kz0_core_107 = ~(input_a[4] | input_a[9]);
  assign popcount29_4kz0_core_108 = input_a[9] | input_a[4];
  assign popcount29_4kz0_core_110 = input_a[1] ^ input_a[26];
  assign popcount29_4kz0_core_111 = ~input_a[17];
  assign popcount29_4kz0_core_112 = input_a[20] & input_a[14];
  assign popcount29_4kz0_core_113 = ~(input_a[5] ^ input_a[22]);
  assign popcount29_4kz0_core_114 = ~input_a[13];
  assign popcount29_4kz0_core_115 = ~(input_a[18] & input_a[11]);
  assign popcount29_4kz0_core_116 = ~(input_a[22] ^ input_a[24]);
  assign popcount29_4kz0_core_117 = ~input_a[28];
  assign popcount29_4kz0_core_118 = input_a[5] ^ input_a[8];
  assign popcount29_4kz0_core_119 = ~input_a[15];
  assign popcount29_4kz0_core_120 = ~input_a[7];
  assign popcount29_4kz0_core_122 = input_a[24] ^ input_a[12];
  assign popcount29_4kz0_core_124 = ~(input_a[11] | input_a[18]);
  assign popcount29_4kz0_core_125 = ~input_a[17];
  assign popcount29_4kz0_core_126 = ~(input_a[0] | input_a[3]);
  assign popcount29_4kz0_core_127 = input_a[1] & input_a[19];
  assign popcount29_4kz0_core_129 = input_a[6] & input_a[18];
  assign popcount29_4kz0_core_132 = ~(input_a[18] ^ input_a[2]);
  assign popcount29_4kz0_core_133 = ~(input_a[17] & input_a[25]);
  assign popcount29_4kz0_core_134 = ~input_a[26];
  assign popcount29_4kz0_core_135 = ~(input_a[7] & input_a[27]);
  assign popcount29_4kz0_core_136 = ~input_a[14];
  assign popcount29_4kz0_core_137 = input_a[24] | input_a[27];
  assign popcount29_4kz0_core_138 = ~(input_a[22] ^ input_a[13]);
  assign popcount29_4kz0_core_140 = ~(input_a[28] | input_a[23]);
  assign popcount29_4kz0_core_141 = input_a[15] ^ input_a[19];
  assign popcount29_4kz0_core_143 = input_a[2] ^ input_a[8];
  assign popcount29_4kz0_core_144 = ~(input_a[9] | input_a[21]);
  assign popcount29_4kz0_core_145 = ~(input_a[16] | input_a[16]);
  assign popcount29_4kz0_core_146 = ~input_a[27];
  assign popcount29_4kz0_core_147 = input_a[13] & input_a[9];
  assign popcount29_4kz0_core_148 = ~(input_a[5] | input_a[17]);
  assign popcount29_4kz0_core_149 = ~(input_a[24] & input_a[18]);
  assign popcount29_4kz0_core_150 = ~(input_a[8] & input_a[14]);
  assign popcount29_4kz0_core_152 = ~(input_a[11] & input_a[3]);
  assign popcount29_4kz0_core_154 = input_a[26] & input_a[12];
  assign popcount29_4kz0_core_157 = ~(input_a[3] ^ input_a[25]);
  assign popcount29_4kz0_core_158 = ~(input_a[12] ^ input_a[8]);
  assign popcount29_4kz0_core_159 = input_a[11] ^ input_a[10];
  assign popcount29_4kz0_core_162 = ~(input_a[10] ^ input_a[26]);
  assign popcount29_4kz0_core_163 = ~(input_a[2] & input_a[14]);
  assign popcount29_4kz0_core_164 = input_a[25] ^ input_a[7];
  assign popcount29_4kz0_core_166 = ~(input_a[21] ^ input_a[16]);
  assign popcount29_4kz0_core_167 = ~(input_a[17] ^ input_a[25]);
  assign popcount29_4kz0_core_169 = input_a[1] & input_a[1];
  assign popcount29_4kz0_core_171 = ~input_a[0];
  assign popcount29_4kz0_core_176_not = ~input_a[5];
  assign popcount29_4kz0_core_177 = ~(input_a[26] | input_a[13]);
  assign popcount29_4kz0_core_179 = ~(input_a[22] | input_a[15]);
  assign popcount29_4kz0_core_180 = ~(input_a[2] | input_a[2]);
  assign popcount29_4kz0_core_181 = input_a[27] ^ input_a[11];
  assign popcount29_4kz0_core_182 = input_a[13] | input_a[26];
  assign popcount29_4kz0_core_183 = ~(input_a[22] ^ input_a[2]);
  assign popcount29_4kz0_core_184 = input_a[24] | input_a[16];
  assign popcount29_4kz0_core_186 = input_a[25] & input_a[27];
  assign popcount29_4kz0_core_188 = ~input_a[2];
  assign popcount29_4kz0_core_189 = input_a[0] ^ input_a[9];
  assign popcount29_4kz0_core_190 = ~(input_a[28] | input_a[18]);
  assign popcount29_4kz0_core_191 = ~input_a[14];
  assign popcount29_4kz0_core_192 = ~input_a[7];
  assign popcount29_4kz0_core_193 = input_a[26] & input_a[16];
  assign popcount29_4kz0_core_194 = ~(input_a[5] | input_a[21]);
  assign popcount29_4kz0_core_198 = ~(input_a[28] ^ input_a[9]);
  assign popcount29_4kz0_core_199 = ~(input_a[28] ^ input_a[0]);
  assign popcount29_4kz0_core_200 = ~(input_a[5] ^ input_a[27]);
  assign popcount29_4kz0_core_201 = input_a[27] | input_a[4];
  assign popcount29_4kz0_core_202 = ~input_a[4];
  assign popcount29_4kz0_core_205 = ~(input_a[22] & input_a[10]);
  assign popcount29_4kz0_core_206 = input_a[27] ^ input_a[14];
  assign popcount29_4kz0_core_207 = input_a[2] ^ input_a[25];

  assign popcount29_4kz0_out[0] = input_a[11];
  assign popcount29_4kz0_out[1] = 1'b0;
  assign popcount29_4kz0_out[2] = popcount29_4kz0_core_093;
  assign popcount29_4kz0_out[3] = popcount29_4kz0_core_093;
  assign popcount29_4kz0_out[4] = input_a[16];
endmodule