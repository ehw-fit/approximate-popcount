// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.14966
// WCE=15.0
// EP=0.854645%
// Printed PDK parameters:
//  Area=96095897.0
//  Delay=87564232.0
//  Power=4145300.0

module popcount43_364m(input [42:0] input_a, output [5:0] popcount43_364m_out);
  wire popcount43_364m_core_045;
  wire popcount43_364m_core_046;
  wire popcount43_364m_core_047;
  wire popcount43_364m_core_048;
  wire popcount43_364m_core_049;
  wire popcount43_364m_core_050;
  wire popcount43_364m_core_051;
  wire popcount43_364m_core_052;
  wire popcount43_364m_core_054;
  wire popcount43_364m_core_055;
  wire popcount43_364m_core_056;
  wire popcount43_364m_core_057;
  wire popcount43_364m_core_058;
  wire popcount43_364m_core_059;
  wire popcount43_364m_core_060;
  wire popcount43_364m_core_062;
  wire popcount43_364m_core_064;
  wire popcount43_364m_core_065;
  wire popcount43_364m_core_066;
  wire popcount43_364m_core_067;
  wire popcount43_364m_core_068;
  wire popcount43_364m_core_069;
  wire popcount43_364m_core_071;
  wire popcount43_364m_core_074;
  wire popcount43_364m_core_075;
  wire popcount43_364m_core_077;
  wire popcount43_364m_core_078;
  wire popcount43_364m_core_081;
  wire popcount43_364m_core_082;
  wire popcount43_364m_core_086;
  wire popcount43_364m_core_087;
  wire popcount43_364m_core_088;
  wire popcount43_364m_core_089;
  wire popcount43_364m_core_090;
  wire popcount43_364m_core_099;
  wire popcount43_364m_core_100;
  wire popcount43_364m_core_101;
  wire popcount43_364m_core_102;
  wire popcount43_364m_core_103;
  wire popcount43_364m_core_104;
  wire popcount43_364m_core_114;
  wire popcount43_364m_core_115;
  wire popcount43_364m_core_118;
  wire popcount43_364m_core_119;
  wire popcount43_364m_core_120;
  wire popcount43_364m_core_121;
  wire popcount43_364m_core_122;
  wire popcount43_364m_core_123;
  wire popcount43_364m_core_125;
  wire popcount43_364m_core_126;
  wire popcount43_364m_core_127;
  wire popcount43_364m_core_128;
  wire popcount43_364m_core_129;
  wire popcount43_364m_core_130;
  wire popcount43_364m_core_131;
  wire popcount43_364m_core_133;
  wire popcount43_364m_core_135;
  wire popcount43_364m_core_136;
  wire popcount43_364m_core_138;
  wire popcount43_364m_core_139;
  wire popcount43_364m_core_143;
  wire popcount43_364m_core_146;
  wire popcount43_364m_core_147;
  wire popcount43_364m_core_152;
  wire popcount43_364m_core_154_not;
  wire popcount43_364m_core_156;
  wire popcount43_364m_core_157;
  wire popcount43_364m_core_158;
  wire popcount43_364m_core_159;
  wire popcount43_364m_core_160;
  wire popcount43_364m_core_161;
  wire popcount43_364m_core_162;
  wire popcount43_364m_core_163;
  wire popcount43_364m_core_164;
  wire popcount43_364m_core_165;
  wire popcount43_364m_core_166;
  wire popcount43_364m_core_167;
  wire popcount43_364m_core_168;
  wire popcount43_364m_core_169;
  wire popcount43_364m_core_170;
  wire popcount43_364m_core_172;
  wire popcount43_364m_core_174;
  wire popcount43_364m_core_175;
  wire popcount43_364m_core_176_not;
  wire popcount43_364m_core_177;
  wire popcount43_364m_core_178;
  wire popcount43_364m_core_179;
  wire popcount43_364m_core_180;
  wire popcount43_364m_core_181;
  wire popcount43_364m_core_182;
  wire popcount43_364m_core_183;
  wire popcount43_364m_core_185;
  wire popcount43_364m_core_186;
  wire popcount43_364m_core_187;
  wire popcount43_364m_core_188;
  wire popcount43_364m_core_189;
  wire popcount43_364m_core_190;
  wire popcount43_364m_core_191;
  wire popcount43_364m_core_192;
  wire popcount43_364m_core_193;
  wire popcount43_364m_core_194;
  wire popcount43_364m_core_195;
  wire popcount43_364m_core_196;
  wire popcount43_364m_core_197;
  wire popcount43_364m_core_198;
  wire popcount43_364m_core_200;
  wire popcount43_364m_core_205;
  wire popcount43_364m_core_206;
  wire popcount43_364m_core_207;
  wire popcount43_364m_core_208;
  wire popcount43_364m_core_209;
  wire popcount43_364m_core_210;
  wire popcount43_364m_core_211;
  wire popcount43_364m_core_214;
  wire popcount43_364m_core_217;
  wire popcount43_364m_core_219;
  wire popcount43_364m_core_220;
  wire popcount43_364m_core_221;
  wire popcount43_364m_core_222;
  wire popcount43_364m_core_223;
  wire popcount43_364m_core_224;
  wire popcount43_364m_core_225;
  wire popcount43_364m_core_226;
  wire popcount43_364m_core_227;
  wire popcount43_364m_core_228;
  wire popcount43_364m_core_234;
  wire popcount43_364m_core_235;
  wire popcount43_364m_core_236;
  wire popcount43_364m_core_237;
  wire popcount43_364m_core_238;
  wire popcount43_364m_core_239;
  wire popcount43_364m_core_240;
  wire popcount43_364m_core_242;
  wire popcount43_364m_core_243;
  wire popcount43_364m_core_244;
  wire popcount43_364m_core_245;
  wire popcount43_364m_core_246;
  wire popcount43_364m_core_247;
  wire popcount43_364m_core_248;
  wire popcount43_364m_core_252;
  wire popcount43_364m_core_256;
  wire popcount43_364m_core_257;
  wire popcount43_364m_core_258;
  wire popcount43_364m_core_259;
  wire popcount43_364m_core_260;
  wire popcount43_364m_core_261;
  wire popcount43_364m_core_262;
  wire popcount43_364m_core_263;
  wire popcount43_364m_core_264;
  wire popcount43_364m_core_265;
  wire popcount43_364m_core_266;
  wire popcount43_364m_core_267;
  wire popcount43_364m_core_268;
  wire popcount43_364m_core_269;
  wire popcount43_364m_core_274;
  wire popcount43_364m_core_275;
  wire popcount43_364m_core_276;
  wire popcount43_364m_core_277;
  wire popcount43_364m_core_278;
  wire popcount43_364m_core_279;
  wire popcount43_364m_core_280;
  wire popcount43_364m_core_281;
  wire popcount43_364m_core_282;
  wire popcount43_364m_core_283;
  wire popcount43_364m_core_284;
  wire popcount43_364m_core_285;
  wire popcount43_364m_core_286;
  wire popcount43_364m_core_288;
  wire popcount43_364m_core_290;
  wire popcount43_364m_core_294;
  wire popcount43_364m_core_295;
  wire popcount43_364m_core_297;
  wire popcount43_364m_core_299;
  wire popcount43_364m_core_300;
  wire popcount43_364m_core_301;
  wire popcount43_364m_core_302;
  wire popcount43_364m_core_303;
  wire popcount43_364m_core_304;
  wire popcount43_364m_core_305;
  wire popcount43_364m_core_306;
  wire popcount43_364m_core_307;
  wire popcount43_364m_core_308;
  wire popcount43_364m_core_310;
  wire popcount43_364m_core_314;
  wire popcount43_364m_core_316;
  wire popcount43_364m_core_317;
  wire popcount43_364m_core_318;
  wire popcount43_364m_core_319;
  wire popcount43_364m_core_320;
  wire popcount43_364m_core_321;
  wire popcount43_364m_core_322;
  wire popcount43_364m_core_323;
  wire popcount43_364m_core_324;
  wire popcount43_364m_core_325;
  wire popcount43_364m_core_326;
  wire popcount43_364m_core_327;
  wire popcount43_364m_core_328;
  wire popcount43_364m_core_329;
  wire popcount43_364m_core_330;
  wire popcount43_364m_core_331;
  wire popcount43_364m_core_332;
  wire popcount43_364m_core_333;
  wire popcount43_364m_core_334;
  wire popcount43_364m_core_335;
  wire popcount43_364m_core_337;
  wire popcount43_364m_core_339;

  assign popcount43_364m_core_045 = input_a[0] ^ input_a[1];
  assign popcount43_364m_core_046 = input_a[0] & input_a[1];
  assign popcount43_364m_core_047 = input_a[3] ^ input_a[4];
  assign popcount43_364m_core_048 = input_a[3] & input_a[4];
  assign popcount43_364m_core_049 = ~(input_a[32] | input_a[41]);
  assign popcount43_364m_core_050 = input_a[2] & popcount43_364m_core_047;
  assign popcount43_364m_core_051 = popcount43_364m_core_048 ^ popcount43_364m_core_050;
  assign popcount43_364m_core_052 = popcount43_364m_core_048 & popcount43_364m_core_050;
  assign popcount43_364m_core_054 = popcount43_364m_core_045 & input_a[15];
  assign popcount43_364m_core_055 = popcount43_364m_core_046 ^ popcount43_364m_core_051;
  assign popcount43_364m_core_056 = popcount43_364m_core_046 & popcount43_364m_core_051;
  assign popcount43_364m_core_057 = popcount43_364m_core_055 ^ popcount43_364m_core_054;
  assign popcount43_364m_core_058 = popcount43_364m_core_055 & popcount43_364m_core_054;
  assign popcount43_364m_core_059 = popcount43_364m_core_056 | popcount43_364m_core_058;
  assign popcount43_364m_core_060 = popcount43_364m_core_052 ^ popcount43_364m_core_059;
  assign popcount43_364m_core_062 = ~(input_a[41] ^ input_a[13]);
  assign popcount43_364m_core_064 = input_a[8] ^ input_a[9];
  assign popcount43_364m_core_065 = input_a[8] & input_a[9];
  assign popcount43_364m_core_066 = input_a[7] ^ popcount43_364m_core_064;
  assign popcount43_364m_core_067 = input_a[7] & popcount43_364m_core_064;
  assign popcount43_364m_core_068 = popcount43_364m_core_065 ^ popcount43_364m_core_067;
  assign popcount43_364m_core_069 = popcount43_364m_core_065 & popcount43_364m_core_067;
  assign popcount43_364m_core_071 = input_a[14] & popcount43_364m_core_066;
  assign popcount43_364m_core_074 = popcount43_364m_core_068 ^ popcount43_364m_core_071;
  assign popcount43_364m_core_075 = popcount43_364m_core_068 & popcount43_364m_core_071;
  assign popcount43_364m_core_077 = popcount43_364m_core_069 ^ popcount43_364m_core_075;
  assign popcount43_364m_core_078 = ~input_a[42];
  assign popcount43_364m_core_081 = popcount43_364m_core_057 ^ popcount43_364m_core_074;
  assign popcount43_364m_core_082 = popcount43_364m_core_057 & popcount43_364m_core_074;
  assign popcount43_364m_core_086 = popcount43_364m_core_060 ^ popcount43_364m_core_077;
  assign popcount43_364m_core_087 = popcount43_364m_core_060 & popcount43_364m_core_077;
  assign popcount43_364m_core_088 = popcount43_364m_core_086 ^ popcount43_364m_core_082;
  assign popcount43_364m_core_089 = popcount43_364m_core_086 & popcount43_364m_core_082;
  assign popcount43_364m_core_090 = popcount43_364m_core_087 | popcount43_364m_core_089;
  assign popcount43_364m_core_099 = ~(input_a[22] ^ input_a[17]);
  assign popcount43_364m_core_100 = input_a[21] ^ input_a[35];
  assign popcount43_364m_core_101 = ~(input_a[5] & input_a[38]);
  assign popcount43_364m_core_102 = input_a[42] & input_a[31];
  assign popcount43_364m_core_103 = input_a[11] ^ input_a[21];
  assign popcount43_364m_core_104 = input_a[22] | input_a[38];
  assign popcount43_364m_core_114 = input_a[2] & input_a[7];
  assign popcount43_364m_core_115 = ~(input_a[1] | input_a[16]);
  assign popcount43_364m_core_118 = ~input_a[26];
  assign popcount43_364m_core_119 = input_a[20] ^ input_a[20];
  assign popcount43_364m_core_120 = input_a[19] & input_a[20];
  assign popcount43_364m_core_121 = input_a[18] ^ popcount43_364m_core_119;
  assign popcount43_364m_core_122 = input_a[18] & popcount43_364m_core_119;
  assign popcount43_364m_core_123 = popcount43_364m_core_120 ^ popcount43_364m_core_122;
  assign popcount43_364m_core_125 = input_a[22] ^ input_a[31];
  assign popcount43_364m_core_126 = input_a[17] & popcount43_364m_core_121;
  assign popcount43_364m_core_127 = input_a[25] ^ popcount43_364m_core_123;
  assign popcount43_364m_core_128 = input_a[25] & popcount43_364m_core_123;
  assign popcount43_364m_core_129 = popcount43_364m_core_127 ^ popcount43_364m_core_126;
  assign popcount43_364m_core_130 = popcount43_364m_core_127 & popcount43_364m_core_126;
  assign popcount43_364m_core_131 = popcount43_364m_core_128 | popcount43_364m_core_130;
  assign popcount43_364m_core_133 = input_a[36] | input_a[18];
  assign popcount43_364m_core_135 = input_a[30] | input_a[21];
  assign popcount43_364m_core_136 = ~(input_a[8] | input_a[30]);
  assign popcount43_364m_core_138 = input_a[7] & input_a[6];
  assign popcount43_364m_core_139 = ~(input_a[32] & input_a[5]);
  assign popcount43_364m_core_143 = popcount43_364m_core_129 | input_a[5];
  assign popcount43_364m_core_146 = popcount43_364m_core_131 ^ popcount43_364m_core_143;
  assign popcount43_364m_core_147 = popcount43_364m_core_131 & input_a[5];
  assign popcount43_364m_core_152 = input_a[10] | input_a[12];
  assign popcount43_364m_core_154_not = ~input_a[5];
  assign popcount43_364m_core_156 = popcount43_364m_core_081 ^ popcount43_364m_core_139;
  assign popcount43_364m_core_157 = popcount43_364m_core_081 & popcount43_364m_core_139;
  assign popcount43_364m_core_158 = popcount43_364m_core_156 ^ input_a[5];
  assign popcount43_364m_core_159 = popcount43_364m_core_156 & input_a[5];
  assign popcount43_364m_core_160 = popcount43_364m_core_157 | popcount43_364m_core_159;
  assign popcount43_364m_core_161 = popcount43_364m_core_088 ^ popcount43_364m_core_146;
  assign popcount43_364m_core_162 = popcount43_364m_core_088 & popcount43_364m_core_146;
  assign popcount43_364m_core_163 = popcount43_364m_core_161 ^ popcount43_364m_core_160;
  assign popcount43_364m_core_164 = popcount43_364m_core_161 & popcount43_364m_core_160;
  assign popcount43_364m_core_165 = popcount43_364m_core_162 | popcount43_364m_core_164;
  assign popcount43_364m_core_166 = popcount43_364m_core_090 ^ popcount43_364m_core_147;
  assign popcount43_364m_core_167 = popcount43_364m_core_090 & popcount43_364m_core_147;
  assign popcount43_364m_core_168 = popcount43_364m_core_166 ^ popcount43_364m_core_165;
  assign popcount43_364m_core_169 = popcount43_364m_core_166 & popcount43_364m_core_165;
  assign popcount43_364m_core_170 = popcount43_364m_core_167 | popcount43_364m_core_169;
  assign popcount43_364m_core_172 = ~(input_a[6] ^ input_a[12]);
  assign popcount43_364m_core_174 = ~(input_a[12] ^ input_a[25]);
  assign popcount43_364m_core_175 = input_a[14] & input_a[31];
  assign popcount43_364m_core_176_not = ~input_a[9];
  assign popcount43_364m_core_177 = input_a[21] & input_a[22];
  assign popcount43_364m_core_178 = input_a[35] & input_a[25];
  assign popcount43_364m_core_179 = input_a[24] & input_a[16];
  assign popcount43_364m_core_180 = input_a[23] ^ popcount43_364m_core_178;
  assign popcount43_364m_core_181 = input_a[23] & popcount43_364m_core_178;
  assign popcount43_364m_core_182 = popcount43_364m_core_179 ^ popcount43_364m_core_181;
  assign popcount43_364m_core_183 = popcount43_364m_core_179 & popcount43_364m_core_181;
  assign popcount43_364m_core_185 = input_a[4] & popcount43_364m_core_180;
  assign popcount43_364m_core_186 = popcount43_364m_core_177 ^ popcount43_364m_core_182;
  assign popcount43_364m_core_187 = popcount43_364m_core_177 & popcount43_364m_core_182;
  assign popcount43_364m_core_188 = popcount43_364m_core_186 ^ popcount43_364m_core_185;
  assign popcount43_364m_core_189 = popcount43_364m_core_186 & popcount43_364m_core_185;
  assign popcount43_364m_core_190 = popcount43_364m_core_187 | popcount43_364m_core_189;
  assign popcount43_364m_core_191 = popcount43_364m_core_183 | popcount43_364m_core_190;
  assign popcount43_364m_core_192 = input_a[14] | input_a[36];
  assign popcount43_364m_core_193 = input_a[27] ^ input_a[28];
  assign popcount43_364m_core_194 = input_a[27] & input_a[28];
  assign popcount43_364m_core_195 = input_a[37] ^ popcount43_364m_core_193;
  assign popcount43_364m_core_196 = input_a[26] & popcount43_364m_core_193;
  assign popcount43_364m_core_197 = popcount43_364m_core_194 ^ popcount43_364m_core_196;
  assign popcount43_364m_core_198 = popcount43_364m_core_194 & popcount43_364m_core_196;
  assign popcount43_364m_core_200 = input_a[30] & input_a[31];
  assign popcount43_364m_core_205 = input_a[6] ^ input_a[18];
  assign popcount43_364m_core_206 = input_a[21] & input_a[29];
  assign popcount43_364m_core_207 = popcount43_364m_core_197 ^ popcount43_364m_core_200;
  assign popcount43_364m_core_208 = popcount43_364m_core_197 & popcount43_364m_core_200;
  assign popcount43_364m_core_209 = popcount43_364m_core_207 ^ popcount43_364m_core_206;
  assign popcount43_364m_core_210 = popcount43_364m_core_207 & popcount43_364m_core_206;
  assign popcount43_364m_core_211 = popcount43_364m_core_208 | popcount43_364m_core_210;
  assign popcount43_364m_core_214 = popcount43_364m_core_198 ^ popcount43_364m_core_211;
  assign popcount43_364m_core_217 = input_a[23] ^ input_a[37];
  assign popcount43_364m_core_219 = popcount43_364m_core_188 ^ popcount43_364m_core_209;
  assign popcount43_364m_core_220 = popcount43_364m_core_188 & popcount43_364m_core_209;
  assign popcount43_364m_core_221 = popcount43_364m_core_219 ^ input_a[11];
  assign popcount43_364m_core_222 = popcount43_364m_core_219 & input_a[11];
  assign popcount43_364m_core_223 = popcount43_364m_core_220 | popcount43_364m_core_222;
  assign popcount43_364m_core_224 = popcount43_364m_core_191 ^ popcount43_364m_core_214;
  assign popcount43_364m_core_225 = popcount43_364m_core_191 & popcount43_364m_core_214;
  assign popcount43_364m_core_226 = popcount43_364m_core_224 ^ popcount43_364m_core_223;
  assign popcount43_364m_core_227 = popcount43_364m_core_224 & popcount43_364m_core_223;
  assign popcount43_364m_core_228 = popcount43_364m_core_225 | popcount43_364m_core_227;
  assign popcount43_364m_core_234 = input_a[32] | input_a[33];
  assign popcount43_364m_core_235 = input_a[32] & input_a[33];
  assign popcount43_364m_core_236 = ~(input_a[35] & input_a[36]);
  assign popcount43_364m_core_237 = input_a[35] & input_a[36];
  assign popcount43_364m_core_238 = input_a[34] ^ popcount43_364m_core_236;
  assign popcount43_364m_core_239 = input_a[34] & popcount43_364m_core_236;
  assign popcount43_364m_core_240 = popcount43_364m_core_237 ^ popcount43_364m_core_239;
  assign popcount43_364m_core_242 = popcount43_364m_core_234 ^ popcount43_364m_core_238;
  assign popcount43_364m_core_243 = popcount43_364m_core_234 & popcount43_364m_core_238;
  assign popcount43_364m_core_244 = popcount43_364m_core_235 ^ popcount43_364m_core_240;
  assign popcount43_364m_core_245 = popcount43_364m_core_235 & popcount43_364m_core_240;
  assign popcount43_364m_core_246 = popcount43_364m_core_244 ^ popcount43_364m_core_243;
  assign popcount43_364m_core_247 = popcount43_364m_core_244 & popcount43_364m_core_243;
  assign popcount43_364m_core_248 = popcount43_364m_core_245 | popcount43_364m_core_247;
  assign popcount43_364m_core_252 = input_a[10] & input_a[39];
  assign popcount43_364m_core_256 = input_a[5] | input_a[40];
  assign popcount43_364m_core_257 = input_a[41] ^ input_a[42];
  assign popcount43_364m_core_258 = input_a[41] & input_a[42];
  assign popcount43_364m_core_259 = input_a[40] ^ popcount43_364m_core_257;
  assign popcount43_364m_core_260 = input_a[40] & popcount43_364m_core_257;
  assign popcount43_364m_core_261 = popcount43_364m_core_258 ^ popcount43_364m_core_260;
  assign popcount43_364m_core_262 = popcount43_364m_core_258 & input_a[35];
  assign popcount43_364m_core_263 = input_a[37] ^ popcount43_364m_core_259;
  assign popcount43_364m_core_264 = input_a[37] & popcount43_364m_core_259;
  assign popcount43_364m_core_265 = popcount43_364m_core_252 ^ popcount43_364m_core_261;
  assign popcount43_364m_core_266 = popcount43_364m_core_252 & popcount43_364m_core_261;
  assign popcount43_364m_core_267 = popcount43_364m_core_265 ^ popcount43_364m_core_264;
  assign popcount43_364m_core_268 = popcount43_364m_core_265 & popcount43_364m_core_264;
  assign popcount43_364m_core_269 = popcount43_364m_core_266 | popcount43_364m_core_268;
  assign popcount43_364m_core_274 = ~(input_a[20] | input_a[34]);
  assign popcount43_364m_core_275 = popcount43_364m_core_242 | input_a[12];
  assign popcount43_364m_core_276 = popcount43_364m_core_242 & popcount43_364m_core_263;
  assign popcount43_364m_core_277 = popcount43_364m_core_246 ^ popcount43_364m_core_267;
  assign popcount43_364m_core_278 = popcount43_364m_core_246 & popcount43_364m_core_267;
  assign popcount43_364m_core_279 = popcount43_364m_core_277 ^ popcount43_364m_core_276;
  assign popcount43_364m_core_280 = popcount43_364m_core_277 & popcount43_364m_core_276;
  assign popcount43_364m_core_281 = popcount43_364m_core_278 | popcount43_364m_core_280;
  assign popcount43_364m_core_282 = popcount43_364m_core_248 ^ popcount43_364m_core_269;
  assign popcount43_364m_core_283 = popcount43_364m_core_248 & popcount43_364m_core_269;
  assign popcount43_364m_core_284 = popcount43_364m_core_282 ^ popcount43_364m_core_281;
  assign popcount43_364m_core_285 = popcount43_364m_core_282 & popcount43_364m_core_281;
  assign popcount43_364m_core_286 = popcount43_364m_core_283 | popcount43_364m_core_285;
  assign popcount43_364m_core_288 = ~(input_a[9] | input_a[9]);
  assign popcount43_364m_core_290 = ~input_a[1];
  assign popcount43_364m_core_294 = popcount43_364m_core_221 ^ popcount43_364m_core_279;
  assign popcount43_364m_core_295 = popcount43_364m_core_221 & popcount43_364m_core_279;
  assign popcount43_364m_core_297 = input_a[10] & input_a[17];
  assign popcount43_364m_core_299 = popcount43_364m_core_226 ^ popcount43_364m_core_284;
  assign popcount43_364m_core_300 = popcount43_364m_core_226 & popcount43_364m_core_284;
  assign popcount43_364m_core_301 = popcount43_364m_core_299 ^ popcount43_364m_core_295;
  assign popcount43_364m_core_302 = popcount43_364m_core_299 & popcount43_364m_core_295;
  assign popcount43_364m_core_303 = popcount43_364m_core_300 | popcount43_364m_core_302;
  assign popcount43_364m_core_304 = popcount43_364m_core_228 ^ popcount43_364m_core_286;
  assign popcount43_364m_core_305 = popcount43_364m_core_228 & popcount43_364m_core_286;
  assign popcount43_364m_core_306 = popcount43_364m_core_304 ^ popcount43_364m_core_303;
  assign popcount43_364m_core_307 = popcount43_364m_core_304 & popcount43_364m_core_303;
  assign popcount43_364m_core_308 = popcount43_364m_core_305 | popcount43_364m_core_307;
  assign popcount43_364m_core_310 = ~(input_a[17] | input_a[7]);
  assign popcount43_364m_core_314 = ~(input_a[1] ^ input_a[21]);
  assign popcount43_364m_core_316 = popcount43_364m_core_158 ^ popcount43_364m_core_294;
  assign popcount43_364m_core_317 = popcount43_364m_core_158 & popcount43_364m_core_294;
  assign popcount43_364m_core_318 = popcount43_364m_core_316 ^ popcount43_364m_core_154_not;
  assign popcount43_364m_core_319 = popcount43_364m_core_316 & popcount43_364m_core_154_not;
  assign popcount43_364m_core_320 = popcount43_364m_core_317 | popcount43_364m_core_319;
  assign popcount43_364m_core_321 = popcount43_364m_core_163 ^ popcount43_364m_core_301;
  assign popcount43_364m_core_322 = popcount43_364m_core_163 & popcount43_364m_core_301;
  assign popcount43_364m_core_323 = popcount43_364m_core_321 ^ popcount43_364m_core_320;
  assign popcount43_364m_core_324 = popcount43_364m_core_321 & popcount43_364m_core_320;
  assign popcount43_364m_core_325 = popcount43_364m_core_322 | popcount43_364m_core_324;
  assign popcount43_364m_core_326 = popcount43_364m_core_168 ^ popcount43_364m_core_306;
  assign popcount43_364m_core_327 = popcount43_364m_core_168 & popcount43_364m_core_306;
  assign popcount43_364m_core_328 = popcount43_364m_core_326 ^ popcount43_364m_core_325;
  assign popcount43_364m_core_329 = popcount43_364m_core_326 & popcount43_364m_core_325;
  assign popcount43_364m_core_330 = popcount43_364m_core_327 | popcount43_364m_core_329;
  assign popcount43_364m_core_331 = popcount43_364m_core_170 ^ popcount43_364m_core_308;
  assign popcount43_364m_core_332 = popcount43_364m_core_170 & popcount43_364m_core_308;
  assign popcount43_364m_core_333 = popcount43_364m_core_331 ^ popcount43_364m_core_330;
  assign popcount43_364m_core_334 = popcount43_364m_core_331 & popcount43_364m_core_330;
  assign popcount43_364m_core_335 = popcount43_364m_core_332 | popcount43_364m_core_334;
  assign popcount43_364m_core_337 = input_a[31] | input_a[22];
  assign popcount43_364m_core_339 = ~input_a[13];

  assign popcount43_364m_out[0] = input_a[12];
  assign popcount43_364m_out[1] = popcount43_364m_core_318;
  assign popcount43_364m_out[2] = popcount43_364m_core_323;
  assign popcount43_364m_out[3] = popcount43_364m_core_328;
  assign popcount43_364m_out[4] = popcount43_364m_core_333;
  assign popcount43_364m_out[5] = popcount43_364m_core_335;
endmodule