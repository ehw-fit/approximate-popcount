// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.68765
// WCE=9.0
// EP=0.816575%
// Printed PDK parameters:
//  Area=80326893.0
//  Delay=87321224.0
//  Power=4173900.0

module popcount45_hpgt(input [44:0] input_a, output [5:0] popcount45_hpgt_out);
  wire popcount45_hpgt_core_047;
  wire popcount45_hpgt_core_048;
  wire popcount45_hpgt_core_049;
  wire popcount45_hpgt_core_050;
  wire popcount45_hpgt_core_051;
  wire popcount45_hpgt_core_052;
  wire popcount45_hpgt_core_053;
  wire popcount45_hpgt_core_055;
  wire popcount45_hpgt_core_056;
  wire popcount45_hpgt_core_057;
  wire popcount45_hpgt_core_058;
  wire popcount45_hpgt_core_059;
  wire popcount45_hpgt_core_060;
  wire popcount45_hpgt_core_061;
  wire popcount45_hpgt_core_064;
  wire popcount45_hpgt_core_065;
  wire popcount45_hpgt_core_067;
  wire popcount45_hpgt_core_069;
  wire popcount45_hpgt_core_070;
  wire popcount45_hpgt_core_071;
  wire popcount45_hpgt_core_072;
  wire popcount45_hpgt_core_073;
  wire popcount45_hpgt_core_074;
  wire popcount45_hpgt_core_075;
  wire popcount45_hpgt_core_076_not;
  wire popcount45_hpgt_core_078;
  wire popcount45_hpgt_core_079;
  wire popcount45_hpgt_core_080;
  wire popcount45_hpgt_core_081;
  wire popcount45_hpgt_core_082;
  wire popcount45_hpgt_core_084;
  wire popcount45_hpgt_core_087;
  wire popcount45_hpgt_core_088;
  wire popcount45_hpgt_core_089;
  wire popcount45_hpgt_core_090;
  wire popcount45_hpgt_core_091;
  wire popcount45_hpgt_core_092;
  wire popcount45_hpgt_core_093;
  wire popcount45_hpgt_core_094;
  wire popcount45_hpgt_core_095;
  wire popcount45_hpgt_core_096;
  wire popcount45_hpgt_core_097;
  wire popcount45_hpgt_core_098;
  wire popcount45_hpgt_core_099;
  wire popcount45_hpgt_core_101;
  wire popcount45_hpgt_core_104;
  wire popcount45_hpgt_core_105;
  wire popcount45_hpgt_core_106;
  wire popcount45_hpgt_core_109;
  wire popcount45_hpgt_core_112;
  wire popcount45_hpgt_core_113;
  wire popcount45_hpgt_core_114;
  wire popcount45_hpgt_core_115;
  wire popcount45_hpgt_core_116;
  wire popcount45_hpgt_core_118;
  wire popcount45_hpgt_core_119;
  wire popcount45_hpgt_core_120;
  wire popcount45_hpgt_core_121;
  wire popcount45_hpgt_core_123;
  wire popcount45_hpgt_core_124;
  wire popcount45_hpgt_core_125;
  wire popcount45_hpgt_core_126;
  wire popcount45_hpgt_core_128;
  wire popcount45_hpgt_core_129;
  wire popcount45_hpgt_core_130;
  wire popcount45_hpgt_core_131;
  wire popcount45_hpgt_core_132;
  wire popcount45_hpgt_core_133;
  wire popcount45_hpgt_core_134;
  wire popcount45_hpgt_core_135;
  wire popcount45_hpgt_core_137;
  wire popcount45_hpgt_core_140;
  wire popcount45_hpgt_core_141;
  wire popcount45_hpgt_core_142;
  wire popcount45_hpgt_core_143;
  wire popcount45_hpgt_core_145;
  wire popcount45_hpgt_core_146;
  wire popcount45_hpgt_core_147;
  wire popcount45_hpgt_core_150;
  wire popcount45_hpgt_core_151;
  wire popcount45_hpgt_core_154;
  wire popcount45_hpgt_core_156;
  wire popcount45_hpgt_core_157;
  wire popcount45_hpgt_core_160;
  wire popcount45_hpgt_core_161;
  wire popcount45_hpgt_core_163;
  wire popcount45_hpgt_core_164;
  wire popcount45_hpgt_core_165;
  wire popcount45_hpgt_core_166;
  wire popcount45_hpgt_core_167;
  wire popcount45_hpgt_core_168;
  wire popcount45_hpgt_core_169;
  wire popcount45_hpgt_core_170;
  wire popcount45_hpgt_core_171;
  wire popcount45_hpgt_core_172;
  wire popcount45_hpgt_core_173;
  wire popcount45_hpgt_core_174;
  wire popcount45_hpgt_core_176;
  wire popcount45_hpgt_core_177;
  wire popcount45_hpgt_core_178;
  wire popcount45_hpgt_core_179;
  wire popcount45_hpgt_core_180;
  wire popcount45_hpgt_core_181;
  wire popcount45_hpgt_core_183;
  wire popcount45_hpgt_core_185;
  wire popcount45_hpgt_core_186;
  wire popcount45_hpgt_core_187;
  wire popcount45_hpgt_core_188;
  wire popcount45_hpgt_core_190;
  wire popcount45_hpgt_core_191;
  wire popcount45_hpgt_core_194;
  wire popcount45_hpgt_core_195;
  wire popcount45_hpgt_core_196;
  wire popcount45_hpgt_core_198;
  wire popcount45_hpgt_core_201;
  wire popcount45_hpgt_core_202;
  wire popcount45_hpgt_core_203;
  wire popcount45_hpgt_core_204;
  wire popcount45_hpgt_core_205;
  wire popcount45_hpgt_core_206;
  wire popcount45_hpgt_core_208;
  wire popcount45_hpgt_core_209;
  wire popcount45_hpgt_core_211_not;
  wire popcount45_hpgt_core_213;
  wire popcount45_hpgt_core_215;
  wire popcount45_hpgt_core_216;
  wire popcount45_hpgt_core_217;
  wire popcount45_hpgt_core_218;
  wire popcount45_hpgt_core_219;
  wire popcount45_hpgt_core_220;
  wire popcount45_hpgt_core_224;
  wire popcount45_hpgt_core_225;
  wire popcount45_hpgt_core_226;
  wire popcount45_hpgt_core_227;
  wire popcount45_hpgt_core_228;
  wire popcount45_hpgt_core_229;
  wire popcount45_hpgt_core_230;
  wire popcount45_hpgt_core_231;
  wire popcount45_hpgt_core_232;
  wire popcount45_hpgt_core_233;
  wire popcount45_hpgt_core_234;
  wire popcount45_hpgt_core_235;
  wire popcount45_hpgt_core_236;
  wire popcount45_hpgt_core_237;
  wire popcount45_hpgt_core_239;
  wire popcount45_hpgt_core_244;
  wire popcount45_hpgt_core_245;
  wire popcount45_hpgt_core_246;
  wire popcount45_hpgt_core_247;
  wire popcount45_hpgt_core_248;
  wire popcount45_hpgt_core_249;
  wire popcount45_hpgt_core_250;
  wire popcount45_hpgt_core_251;
  wire popcount45_hpgt_core_252;
  wire popcount45_hpgt_core_253;
  wire popcount45_hpgt_core_254;
  wire popcount45_hpgt_core_255;
  wire popcount45_hpgt_core_256;
  wire popcount45_hpgt_core_257;
  wire popcount45_hpgt_core_258;
  wire popcount45_hpgt_core_260;
  wire popcount45_hpgt_core_263;
  wire popcount45_hpgt_core_265;
  wire popcount45_hpgt_core_270;
  wire popcount45_hpgt_core_271;
  wire popcount45_hpgt_core_272;
  wire popcount45_hpgt_core_273;
  wire popcount45_hpgt_core_274_not;
  wire popcount45_hpgt_core_277;
  wire popcount45_hpgt_core_278;
  wire popcount45_hpgt_core_281;
  wire popcount45_hpgt_core_283;
  wire popcount45_hpgt_core_284;
  wire popcount45_hpgt_core_285;
  wire popcount45_hpgt_core_286;
  wire popcount45_hpgt_core_288;
  wire popcount45_hpgt_core_289;
  wire popcount45_hpgt_core_290;
  wire popcount45_hpgt_core_291;
  wire popcount45_hpgt_core_292;
  wire popcount45_hpgt_core_295;
  wire popcount45_hpgt_core_296;
  wire popcount45_hpgt_core_300;
  wire popcount45_hpgt_core_301;
  wire popcount45_hpgt_core_302;
  wire popcount45_hpgt_core_304;
  wire popcount45_hpgt_core_306;
  wire popcount45_hpgt_core_307;
  wire popcount45_hpgt_core_309;
  wire popcount45_hpgt_core_310;
  wire popcount45_hpgt_core_311;
  wire popcount45_hpgt_core_312;
  wire popcount45_hpgt_core_313;
  wire popcount45_hpgt_core_314;
  wire popcount45_hpgt_core_315;
  wire popcount45_hpgt_core_316;
  wire popcount45_hpgt_core_317;
  wire popcount45_hpgt_core_318;
  wire popcount45_hpgt_core_319;
  wire popcount45_hpgt_core_320;
  wire popcount45_hpgt_core_322;
  wire popcount45_hpgt_core_323;
  wire popcount45_hpgt_core_324;
  wire popcount45_hpgt_core_326;
  wire popcount45_hpgt_core_328;
  wire popcount45_hpgt_core_331;
  wire popcount45_hpgt_core_332;
  wire popcount45_hpgt_core_333;
  wire popcount45_hpgt_core_334;
  wire popcount45_hpgt_core_335;
  wire popcount45_hpgt_core_336;
  wire popcount45_hpgt_core_337;
  wire popcount45_hpgt_core_338;
  wire popcount45_hpgt_core_339;
  wire popcount45_hpgt_core_340;
  wire popcount45_hpgt_core_341;
  wire popcount45_hpgt_core_342;
  wire popcount45_hpgt_core_343;
  wire popcount45_hpgt_core_344;
  wire popcount45_hpgt_core_345;
  wire popcount45_hpgt_core_346;
  wire popcount45_hpgt_core_348;
  wire popcount45_hpgt_core_349;
  wire popcount45_hpgt_core_350;
  wire popcount45_hpgt_core_351;
  wire popcount45_hpgt_core_353;
  wire popcount45_hpgt_core_355;
  wire popcount45_hpgt_core_356;

  assign popcount45_hpgt_core_047 = input_a[0] ^ input_a[1];
  assign popcount45_hpgt_core_048 = input_a[0] & input_a[1];
  assign popcount45_hpgt_core_049 = input_a[3] ^ input_a[4];
  assign popcount45_hpgt_core_050 = input_a[3] & input_a[4];
  assign popcount45_hpgt_core_051 = input_a[2] ^ popcount45_hpgt_core_049;
  assign popcount45_hpgt_core_052 = input_a[2] & popcount45_hpgt_core_049;
  assign popcount45_hpgt_core_053 = popcount45_hpgt_core_050 | popcount45_hpgt_core_052;
  assign popcount45_hpgt_core_055 = popcount45_hpgt_core_047 ^ popcount45_hpgt_core_051;
  assign popcount45_hpgt_core_056 = popcount45_hpgt_core_047 & popcount45_hpgt_core_051;
  assign popcount45_hpgt_core_057 = popcount45_hpgt_core_048 ^ popcount45_hpgt_core_053;
  assign popcount45_hpgt_core_058 = popcount45_hpgt_core_048 & popcount45_hpgt_core_053;
  assign popcount45_hpgt_core_059 = popcount45_hpgt_core_057 ^ popcount45_hpgt_core_056;
  assign popcount45_hpgt_core_060 = popcount45_hpgt_core_057 & popcount45_hpgt_core_056;
  assign popcount45_hpgt_core_061 = popcount45_hpgt_core_058 | popcount45_hpgt_core_060;
  assign popcount45_hpgt_core_064 = input_a[20] & input_a[23];
  assign popcount45_hpgt_core_065 = input_a[12] & input_a[7];
  assign popcount45_hpgt_core_067 = ~(input_a[23] | input_a[37]);
  assign popcount45_hpgt_core_069 = ~(input_a[7] & input_a[44]);
  assign popcount45_hpgt_core_070 = input_a[9] ^ input_a[10];
  assign popcount45_hpgt_core_071 = input_a[9] & input_a[10];
  assign popcount45_hpgt_core_072 = input_a[8] ^ popcount45_hpgt_core_070;
  assign popcount45_hpgt_core_073 = input_a[8] & popcount45_hpgt_core_070;
  assign popcount45_hpgt_core_074 = popcount45_hpgt_core_071 | popcount45_hpgt_core_073;
  assign popcount45_hpgt_core_075 = input_a[44] ^ input_a[30];
  assign popcount45_hpgt_core_076_not = ~popcount45_hpgt_core_072;
  assign popcount45_hpgt_core_078 = popcount45_hpgt_core_065 ^ popcount45_hpgt_core_074;
  assign popcount45_hpgt_core_079 = popcount45_hpgt_core_065 & popcount45_hpgt_core_074;
  assign popcount45_hpgt_core_080 = popcount45_hpgt_core_078 ^ popcount45_hpgt_core_072;
  assign popcount45_hpgt_core_081 = popcount45_hpgt_core_078 & popcount45_hpgt_core_072;
  assign popcount45_hpgt_core_082 = popcount45_hpgt_core_079 | popcount45_hpgt_core_081;
  assign popcount45_hpgt_core_084 = ~(input_a[3] & input_a[18]);
  assign popcount45_hpgt_core_087 = input_a[20] | input_a[33];
  assign popcount45_hpgt_core_088 = ~input_a[24];
  assign popcount45_hpgt_core_089 = popcount45_hpgt_core_055 & popcount45_hpgt_core_076_not;
  assign popcount45_hpgt_core_090 = popcount45_hpgt_core_059 ^ popcount45_hpgt_core_080;
  assign popcount45_hpgt_core_091 = popcount45_hpgt_core_059 & popcount45_hpgt_core_080;
  assign popcount45_hpgt_core_092 = popcount45_hpgt_core_090 ^ popcount45_hpgt_core_089;
  assign popcount45_hpgt_core_093 = popcount45_hpgt_core_090 & popcount45_hpgt_core_089;
  assign popcount45_hpgt_core_094 = popcount45_hpgt_core_091 | popcount45_hpgt_core_093;
  assign popcount45_hpgt_core_095 = popcount45_hpgt_core_061 ^ popcount45_hpgt_core_082;
  assign popcount45_hpgt_core_096 = popcount45_hpgt_core_061 & popcount45_hpgt_core_082;
  assign popcount45_hpgt_core_097 = popcount45_hpgt_core_095 ^ popcount45_hpgt_core_094;
  assign popcount45_hpgt_core_098 = popcount45_hpgt_core_095 & popcount45_hpgt_core_094;
  assign popcount45_hpgt_core_099 = popcount45_hpgt_core_096 | popcount45_hpgt_core_098;
  assign popcount45_hpgt_core_101 = input_a[26] & input_a[0];
  assign popcount45_hpgt_core_104 = ~(input_a[17] & input_a[8]);
  assign popcount45_hpgt_core_105 = input_a[2] & input_a[8];
  assign popcount45_hpgt_core_106 = input_a[31] | input_a[10];
  assign popcount45_hpgt_core_109 = ~(input_a[20] | input_a[6]);
  assign popcount45_hpgt_core_112 = input_a[29] | input_a[12];
  assign popcount45_hpgt_core_113 = ~input_a[0];
  assign popcount45_hpgt_core_114 = ~input_a[10];
  assign popcount45_hpgt_core_115 = input_a[23] ^ input_a[4];
  assign popcount45_hpgt_core_116 = input_a[10] & input_a[37];
  assign popcount45_hpgt_core_118 = ~(input_a[35] & input_a[20]);
  assign popcount45_hpgt_core_119 = input_a[21] & input_a[30];
  assign popcount45_hpgt_core_120 = ~(input_a[42] | input_a[6]);
  assign popcount45_hpgt_core_121 = ~(input_a[14] & input_a[26]);
  assign popcount45_hpgt_core_123 = ~(input_a[11] | input_a[0]);
  assign popcount45_hpgt_core_124 = input_a[11] ^ input_a[12];
  assign popcount45_hpgt_core_125 = ~(input_a[13] | input_a[4]);
  assign popcount45_hpgt_core_126 = ~(input_a[17] ^ input_a[26]);
  assign popcount45_hpgt_core_128 = input_a[34] | input_a[32];
  assign popcount45_hpgt_core_129 = ~(input_a[7] | input_a[30]);
  assign popcount45_hpgt_core_130 = ~input_a[12];
  assign popcount45_hpgt_core_131 = ~(input_a[39] & input_a[9]);
  assign popcount45_hpgt_core_132 = input_a[15] & input_a[7];
  assign popcount45_hpgt_core_133 = ~(input_a[13] & input_a[37]);
  assign popcount45_hpgt_core_134 = input_a[37] & input_a[44];
  assign popcount45_hpgt_core_135 = input_a[14] & input_a[19];
  assign popcount45_hpgt_core_137 = ~(input_a[44] & input_a[38]);
  assign popcount45_hpgt_core_140 = ~(input_a[10] & input_a[38]);
  assign popcount45_hpgt_core_141 = ~input_a[25];
  assign popcount45_hpgt_core_142 = input_a[1] & input_a[11];
  assign popcount45_hpgt_core_143 = ~(input_a[11] & input_a[33]);
  assign popcount45_hpgt_core_145 = input_a[1] & input_a[20];
  assign popcount45_hpgt_core_146 = input_a[37] ^ input_a[41];
  assign popcount45_hpgt_core_147 = input_a[37] & input_a[41];
  assign popcount45_hpgt_core_150 = popcount45_hpgt_core_135 ^ popcount45_hpgt_core_147;
  assign popcount45_hpgt_core_151 = popcount45_hpgt_core_135 & popcount45_hpgt_core_147;
  assign popcount45_hpgt_core_154 = ~(input_a[24] ^ input_a[22]);
  assign popcount45_hpgt_core_156 = input_a[32] ^ input_a[35];
  assign popcount45_hpgt_core_157 = ~(input_a[32] | input_a[25]);
  assign popcount45_hpgt_core_160 = ~input_a[18];
  assign popcount45_hpgt_core_161 = ~(input_a[39] ^ input_a[27]);
  assign popcount45_hpgt_core_163 = ~(input_a[37] | input_a[6]);
  assign popcount45_hpgt_core_164 = input_a[38] & popcount45_hpgt_core_146;
  assign popcount45_hpgt_core_165 = popcount45_hpgt_core_092 ^ popcount45_hpgt_core_150;
  assign popcount45_hpgt_core_166 = popcount45_hpgt_core_092 & popcount45_hpgt_core_150;
  assign popcount45_hpgt_core_167 = popcount45_hpgt_core_165 ^ popcount45_hpgt_core_164;
  assign popcount45_hpgt_core_168 = popcount45_hpgt_core_165 & popcount45_hpgt_core_164;
  assign popcount45_hpgt_core_169 = popcount45_hpgt_core_166 | popcount45_hpgt_core_168;
  assign popcount45_hpgt_core_170 = popcount45_hpgt_core_097 ^ popcount45_hpgt_core_151;
  assign popcount45_hpgt_core_171 = popcount45_hpgt_core_097 & popcount45_hpgt_core_151;
  assign popcount45_hpgt_core_172 = popcount45_hpgt_core_170 ^ popcount45_hpgt_core_169;
  assign popcount45_hpgt_core_173 = popcount45_hpgt_core_170 & popcount45_hpgt_core_169;
  assign popcount45_hpgt_core_174 = popcount45_hpgt_core_171 | popcount45_hpgt_core_173;
  assign popcount45_hpgt_core_176 = ~(input_a[14] & input_a[20]);
  assign popcount45_hpgt_core_177 = popcount45_hpgt_core_099 | popcount45_hpgt_core_174;
  assign popcount45_hpgt_core_178 = input_a[2] ^ input_a[17];
  assign popcount45_hpgt_core_179 = input_a[20] & input_a[1];
  assign popcount45_hpgt_core_180 = input_a[41] | input_a[43];
  assign popcount45_hpgt_core_181 = ~input_a[38];
  assign popcount45_hpgt_core_183 = input_a[35] | input_a[10];
  assign popcount45_hpgt_core_185 = input_a[25] ^ input_a[26];
  assign popcount45_hpgt_core_186 = input_a[22] & input_a[5];
  assign popcount45_hpgt_core_187 = ~(input_a[43] ^ input_a[29]);
  assign popcount45_hpgt_core_188 = input_a[25] & input_a[20];
  assign popcount45_hpgt_core_190 = input_a[43] & input_a[34];
  assign popcount45_hpgt_core_191 = popcount45_hpgt_core_188 | popcount45_hpgt_core_190;
  assign popcount45_hpgt_core_194 = ~(input_a[38] | input_a[7]);
  assign popcount45_hpgt_core_195 = popcount45_hpgt_core_186 ^ popcount45_hpgt_core_191;
  assign popcount45_hpgt_core_196 = popcount45_hpgt_core_186 & popcount45_hpgt_core_191;
  assign popcount45_hpgt_core_198 = input_a[16] ^ input_a[29];
  assign popcount45_hpgt_core_201 = ~(input_a[7] ^ input_a[31]);
  assign popcount45_hpgt_core_202 = input_a[28] | input_a[29];
  assign popcount45_hpgt_core_203 = input_a[28] & input_a[29];
  assign popcount45_hpgt_core_204 = input_a[44] & input_a[4];
  assign popcount45_hpgt_core_205 = input_a[27] & popcount45_hpgt_core_202;
  assign popcount45_hpgt_core_206 = popcount45_hpgt_core_203 | popcount45_hpgt_core_205;
  assign popcount45_hpgt_core_208 = input_a[5] | input_a[15];
  assign popcount45_hpgt_core_209 = input_a[11] & input_a[26];
  assign popcount45_hpgt_core_211_not = ~input_a[32];
  assign popcount45_hpgt_core_213 = ~(input_a[30] & input_a[40]);
  assign popcount45_hpgt_core_215 = input_a[6] & input_a[40];
  assign popcount45_hpgt_core_216 = popcount45_hpgt_core_206 ^ popcount45_hpgt_core_209;
  assign popcount45_hpgt_core_217 = popcount45_hpgt_core_206 & popcount45_hpgt_core_209;
  assign popcount45_hpgt_core_218 = popcount45_hpgt_core_216 ^ popcount45_hpgt_core_215;
  assign popcount45_hpgt_core_219 = popcount45_hpgt_core_216 & popcount45_hpgt_core_215;
  assign popcount45_hpgt_core_220 = popcount45_hpgt_core_217 | popcount45_hpgt_core_219;
  assign popcount45_hpgt_core_224 = ~(input_a[44] ^ input_a[41]);
  assign popcount45_hpgt_core_225 = ~(input_a[30] ^ input_a[28]);
  assign popcount45_hpgt_core_226 = input_a[23] & input_a[24];
  assign popcount45_hpgt_core_227 = input_a[18] & input_a[13];
  assign popcount45_hpgt_core_228 = popcount45_hpgt_core_195 ^ popcount45_hpgt_core_218;
  assign popcount45_hpgt_core_229 = popcount45_hpgt_core_195 & popcount45_hpgt_core_218;
  assign popcount45_hpgt_core_230 = popcount45_hpgt_core_228 ^ popcount45_hpgt_core_227;
  assign popcount45_hpgt_core_231 = popcount45_hpgt_core_228 & popcount45_hpgt_core_227;
  assign popcount45_hpgt_core_232 = popcount45_hpgt_core_229 | popcount45_hpgt_core_231;
  assign popcount45_hpgt_core_233 = popcount45_hpgt_core_196 ^ popcount45_hpgt_core_220;
  assign popcount45_hpgt_core_234 = popcount45_hpgt_core_196 & popcount45_hpgt_core_220;
  assign popcount45_hpgt_core_235 = popcount45_hpgt_core_233 ^ popcount45_hpgt_core_232;
  assign popcount45_hpgt_core_236 = popcount45_hpgt_core_233 & popcount45_hpgt_core_232;
  assign popcount45_hpgt_core_237 = popcount45_hpgt_core_234 | popcount45_hpgt_core_236;
  assign popcount45_hpgt_core_239 = ~(input_a[32] & input_a[14]);
  assign popcount45_hpgt_core_244 = input_a[33] & input_a[21];
  assign popcount45_hpgt_core_245 = ~(input_a[18] & input_a[41]);
  assign popcount45_hpgt_core_246 = input_a[24] & input_a[30];
  assign popcount45_hpgt_core_247 = popcount45_hpgt_core_244 | popcount45_hpgt_core_246;
  assign popcount45_hpgt_core_248 = ~(input_a[10] & input_a[35]);
  assign popcount45_hpgt_core_249 = ~(input_a[35] & input_a[31]);
  assign popcount45_hpgt_core_250 = input_a[42] & input_a[31];
  assign popcount45_hpgt_core_251 = input_a[15] | input_a[31];
  assign popcount45_hpgt_core_252 = input_a[15] & input_a[36];
  assign popcount45_hpgt_core_253 = popcount45_hpgt_core_250 | popcount45_hpgt_core_252;
  assign popcount45_hpgt_core_254 = ~(input_a[5] | input_a[25]);
  assign popcount45_hpgt_core_255 = input_a[30] & input_a[11];
  assign popcount45_hpgt_core_256 = input_a[5] ^ input_a[22];
  assign popcount45_hpgt_core_257 = popcount45_hpgt_core_247 ^ popcount45_hpgt_core_253;
  assign popcount45_hpgt_core_258 = popcount45_hpgt_core_247 & popcount45_hpgt_core_253;
  assign popcount45_hpgt_core_260 = input_a[26] & input_a[38];
  assign popcount45_hpgt_core_263 = ~(input_a[12] ^ input_a[43]);
  assign popcount45_hpgt_core_265 = input_a[19] | input_a[16];
  assign popcount45_hpgt_core_270 = ~(input_a[23] | input_a[2]);
  assign popcount45_hpgt_core_271 = input_a[11] ^ input_a[44];
  assign popcount45_hpgt_core_272 = ~input_a[43];
  assign popcount45_hpgt_core_273 = input_a[41] ^ input_a[19];
  assign popcount45_hpgt_core_274_not = ~input_a[37];
  assign popcount45_hpgt_core_277 = ~(input_a[17] & input_a[22]);
  assign popcount45_hpgt_core_278 = input_a[22] | input_a[24];
  assign popcount45_hpgt_core_281 = ~input_a[25];
  assign popcount45_hpgt_core_283 = ~input_a[7];
  assign popcount45_hpgt_core_284 = ~input_a[38];
  assign popcount45_hpgt_core_285 = input_a[25] & input_a[40];
  assign popcount45_hpgt_core_286 = ~(input_a[36] ^ input_a[8]);
  assign popcount45_hpgt_core_288 = ~(input_a[35] | input_a[39]);
  assign popcount45_hpgt_core_289 = input_a[0] ^ input_a[40];
  assign popcount45_hpgt_core_290 = ~(input_a[8] | input_a[8]);
  assign popcount45_hpgt_core_291 = ~(input_a[16] ^ input_a[3]);
  assign popcount45_hpgt_core_292 = input_a[35] & input_a[17];
  assign popcount45_hpgt_core_295 = popcount45_hpgt_core_257 ^ popcount45_hpgt_core_292;
  assign popcount45_hpgt_core_296 = popcount45_hpgt_core_257 & popcount45_hpgt_core_292;
  assign popcount45_hpgt_core_300 = popcount45_hpgt_core_258 | popcount45_hpgt_core_296;
  assign popcount45_hpgt_core_301 = ~input_a[5];
  assign popcount45_hpgt_core_302 = input_a[8] & input_a[11];
  assign popcount45_hpgt_core_304 = input_a[18] ^ input_a[36];
  assign popcount45_hpgt_core_306 = ~(input_a[38] & input_a[41]);
  assign popcount45_hpgt_core_307 = ~(input_a[32] | input_a[29]);
  assign popcount45_hpgt_core_309 = input_a[32] & input_a[39];
  assign popcount45_hpgt_core_310 = popcount45_hpgt_core_230 ^ popcount45_hpgt_core_295;
  assign popcount45_hpgt_core_311 = popcount45_hpgt_core_230 & popcount45_hpgt_core_295;
  assign popcount45_hpgt_core_312 = popcount45_hpgt_core_310 ^ popcount45_hpgt_core_309;
  assign popcount45_hpgt_core_313 = popcount45_hpgt_core_310 & popcount45_hpgt_core_309;
  assign popcount45_hpgt_core_314 = popcount45_hpgt_core_311 | popcount45_hpgt_core_313;
  assign popcount45_hpgt_core_315 = popcount45_hpgt_core_235 ^ popcount45_hpgt_core_300;
  assign popcount45_hpgt_core_316 = popcount45_hpgt_core_235 & popcount45_hpgt_core_300;
  assign popcount45_hpgt_core_317 = popcount45_hpgt_core_315 ^ popcount45_hpgt_core_314;
  assign popcount45_hpgt_core_318 = popcount45_hpgt_core_315 & popcount45_hpgt_core_314;
  assign popcount45_hpgt_core_319 = popcount45_hpgt_core_316 | popcount45_hpgt_core_318;
  assign popcount45_hpgt_core_320 = ~popcount45_hpgt_core_237;
  assign popcount45_hpgt_core_322 = popcount45_hpgt_core_320 ^ popcount45_hpgt_core_319;
  assign popcount45_hpgt_core_323 = popcount45_hpgt_core_320 & popcount45_hpgt_core_319;
  assign popcount45_hpgt_core_324 = popcount45_hpgt_core_237 | popcount45_hpgt_core_323;
  assign popcount45_hpgt_core_326 = input_a[24] | input_a[3];
  assign popcount45_hpgt_core_328 = ~(input_a[20] ^ input_a[25]);
  assign popcount45_hpgt_core_331 = input_a[16] & input_a[44];
  assign popcount45_hpgt_core_332 = popcount45_hpgt_core_167 ^ popcount45_hpgt_core_312;
  assign popcount45_hpgt_core_333 = popcount45_hpgt_core_167 & popcount45_hpgt_core_312;
  assign popcount45_hpgt_core_334 = popcount45_hpgt_core_332 ^ popcount45_hpgt_core_331;
  assign popcount45_hpgt_core_335 = popcount45_hpgt_core_332 & popcount45_hpgt_core_331;
  assign popcount45_hpgt_core_336 = popcount45_hpgt_core_333 | popcount45_hpgt_core_335;
  assign popcount45_hpgt_core_337 = popcount45_hpgt_core_172 ^ popcount45_hpgt_core_317;
  assign popcount45_hpgt_core_338 = popcount45_hpgt_core_172 & popcount45_hpgt_core_317;
  assign popcount45_hpgt_core_339 = popcount45_hpgt_core_337 ^ popcount45_hpgt_core_336;
  assign popcount45_hpgt_core_340 = popcount45_hpgt_core_337 & popcount45_hpgt_core_336;
  assign popcount45_hpgt_core_341 = popcount45_hpgt_core_338 | popcount45_hpgt_core_340;
  assign popcount45_hpgt_core_342 = popcount45_hpgt_core_177 ^ popcount45_hpgt_core_322;
  assign popcount45_hpgt_core_343 = popcount45_hpgt_core_177 & popcount45_hpgt_core_322;
  assign popcount45_hpgt_core_344 = popcount45_hpgt_core_342 ^ popcount45_hpgt_core_341;
  assign popcount45_hpgt_core_345 = popcount45_hpgt_core_342 & popcount45_hpgt_core_341;
  assign popcount45_hpgt_core_346 = popcount45_hpgt_core_343 | popcount45_hpgt_core_345;
  assign popcount45_hpgt_core_348 = input_a[37] & input_a[18];
  assign popcount45_hpgt_core_349 = popcount45_hpgt_core_324 ^ popcount45_hpgt_core_346;
  assign popcount45_hpgt_core_350 = popcount45_hpgt_core_324 & popcount45_hpgt_core_346;
  assign popcount45_hpgt_core_351 = ~input_a[36];
  assign popcount45_hpgt_core_353 = ~(input_a[8] | input_a[10]);
  assign popcount45_hpgt_core_355 = input_a[6] ^ input_a[35];
  assign popcount45_hpgt_core_356 = input_a[33] | input_a[8];

  assign popcount45_hpgt_out[0] = input_a[23];
  assign popcount45_hpgt_out[1] = popcount45_hpgt_core_334;
  assign popcount45_hpgt_out[2] = popcount45_hpgt_core_339;
  assign popcount45_hpgt_out[3] = popcount45_hpgt_core_344;
  assign popcount45_hpgt_out[4] = popcount45_hpgt_core_349;
  assign popcount45_hpgt_out[5] = popcount45_hpgt_core_350;
endmodule