// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.64904
// WCE=19.0
// EP=0.955523%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_vbgj(input [27:0] input_a, output [4:0] popcount28_vbgj_out);
  wire popcount28_vbgj_core_032;
  wire popcount28_vbgj_core_034;
  wire popcount28_vbgj_core_035;
  wire popcount28_vbgj_core_036;
  wire popcount28_vbgj_core_037;
  wire popcount28_vbgj_core_038;
  wire popcount28_vbgj_core_039_not;
  wire popcount28_vbgj_core_041;
  wire popcount28_vbgj_core_042;
  wire popcount28_vbgj_core_043;
  wire popcount28_vbgj_core_049;
  wire popcount28_vbgj_core_050;
  wire popcount28_vbgj_core_052;
  wire popcount28_vbgj_core_054;
  wire popcount28_vbgj_core_055;
  wire popcount28_vbgj_core_057;
  wire popcount28_vbgj_core_058;
  wire popcount28_vbgj_core_061;
  wire popcount28_vbgj_core_063;
  wire popcount28_vbgj_core_065;
  wire popcount28_vbgj_core_069;
  wire popcount28_vbgj_core_070;
  wire popcount28_vbgj_core_072;
  wire popcount28_vbgj_core_073;
  wire popcount28_vbgj_core_074;
  wire popcount28_vbgj_core_075;
  wire popcount28_vbgj_core_076;
  wire popcount28_vbgj_core_077;
  wire popcount28_vbgj_core_078;
  wire popcount28_vbgj_core_079;
  wire popcount28_vbgj_core_081;
  wire popcount28_vbgj_core_082;
  wire popcount28_vbgj_core_083;
  wire popcount28_vbgj_core_084;
  wire popcount28_vbgj_core_085;
  wire popcount28_vbgj_core_086;
  wire popcount28_vbgj_core_087;
  wire popcount28_vbgj_core_088;
  wire popcount28_vbgj_core_090;
  wire popcount28_vbgj_core_091;
  wire popcount28_vbgj_core_092;
  wire popcount28_vbgj_core_093;
  wire popcount28_vbgj_core_095;
  wire popcount28_vbgj_core_096;
  wire popcount28_vbgj_core_097;
  wire popcount28_vbgj_core_098;
  wire popcount28_vbgj_core_099;
  wire popcount28_vbgj_core_101;
  wire popcount28_vbgj_core_102;
  wire popcount28_vbgj_core_104;
  wire popcount28_vbgj_core_105;
  wire popcount28_vbgj_core_106;
  wire popcount28_vbgj_core_107;
  wire popcount28_vbgj_core_109;
  wire popcount28_vbgj_core_112;
  wire popcount28_vbgj_core_113;
  wire popcount28_vbgj_core_114;
  wire popcount28_vbgj_core_115;
  wire popcount28_vbgj_core_116;
  wire popcount28_vbgj_core_117;
  wire popcount28_vbgj_core_118;
  wire popcount28_vbgj_core_119;
  wire popcount28_vbgj_core_120;
  wire popcount28_vbgj_core_122;
  wire popcount28_vbgj_core_124;
  wire popcount28_vbgj_core_125_not;
  wire popcount28_vbgj_core_126;
  wire popcount28_vbgj_core_127;
  wire popcount28_vbgj_core_131;
  wire popcount28_vbgj_core_132_not;
  wire popcount28_vbgj_core_133;
  wire popcount28_vbgj_core_134;
  wire popcount28_vbgj_core_136;
  wire popcount28_vbgj_core_137;
  wire popcount28_vbgj_core_138;
  wire popcount28_vbgj_core_142;
  wire popcount28_vbgj_core_145;
  wire popcount28_vbgj_core_146;
  wire popcount28_vbgj_core_147;
  wire popcount28_vbgj_core_148;
  wire popcount28_vbgj_core_149;
  wire popcount28_vbgj_core_151;
  wire popcount28_vbgj_core_154;
  wire popcount28_vbgj_core_157;
  wire popcount28_vbgj_core_158;
  wire popcount28_vbgj_core_160;
  wire popcount28_vbgj_core_166;
  wire popcount28_vbgj_core_168;
  wire popcount28_vbgj_core_169;
  wire popcount28_vbgj_core_173;
  wire popcount28_vbgj_core_174;
  wire popcount28_vbgj_core_177;
  wire popcount28_vbgj_core_178;
  wire popcount28_vbgj_core_180;
  wire popcount28_vbgj_core_181;
  wire popcount28_vbgj_core_182;
  wire popcount28_vbgj_core_183;
  wire popcount28_vbgj_core_184;
  wire popcount28_vbgj_core_185;
  wire popcount28_vbgj_core_187_not;
  wire popcount28_vbgj_core_191;
  wire popcount28_vbgj_core_193;
  wire popcount28_vbgj_core_194;
  wire popcount28_vbgj_core_196;
  wire popcount28_vbgj_core_199;
  wire popcount28_vbgj_core_200;
  wire popcount28_vbgj_core_201;

  assign popcount28_vbgj_core_032 = input_a[22] | input_a[4];
  assign popcount28_vbgj_core_034 = ~input_a[9];
  assign popcount28_vbgj_core_035 = input_a[19] ^ input_a[2];
  assign popcount28_vbgj_core_036 = ~input_a[27];
  assign popcount28_vbgj_core_037 = ~(input_a[14] & input_a[9]);
  assign popcount28_vbgj_core_038 = input_a[4] ^ input_a[12];
  assign popcount28_vbgj_core_039_not = ~input_a[26];
  assign popcount28_vbgj_core_041 = input_a[27] ^ input_a[6];
  assign popcount28_vbgj_core_042 = input_a[9] ^ input_a[1];
  assign popcount28_vbgj_core_043 = input_a[3] ^ input_a[18];
  assign popcount28_vbgj_core_049 = ~input_a[13];
  assign popcount28_vbgj_core_050 = ~(input_a[1] | input_a[8]);
  assign popcount28_vbgj_core_052 = input_a[2] | input_a[22];
  assign popcount28_vbgj_core_054 = ~(input_a[3] | input_a[4]);
  assign popcount28_vbgj_core_055 = ~input_a[3];
  assign popcount28_vbgj_core_057 = input_a[2] ^ input_a[0];
  assign popcount28_vbgj_core_058 = ~(input_a[21] ^ input_a[18]);
  assign popcount28_vbgj_core_061 = input_a[13] ^ input_a[14];
  assign popcount28_vbgj_core_063 = ~input_a[13];
  assign popcount28_vbgj_core_065 = ~(input_a[12] ^ input_a[27]);
  assign popcount28_vbgj_core_069 = ~input_a[22];
  assign popcount28_vbgj_core_070 = ~input_a[4];
  assign popcount28_vbgj_core_072 = ~(input_a[3] | input_a[0]);
  assign popcount28_vbgj_core_073 = ~(input_a[2] | input_a[20]);
  assign popcount28_vbgj_core_074 = input_a[16] | input_a[21];
  assign popcount28_vbgj_core_075 = ~input_a[12];
  assign popcount28_vbgj_core_076 = ~(input_a[27] & input_a[4]);
  assign popcount28_vbgj_core_077 = ~(input_a[21] & input_a[8]);
  assign popcount28_vbgj_core_078 = ~input_a[15];
  assign popcount28_vbgj_core_079 = input_a[19] ^ input_a[11];
  assign popcount28_vbgj_core_081 = input_a[2] ^ input_a[20];
  assign popcount28_vbgj_core_082 = input_a[19] & input_a[0];
  assign popcount28_vbgj_core_083 = ~input_a[9];
  assign popcount28_vbgj_core_084 = input_a[18] | input_a[0];
  assign popcount28_vbgj_core_085 = ~(input_a[9] ^ input_a[7]);
  assign popcount28_vbgj_core_086 = ~(input_a[17] ^ input_a[21]);
  assign popcount28_vbgj_core_087 = input_a[11] | input_a[4];
  assign popcount28_vbgj_core_088 = ~(input_a[27] & input_a[8]);
  assign popcount28_vbgj_core_090 = input_a[5] | input_a[0];
  assign popcount28_vbgj_core_091 = input_a[14] & input_a[22];
  assign popcount28_vbgj_core_092 = ~(input_a[9] & input_a[19]);
  assign popcount28_vbgj_core_093 = input_a[25] & input_a[27];
  assign popcount28_vbgj_core_095 = input_a[24] ^ input_a[4];
  assign popcount28_vbgj_core_096 = input_a[9] | input_a[4];
  assign popcount28_vbgj_core_097 = ~input_a[4];
  assign popcount28_vbgj_core_098 = input_a[8] ^ input_a[13];
  assign popcount28_vbgj_core_099 = ~(input_a[0] ^ input_a[3]);
  assign popcount28_vbgj_core_101 = input_a[26] ^ input_a[10];
  assign popcount28_vbgj_core_102 = input_a[5] ^ input_a[1];
  assign popcount28_vbgj_core_104 = input_a[11] ^ input_a[22];
  assign popcount28_vbgj_core_105 = ~input_a[9];
  assign popcount28_vbgj_core_106 = input_a[14] ^ input_a[10];
  assign popcount28_vbgj_core_107 = ~(input_a[15] ^ input_a[2]);
  assign popcount28_vbgj_core_109 = ~(input_a[10] | input_a[15]);
  assign popcount28_vbgj_core_112 = ~(input_a[26] ^ input_a[7]);
  assign popcount28_vbgj_core_113 = ~input_a[18];
  assign popcount28_vbgj_core_114 = ~(input_a[23] ^ input_a[20]);
  assign popcount28_vbgj_core_115 = input_a[0] ^ input_a[11];
  assign popcount28_vbgj_core_116 = ~input_a[9];
  assign popcount28_vbgj_core_117 = ~input_a[19];
  assign popcount28_vbgj_core_118 = ~(input_a[9] | input_a[2]);
  assign popcount28_vbgj_core_119 = input_a[13] ^ input_a[8];
  assign popcount28_vbgj_core_120 = ~(input_a[26] & input_a[19]);
  assign popcount28_vbgj_core_122 = input_a[23] ^ input_a[4];
  assign popcount28_vbgj_core_124 = ~(input_a[12] | input_a[15]);
  assign popcount28_vbgj_core_125_not = ~input_a[23];
  assign popcount28_vbgj_core_126 = ~(input_a[0] | input_a[12]);
  assign popcount28_vbgj_core_127 = input_a[20] | input_a[20];
  assign popcount28_vbgj_core_131 = input_a[11] & input_a[20];
  assign popcount28_vbgj_core_132_not = ~input_a[7];
  assign popcount28_vbgj_core_133 = input_a[19] ^ input_a[17];
  assign popcount28_vbgj_core_134 = input_a[13] & input_a[8];
  assign popcount28_vbgj_core_136 = input_a[17] & input_a[6];
  assign popcount28_vbgj_core_137 = ~(input_a[0] & input_a[16]);
  assign popcount28_vbgj_core_138 = input_a[0] & input_a[9];
  assign popcount28_vbgj_core_142 = input_a[2] ^ input_a[5];
  assign popcount28_vbgj_core_145 = ~input_a[9];
  assign popcount28_vbgj_core_146 = ~(input_a[14] ^ input_a[17]);
  assign popcount28_vbgj_core_147 = ~input_a[26];
  assign popcount28_vbgj_core_148 = ~(input_a[15] & input_a[9]);
  assign popcount28_vbgj_core_149 = ~(input_a[21] ^ input_a[27]);
  assign popcount28_vbgj_core_151 = ~input_a[11];
  assign popcount28_vbgj_core_154 = input_a[10] | input_a[27];
  assign popcount28_vbgj_core_157 = ~input_a[3];
  assign popcount28_vbgj_core_158 = input_a[7] & input_a[12];
  assign popcount28_vbgj_core_160 = input_a[15] ^ input_a[11];
  assign popcount28_vbgj_core_166 = input_a[27] | input_a[6];
  assign popcount28_vbgj_core_168 = ~(input_a[7] ^ input_a[1]);
  assign popcount28_vbgj_core_169 = ~(input_a[11] | input_a[5]);
  assign popcount28_vbgj_core_173 = input_a[17] & input_a[3];
  assign popcount28_vbgj_core_174 = ~(input_a[11] & input_a[0]);
  assign popcount28_vbgj_core_177 = input_a[20] ^ input_a[6];
  assign popcount28_vbgj_core_178 = ~input_a[23];
  assign popcount28_vbgj_core_180 = input_a[0] | input_a[4];
  assign popcount28_vbgj_core_181 = input_a[8] & input_a[12];
  assign popcount28_vbgj_core_182 = input_a[12] & input_a[10];
  assign popcount28_vbgj_core_183 = input_a[10] & input_a[19];
  assign popcount28_vbgj_core_184 = ~(input_a[22] | input_a[2]);
  assign popcount28_vbgj_core_185 = ~(input_a[2] | input_a[18]);
  assign popcount28_vbgj_core_187_not = ~input_a[6];
  assign popcount28_vbgj_core_191 = ~(input_a[20] ^ input_a[5]);
  assign popcount28_vbgj_core_193 = input_a[2] | input_a[0];
  assign popcount28_vbgj_core_194 = input_a[22] ^ input_a[7];
  assign popcount28_vbgj_core_196 = ~(input_a[11] ^ input_a[10]);
  assign popcount28_vbgj_core_199 = ~(input_a[14] & input_a[0]);
  assign popcount28_vbgj_core_200 = input_a[12] & input_a[14];
  assign popcount28_vbgj_core_201 = input_a[7] & input_a[10];

  assign popcount28_vbgj_out[0] = input_a[13];
  assign popcount28_vbgj_out[1] = 1'b0;
  assign popcount28_vbgj_out[2] = input_a[19];
  assign popcount28_vbgj_out[3] = 1'b0;
  assign popcount28_vbgj_out[4] = 1'b1;
endmodule