// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.4559
// WCE=16.0
// EP=0.873594%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_96cy(input [29:0] input_a, output [4:0] popcount30_96cy_out);
  wire popcount30_96cy_core_032;
  wire popcount30_96cy_core_033;
  wire popcount30_96cy_core_034;
  wire popcount30_96cy_core_035;
  wire popcount30_96cy_core_036;
  wire popcount30_96cy_core_038;
  wire popcount30_96cy_core_041;
  wire popcount30_96cy_core_043;
  wire popcount30_96cy_core_044;
  wire popcount30_96cy_core_045;
  wire popcount30_96cy_core_046;
  wire popcount30_96cy_core_048;
  wire popcount30_96cy_core_049;
  wire popcount30_96cy_core_050;
  wire popcount30_96cy_core_051;
  wire popcount30_96cy_core_053;
  wire popcount30_96cy_core_054;
  wire popcount30_96cy_core_058;
  wire popcount30_96cy_core_061;
  wire popcount30_96cy_core_065;
  wire popcount30_96cy_core_068;
  wire popcount30_96cy_core_069;
  wire popcount30_96cy_core_070;
  wire popcount30_96cy_core_071;
  wire popcount30_96cy_core_072;
  wire popcount30_96cy_core_073;
  wire popcount30_96cy_core_074;
  wire popcount30_96cy_core_075;
  wire popcount30_96cy_core_078;
  wire popcount30_96cy_core_079;
  wire popcount30_96cy_core_080;
  wire popcount30_96cy_core_090;
  wire popcount30_96cy_core_093;
  wire popcount30_96cy_core_094;
  wire popcount30_96cy_core_096;
  wire popcount30_96cy_core_097;
  wire popcount30_96cy_core_098;
  wire popcount30_96cy_core_102;
  wire popcount30_96cy_core_105;
  wire popcount30_96cy_core_106;
  wire popcount30_96cy_core_109;
  wire popcount30_96cy_core_110;
  wire popcount30_96cy_core_111;
  wire popcount30_96cy_core_112;
  wire popcount30_96cy_core_114;
  wire popcount30_96cy_core_115;
  wire popcount30_96cy_core_116;
  wire popcount30_96cy_core_118;
  wire popcount30_96cy_core_119;
  wire popcount30_96cy_core_121;
  wire popcount30_96cy_core_122_not;
  wire popcount30_96cy_core_123;
  wire popcount30_96cy_core_124;
  wire popcount30_96cy_core_125;
  wire popcount30_96cy_core_126;
  wire popcount30_96cy_core_128;
  wire popcount30_96cy_core_129;
  wire popcount30_96cy_core_130;
  wire popcount30_96cy_core_131;
  wire popcount30_96cy_core_132;
  wire popcount30_96cy_core_133;
  wire popcount30_96cy_core_136;
  wire popcount30_96cy_core_139;
  wire popcount30_96cy_core_140;
  wire popcount30_96cy_core_141;
  wire popcount30_96cy_core_142;
  wire popcount30_96cy_core_145;
  wire popcount30_96cy_core_146;
  wire popcount30_96cy_core_147_not;
  wire popcount30_96cy_core_148;
  wire popcount30_96cy_core_152;
  wire popcount30_96cy_core_153;
  wire popcount30_96cy_core_154;
  wire popcount30_96cy_core_156;
  wire popcount30_96cy_core_157;
  wire popcount30_96cy_core_158;
  wire popcount30_96cy_core_159;
  wire popcount30_96cy_core_160;
  wire popcount30_96cy_core_163;
  wire popcount30_96cy_core_166;
  wire popcount30_96cy_core_168;
  wire popcount30_96cy_core_171;
  wire popcount30_96cy_core_172;
  wire popcount30_96cy_core_173_not;
  wire popcount30_96cy_core_174_not;
  wire popcount30_96cy_core_175;
  wire popcount30_96cy_core_176;
  wire popcount30_96cy_core_179;
  wire popcount30_96cy_core_180;
  wire popcount30_96cy_core_181_not;
  wire popcount30_96cy_core_182;
  wire popcount30_96cy_core_183;
  wire popcount30_96cy_core_184;
  wire popcount30_96cy_core_185;
  wire popcount30_96cy_core_186;
  wire popcount30_96cy_core_189;
  wire popcount30_96cy_core_190;
  wire popcount30_96cy_core_191;
  wire popcount30_96cy_core_193;
  wire popcount30_96cy_core_194;
  wire popcount30_96cy_core_195;
  wire popcount30_96cy_core_197;
  wire popcount30_96cy_core_199;
  wire popcount30_96cy_core_202;
  wire popcount30_96cy_core_204;
  wire popcount30_96cy_core_205;
  wire popcount30_96cy_core_206;
  wire popcount30_96cy_core_208;
  wire popcount30_96cy_core_209;
  wire popcount30_96cy_core_210;
  wire popcount30_96cy_core_211;
  wire popcount30_96cy_core_213;

  assign popcount30_96cy_core_032 = ~(input_a[24] ^ input_a[19]);
  assign popcount30_96cy_core_033 = ~(input_a[16] | input_a[2]);
  assign popcount30_96cy_core_034 = ~(input_a[28] & input_a[13]);
  assign popcount30_96cy_core_035 = input_a[5] & input_a[22];
  assign popcount30_96cy_core_036 = input_a[16] & input_a[18];
  assign popcount30_96cy_core_038 = ~input_a[24];
  assign popcount30_96cy_core_041 = ~(input_a[20] & input_a[27]);
  assign popcount30_96cy_core_043 = input_a[12] | input_a[23];
  assign popcount30_96cy_core_044 = input_a[26] ^ input_a[21];
  assign popcount30_96cy_core_045 = ~(input_a[27] ^ input_a[22]);
  assign popcount30_96cy_core_046 = ~(input_a[28] & input_a[1]);
  assign popcount30_96cy_core_048 = ~(input_a[10] & input_a[29]);
  assign popcount30_96cy_core_049 = ~(input_a[3] ^ input_a[10]);
  assign popcount30_96cy_core_050 = input_a[21] | input_a[20];
  assign popcount30_96cy_core_051 = ~(input_a[15] & input_a[24]);
  assign popcount30_96cy_core_053 = ~input_a[20];
  assign popcount30_96cy_core_054 = ~input_a[24];
  assign popcount30_96cy_core_058 = input_a[22] & input_a[26];
  assign popcount30_96cy_core_061 = input_a[8] ^ input_a[6];
  assign popcount30_96cy_core_065 = ~(input_a[11] & input_a[14]);
  assign popcount30_96cy_core_068 = input_a[11] ^ input_a[28];
  assign popcount30_96cy_core_069 = ~(input_a[28] & input_a[0]);
  assign popcount30_96cy_core_070 = ~input_a[17];
  assign popcount30_96cy_core_071 = ~(input_a[2] | input_a[10]);
  assign popcount30_96cy_core_072 = ~(input_a[20] | input_a[19]);
  assign popcount30_96cy_core_073 = ~input_a[5];
  assign popcount30_96cy_core_074 = ~(input_a[27] ^ input_a[0]);
  assign popcount30_96cy_core_075 = ~(input_a[24] & input_a[0]);
  assign popcount30_96cy_core_078 = ~(input_a[6] & input_a[13]);
  assign popcount30_96cy_core_079 = input_a[24] ^ input_a[14];
  assign popcount30_96cy_core_080 = ~(input_a[0] ^ input_a[7]);
  assign popcount30_96cy_core_090 = ~(input_a[5] ^ input_a[0]);
  assign popcount30_96cy_core_093 = input_a[26] & input_a[9];
  assign popcount30_96cy_core_094 = input_a[2] ^ input_a[26];
  assign popcount30_96cy_core_096 = ~(input_a[16] | input_a[22]);
  assign popcount30_96cy_core_097 = ~(input_a[6] | input_a[6]);
  assign popcount30_96cy_core_098 = ~(input_a[18] ^ input_a[20]);
  assign popcount30_96cy_core_102 = ~(input_a[20] & input_a[20]);
  assign popcount30_96cy_core_105 = ~(input_a[5] ^ input_a[16]);
  assign popcount30_96cy_core_106 = ~(input_a[27] | input_a[27]);
  assign popcount30_96cy_core_109 = input_a[17] & input_a[16];
  assign popcount30_96cy_core_110 = ~input_a[19];
  assign popcount30_96cy_core_111 = ~input_a[20];
  assign popcount30_96cy_core_112 = ~(input_a[19] ^ input_a[6]);
  assign popcount30_96cy_core_114 = ~input_a[16];
  assign popcount30_96cy_core_115 = ~(input_a[28] | input_a[8]);
  assign popcount30_96cy_core_116 = input_a[19] ^ input_a[22];
  assign popcount30_96cy_core_118 = input_a[20] | input_a[4];
  assign popcount30_96cy_core_119 = input_a[21] ^ input_a[7];
  assign popcount30_96cy_core_121 = input_a[2] ^ input_a[22];
  assign popcount30_96cy_core_122_not = ~input_a[20];
  assign popcount30_96cy_core_123 = ~(input_a[20] & input_a[20]);
  assign popcount30_96cy_core_124 = ~(input_a[7] | input_a[29]);
  assign popcount30_96cy_core_125 = ~(input_a[12] | input_a[17]);
  assign popcount30_96cy_core_126 = ~(input_a[18] | input_a[24]);
  assign popcount30_96cy_core_128 = ~input_a[23];
  assign popcount30_96cy_core_129 = input_a[0] ^ input_a[24];
  assign popcount30_96cy_core_130 = ~(input_a[28] & input_a[17]);
  assign popcount30_96cy_core_131 = input_a[19] ^ input_a[25];
  assign popcount30_96cy_core_132 = ~input_a[17];
  assign popcount30_96cy_core_133 = input_a[21] | input_a[28];
  assign popcount30_96cy_core_136 = ~input_a[9];
  assign popcount30_96cy_core_139 = ~(input_a[11] | input_a[29]);
  assign popcount30_96cy_core_140 = ~(input_a[14] & input_a[18]);
  assign popcount30_96cy_core_141 = input_a[0] ^ input_a[0];
  assign popcount30_96cy_core_142 = ~(input_a[17] ^ input_a[3]);
  assign popcount30_96cy_core_145 = ~(input_a[18] & input_a[8]);
  assign popcount30_96cy_core_146 = ~(input_a[24] ^ input_a[25]);
  assign popcount30_96cy_core_147_not = ~input_a[3];
  assign popcount30_96cy_core_148 = ~input_a[19];
  assign popcount30_96cy_core_152 = input_a[14] | input_a[17];
  assign popcount30_96cy_core_153 = input_a[9] & input_a[16];
  assign popcount30_96cy_core_154 = input_a[12] | input_a[29];
  assign popcount30_96cy_core_156 = ~(input_a[6] & input_a[23]);
  assign popcount30_96cy_core_157 = ~(input_a[1] ^ input_a[5]);
  assign popcount30_96cy_core_158 = input_a[4] | input_a[25];
  assign popcount30_96cy_core_159 = input_a[16] & input_a[5];
  assign popcount30_96cy_core_160 = ~(input_a[12] | input_a[24]);
  assign popcount30_96cy_core_163 = input_a[27] ^ input_a[17];
  assign popcount30_96cy_core_166 = ~(input_a[2] & input_a[17]);
  assign popcount30_96cy_core_168 = ~(input_a[18] & input_a[17]);
  assign popcount30_96cy_core_171 = ~(input_a[18] | input_a[10]);
  assign popcount30_96cy_core_172 = input_a[7] & input_a[28];
  assign popcount30_96cy_core_173_not = ~input_a[6];
  assign popcount30_96cy_core_174_not = ~input_a[22];
  assign popcount30_96cy_core_175 = ~(input_a[17] | input_a[1]);
  assign popcount30_96cy_core_176 = ~(input_a[3] & input_a[11]);
  assign popcount30_96cy_core_179 = ~(input_a[26] | input_a[9]);
  assign popcount30_96cy_core_180 = ~(input_a[21] | input_a[18]);
  assign popcount30_96cy_core_181_not = ~input_a[10];
  assign popcount30_96cy_core_182 = ~(input_a[18] | input_a[21]);
  assign popcount30_96cy_core_183 = input_a[3] & input_a[18];
  assign popcount30_96cy_core_184 = ~(input_a[19] ^ input_a[13]);
  assign popcount30_96cy_core_185 = ~(input_a[27] | input_a[3]);
  assign popcount30_96cy_core_186 = ~(input_a[26] ^ input_a[17]);
  assign popcount30_96cy_core_189 = ~(input_a[23] ^ input_a[4]);
  assign popcount30_96cy_core_190 = ~(input_a[29] ^ input_a[7]);
  assign popcount30_96cy_core_191 = ~(input_a[16] & input_a[0]);
  assign popcount30_96cy_core_193 = input_a[3] & input_a[28];
  assign popcount30_96cy_core_194 = input_a[15] & input_a[28];
  assign popcount30_96cy_core_195 = ~(input_a[15] | input_a[9]);
  assign popcount30_96cy_core_197 = ~(input_a[5] ^ input_a[17]);
  assign popcount30_96cy_core_199 = ~input_a[7];
  assign popcount30_96cy_core_202 = input_a[4] | input_a[3];
  assign popcount30_96cy_core_204 = ~(input_a[16] & input_a[26]);
  assign popcount30_96cy_core_205 = ~(input_a[0] & input_a[14]);
  assign popcount30_96cy_core_206 = ~(input_a[25] | input_a[18]);
  assign popcount30_96cy_core_208 = input_a[8] & input_a[23];
  assign popcount30_96cy_core_209 = ~(input_a[7] & input_a[1]);
  assign popcount30_96cy_core_210 = ~(input_a[29] ^ input_a[28]);
  assign popcount30_96cy_core_211 = ~(input_a[26] | input_a[7]);
  assign popcount30_96cy_core_213 = input_a[10] & input_a[7];

  assign popcount30_96cy_out[0] = input_a[23];
  assign popcount30_96cy_out[1] = 1'b0;
  assign popcount30_96cy_out[2] = 1'b0;
  assign popcount30_96cy_out[3] = 1'b0;
  assign popcount30_96cy_out[4] = 1'b1;
endmodule