// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.84587
// WCE=20.0
// EP=0.830224%
// Printed PDK parameters:
//  Area=45819608.0
//  Delay=77341296.0
//  Power=2410400.0

module popcount38_akwm(input [37:0] input_a, output [5:0] popcount38_akwm_out);
  wire popcount38_akwm_core_040;
  wire popcount38_akwm_core_041;
  wire popcount38_akwm_core_042;
  wire popcount38_akwm_core_043;
  wire popcount38_akwm_core_045;
  wire popcount38_akwm_core_047;
  wire popcount38_akwm_core_049;
  wire popcount38_akwm_core_051;
  wire popcount38_akwm_core_053_not;
  wire popcount38_akwm_core_055;
  wire popcount38_akwm_core_059;
  wire popcount38_akwm_core_061;
  wire popcount38_akwm_core_063;
  wire popcount38_akwm_core_064;
  wire popcount38_akwm_core_065;
  wire popcount38_akwm_core_068;
  wire popcount38_akwm_core_070;
  wire popcount38_akwm_core_071;
  wire popcount38_akwm_core_073;
  wire popcount38_akwm_core_074;
  wire popcount38_akwm_core_075;
  wire popcount38_akwm_core_076;
  wire popcount38_akwm_core_078_not;
  wire popcount38_akwm_core_079;
  wire popcount38_akwm_core_082;
  wire popcount38_akwm_core_083;
  wire popcount38_akwm_core_084;
  wire popcount38_akwm_core_085;
  wire popcount38_akwm_core_086;
  wire popcount38_akwm_core_087;
  wire popcount38_akwm_core_088;
  wire popcount38_akwm_core_091;
  wire popcount38_akwm_core_092;
  wire popcount38_akwm_core_093;
  wire popcount38_akwm_core_094;
  wire popcount38_akwm_core_095;
  wire popcount38_akwm_core_096;
  wire popcount38_akwm_core_098;
  wire popcount38_akwm_core_100;
  wire popcount38_akwm_core_101;
  wire popcount38_akwm_core_102;
  wire popcount38_akwm_core_104;
  wire popcount38_akwm_core_105;
  wire popcount38_akwm_core_108;
  wire popcount38_akwm_core_109;
  wire popcount38_akwm_core_110;
  wire popcount38_akwm_core_111;
  wire popcount38_akwm_core_112;
  wire popcount38_akwm_core_113;
  wire popcount38_akwm_core_115;
  wire popcount38_akwm_core_116;
  wire popcount38_akwm_core_117;
  wire popcount38_akwm_core_118;
  wire popcount38_akwm_core_119;
  wire popcount38_akwm_core_120;
  wire popcount38_akwm_core_121;
  wire popcount38_akwm_core_122;
  wire popcount38_akwm_core_123;
  wire popcount38_akwm_core_125;
  wire popcount38_akwm_core_127;
  wire popcount38_akwm_core_129;
  wire popcount38_akwm_core_131;
  wire popcount38_akwm_core_132;
  wire popcount38_akwm_core_134;
  wire popcount38_akwm_core_137;
  wire popcount38_akwm_core_138;
  wire popcount38_akwm_core_140_not;
  wire popcount38_akwm_core_142;
  wire popcount38_akwm_core_143;
  wire popcount38_akwm_core_144;
  wire popcount38_akwm_core_147;
  wire popcount38_akwm_core_148;
  wire popcount38_akwm_core_149;
  wire popcount38_akwm_core_150;
  wire popcount38_akwm_core_151;
  wire popcount38_akwm_core_153;
  wire popcount38_akwm_core_154;
  wire popcount38_akwm_core_155;
  wire popcount38_akwm_core_157;
  wire popcount38_akwm_core_158;
  wire popcount38_akwm_core_159;
  wire popcount38_akwm_core_160;
  wire popcount38_akwm_core_161;
  wire popcount38_akwm_core_162;
  wire popcount38_akwm_core_163;
  wire popcount38_akwm_core_164;
  wire popcount38_akwm_core_166;
  wire popcount38_akwm_core_167;
  wire popcount38_akwm_core_168;
  wire popcount38_akwm_core_169;
  wire popcount38_akwm_core_172;
  wire popcount38_akwm_core_174;
  wire popcount38_akwm_core_175;
  wire popcount38_akwm_core_176;
  wire popcount38_akwm_core_177;
  wire popcount38_akwm_core_178;
  wire popcount38_akwm_core_179;
  wire popcount38_akwm_core_180;
  wire popcount38_akwm_core_183;
  wire popcount38_akwm_core_185;
  wire popcount38_akwm_core_186;
  wire popcount38_akwm_core_187;
  wire popcount38_akwm_core_188;
  wire popcount38_akwm_core_189;
  wire popcount38_akwm_core_190;
  wire popcount38_akwm_core_191;
  wire popcount38_akwm_core_192;
  wire popcount38_akwm_core_193;
  wire popcount38_akwm_core_194;
  wire popcount38_akwm_core_196;
  wire popcount38_akwm_core_198;
  wire popcount38_akwm_core_200;
  wire popcount38_akwm_core_202;
  wire popcount38_akwm_core_204;
  wire popcount38_akwm_core_208;
  wire popcount38_akwm_core_211;
  wire popcount38_akwm_core_213;
  wire popcount38_akwm_core_214;
  wire popcount38_akwm_core_215;
  wire popcount38_akwm_core_218;
  wire popcount38_akwm_core_219;
  wire popcount38_akwm_core_220;
  wire popcount38_akwm_core_221;
  wire popcount38_akwm_core_224;
  wire popcount38_akwm_core_226;
  wire popcount38_akwm_core_227;
  wire popcount38_akwm_core_229;
  wire popcount38_akwm_core_232;
  wire popcount38_akwm_core_236;
  wire popcount38_akwm_core_237;
  wire popcount38_akwm_core_243;
  wire popcount38_akwm_core_244;
  wire popcount38_akwm_core_247;
  wire popcount38_akwm_core_248;
  wire popcount38_akwm_core_251;
  wire popcount38_akwm_core_253;
  wire popcount38_akwm_core_254;
  wire popcount38_akwm_core_255;
  wire popcount38_akwm_core_258_not;
  wire popcount38_akwm_core_261;
  wire popcount38_akwm_core_262;
  wire popcount38_akwm_core_263;
  wire popcount38_akwm_core_264;
  wire popcount38_akwm_core_265;
  wire popcount38_akwm_core_266;
  wire popcount38_akwm_core_268;
  wire popcount38_akwm_core_269;
  wire popcount38_akwm_core_270;
  wire popcount38_akwm_core_271;
  wire popcount38_akwm_core_272;
  wire popcount38_akwm_core_273;
  wire popcount38_akwm_core_274;
  wire popcount38_akwm_core_275;
  wire popcount38_akwm_core_276;
  wire popcount38_akwm_core_277;
  wire popcount38_akwm_core_278;
  wire popcount38_akwm_core_279;
  wire popcount38_akwm_core_280;
  wire popcount38_akwm_core_281;
  wire popcount38_akwm_core_282;
  wire popcount38_akwm_core_283;
  wire popcount38_akwm_core_284;
  wire popcount38_akwm_core_285;
  wire popcount38_akwm_core_286;
  wire popcount38_akwm_core_290;
  wire popcount38_akwm_core_291;
  wire popcount38_akwm_core_294;
  wire popcount38_akwm_core_295;

  assign popcount38_akwm_core_040 = ~(input_a[27] & input_a[32]);
  assign popcount38_akwm_core_041 = input_a[14] & input_a[15];
  assign popcount38_akwm_core_042 = ~(input_a[20] | input_a[14]);
  assign popcount38_akwm_core_043 = input_a[4] & input_a[24];
  assign popcount38_akwm_core_045 = ~(input_a[1] ^ input_a[16]);
  assign popcount38_akwm_core_047 = input_a[22] | input_a[16];
  assign popcount38_akwm_core_049 = ~(input_a[15] & input_a[36]);
  assign popcount38_akwm_core_051 = input_a[12] ^ input_a[22];
  assign popcount38_akwm_core_053_not = ~input_a[3];
  assign popcount38_akwm_core_055 = input_a[36] ^ input_a[26];
  assign popcount38_akwm_core_059 = ~(input_a[35] | input_a[35]);
  assign popcount38_akwm_core_061 = ~(input_a[31] | input_a[32]);
  assign popcount38_akwm_core_063 = input_a[35] & input_a[2];
  assign popcount38_akwm_core_064 = input_a[13] ^ input_a[6];
  assign popcount38_akwm_core_065 = input_a[24] ^ input_a[8];
  assign popcount38_akwm_core_068 = ~(input_a[18] ^ input_a[25]);
  assign popcount38_akwm_core_070 = ~input_a[16];
  assign popcount38_akwm_core_071 = input_a[19] ^ input_a[32];
  assign popcount38_akwm_core_073 = input_a[0] & input_a[10];
  assign popcount38_akwm_core_074 = ~(input_a[6] & input_a[30]);
  assign popcount38_akwm_core_075 = input_a[9] | input_a[25];
  assign popcount38_akwm_core_076 = ~(input_a[23] ^ input_a[0]);
  assign popcount38_akwm_core_078_not = ~input_a[20];
  assign popcount38_akwm_core_079 = input_a[19] | input_a[34];
  assign popcount38_akwm_core_082 = input_a[18] & input_a[37];
  assign popcount38_akwm_core_083 = input_a[9] & input_a[10];
  assign popcount38_akwm_core_084 = input_a[12] ^ input_a[34];
  assign popcount38_akwm_core_085 = input_a[5] & input_a[25];
  assign popcount38_akwm_core_086 = ~(input_a[29] | input_a[6]);
  assign popcount38_akwm_core_087 = input_a[11] & input_a[31];
  assign popcount38_akwm_core_088 = popcount38_akwm_core_085 | popcount38_akwm_core_087;
  assign popcount38_akwm_core_091 = input_a[13] & input_a[24];
  assign popcount38_akwm_core_092 = popcount38_akwm_core_083 ^ popcount38_akwm_core_088;
  assign popcount38_akwm_core_093 = popcount38_akwm_core_083 & popcount38_akwm_core_088;
  assign popcount38_akwm_core_094 = popcount38_akwm_core_092 ^ popcount38_akwm_core_091;
  assign popcount38_akwm_core_095 = popcount38_akwm_core_092 & popcount38_akwm_core_091;
  assign popcount38_akwm_core_096 = popcount38_akwm_core_093 | popcount38_akwm_core_095;
  assign popcount38_akwm_core_098 = ~(input_a[28] & input_a[29]);
  assign popcount38_akwm_core_100 = input_a[14] & input_a[34];
  assign popcount38_akwm_core_101 = input_a[17] ^ input_a[18];
  assign popcount38_akwm_core_102 = input_a[17] & input_a[18];
  assign popcount38_akwm_core_104 = input_a[4] & input_a[16];
  assign popcount38_akwm_core_105 = popcount38_akwm_core_102 | popcount38_akwm_core_104;
  assign popcount38_akwm_core_108 = input_a[6] & input_a[28];
  assign popcount38_akwm_core_109 = popcount38_akwm_core_100 ^ popcount38_akwm_core_105;
  assign popcount38_akwm_core_110 = popcount38_akwm_core_100 & popcount38_akwm_core_105;
  assign popcount38_akwm_core_111 = popcount38_akwm_core_109 ^ popcount38_akwm_core_108;
  assign popcount38_akwm_core_112 = popcount38_akwm_core_109 & popcount38_akwm_core_108;
  assign popcount38_akwm_core_113 = popcount38_akwm_core_110 | popcount38_akwm_core_112;
  assign popcount38_akwm_core_115 = ~(input_a[9] | input_a[32]);
  assign popcount38_akwm_core_116 = ~(input_a[33] | input_a[32]);
  assign popcount38_akwm_core_117 = input_a[36] & input_a[12];
  assign popcount38_akwm_core_118 = popcount38_akwm_core_094 ^ popcount38_akwm_core_111;
  assign popcount38_akwm_core_119 = popcount38_akwm_core_094 & popcount38_akwm_core_111;
  assign popcount38_akwm_core_120 = popcount38_akwm_core_118 ^ popcount38_akwm_core_117;
  assign popcount38_akwm_core_121 = popcount38_akwm_core_118 & popcount38_akwm_core_117;
  assign popcount38_akwm_core_122 = popcount38_akwm_core_119 | popcount38_akwm_core_121;
  assign popcount38_akwm_core_123 = popcount38_akwm_core_096 | popcount38_akwm_core_113;
  assign popcount38_akwm_core_125 = popcount38_akwm_core_123 ^ popcount38_akwm_core_122;
  assign popcount38_akwm_core_127 = popcount38_akwm_core_096 | popcount38_akwm_core_123;
  assign popcount38_akwm_core_129 = ~(input_a[16] ^ input_a[29]);
  assign popcount38_akwm_core_131 = ~(input_a[36] ^ input_a[5]);
  assign popcount38_akwm_core_132 = ~(input_a[14] ^ input_a[32]);
  assign popcount38_akwm_core_134 = input_a[29] & input_a[20];
  assign popcount38_akwm_core_137 = popcount38_akwm_core_120 ^ popcount38_akwm_core_134;
  assign popcount38_akwm_core_138 = popcount38_akwm_core_120 & popcount38_akwm_core_134;
  assign popcount38_akwm_core_140_not = ~popcount38_akwm_core_125;
  assign popcount38_akwm_core_142 = popcount38_akwm_core_140_not ^ popcount38_akwm_core_138;
  assign popcount38_akwm_core_143 = input_a[20] & popcount38_akwm_core_138;
  assign popcount38_akwm_core_144 = popcount38_akwm_core_125 | popcount38_akwm_core_143;
  assign popcount38_akwm_core_147 = popcount38_akwm_core_127 | popcount38_akwm_core_144;
  assign popcount38_akwm_core_148 = ~(input_a[22] | input_a[22]);
  assign popcount38_akwm_core_149 = ~(input_a[16] ^ input_a[32]);
  assign popcount38_akwm_core_150 = ~(input_a[13] ^ input_a[28]);
  assign popcount38_akwm_core_151 = ~(input_a[13] | input_a[14]);
  assign popcount38_akwm_core_153 = input_a[29] & input_a[37];
  assign popcount38_akwm_core_154 = ~input_a[1];
  assign popcount38_akwm_core_155 = ~input_a[35];
  assign popcount38_akwm_core_157 = ~(input_a[21] & input_a[22]);
  assign popcount38_akwm_core_158 = input_a[21] & input_a[22];
  assign popcount38_akwm_core_159 = ~(input_a[15] & input_a[8]);
  assign popcount38_akwm_core_160 = input_a[19] & popcount38_akwm_core_157;
  assign popcount38_akwm_core_161 = input_a[7] ^ popcount38_akwm_core_158;
  assign popcount38_akwm_core_162 = input_a[7] & popcount38_akwm_core_158;
  assign popcount38_akwm_core_163 = popcount38_akwm_core_161 | popcount38_akwm_core_160;
  assign popcount38_akwm_core_164 = input_a[14] | input_a[23];
  assign popcount38_akwm_core_166 = input_a[12] | input_a[14];
  assign popcount38_akwm_core_167 = input_a[2] & input_a[30];
  assign popcount38_akwm_core_168 = ~(input_a[9] ^ input_a[26]);
  assign popcount38_akwm_core_169 = input_a[33] & input_a[27];
  assign popcount38_akwm_core_172 = input_a[27] | input_a[1];
  assign popcount38_akwm_core_174 = ~(input_a[4] & input_a[20]);
  assign popcount38_akwm_core_175 = input_a[33] & input_a[8];
  assign popcount38_akwm_core_176 = popcount38_akwm_core_167 ^ popcount38_akwm_core_172;
  assign popcount38_akwm_core_177 = popcount38_akwm_core_167 & popcount38_akwm_core_172;
  assign popcount38_akwm_core_178 = popcount38_akwm_core_176 ^ popcount38_akwm_core_175;
  assign popcount38_akwm_core_179 = popcount38_akwm_core_176 & popcount38_akwm_core_175;
  assign popcount38_akwm_core_180 = popcount38_akwm_core_177 | popcount38_akwm_core_179;
  assign popcount38_akwm_core_183 = ~input_a[3];
  assign popcount38_akwm_core_185 = popcount38_akwm_core_163 ^ popcount38_akwm_core_178;
  assign popcount38_akwm_core_186 = popcount38_akwm_core_163 & popcount38_akwm_core_178;
  assign popcount38_akwm_core_187 = popcount38_akwm_core_185 ^ input_a[35];
  assign popcount38_akwm_core_188 = popcount38_akwm_core_185 & input_a[35];
  assign popcount38_akwm_core_189 = popcount38_akwm_core_186 | popcount38_akwm_core_188;
  assign popcount38_akwm_core_190 = popcount38_akwm_core_162 ^ popcount38_akwm_core_180;
  assign popcount38_akwm_core_191 = popcount38_akwm_core_162 & input_a[21];
  assign popcount38_akwm_core_192 = popcount38_akwm_core_190 ^ popcount38_akwm_core_189;
  assign popcount38_akwm_core_193 = popcount38_akwm_core_190 & popcount38_akwm_core_189;
  assign popcount38_akwm_core_194 = popcount38_akwm_core_191 | popcount38_akwm_core_193;
  assign popcount38_akwm_core_196 = ~(input_a[5] ^ input_a[12]);
  assign popcount38_akwm_core_198 = ~input_a[22];
  assign popcount38_akwm_core_200 = input_a[12] | input_a[18];
  assign popcount38_akwm_core_202 = ~(input_a[35] ^ input_a[3]);
  assign popcount38_akwm_core_204 = ~input_a[1];
  assign popcount38_akwm_core_208 = input_a[34] ^ input_a[22];
  assign popcount38_akwm_core_211 = input_a[16] | input_a[32];
  assign popcount38_akwm_core_213 = input_a[7] & input_a[7];
  assign popcount38_akwm_core_214 = ~input_a[6];
  assign popcount38_akwm_core_215 = ~(input_a[36] & input_a[4]);
  assign popcount38_akwm_core_218 = ~input_a[18];
  assign popcount38_akwm_core_219 = input_a[0] | input_a[22];
  assign popcount38_akwm_core_220 = input_a[18] | input_a[23];
  assign popcount38_akwm_core_221 = ~(input_a[0] ^ input_a[15]);
  assign popcount38_akwm_core_224 = ~(input_a[1] | input_a[6]);
  assign popcount38_akwm_core_226 = input_a[6] & input_a[20];
  assign popcount38_akwm_core_227 = input_a[5] ^ input_a[7];
  assign popcount38_akwm_core_229 = ~(input_a[36] | input_a[1]);
  assign popcount38_akwm_core_232 = ~(input_a[28] ^ input_a[19]);
  assign popcount38_akwm_core_236 = ~(input_a[1] & input_a[5]);
  assign popcount38_akwm_core_237 = input_a[6] & input_a[7];
  assign popcount38_akwm_core_243 = ~(input_a[26] & input_a[10]);
  assign popcount38_akwm_core_244 = ~(input_a[17] | input_a[0]);
  assign popcount38_akwm_core_247 = input_a[11] | input_a[1];
  assign popcount38_akwm_core_248 = ~popcount38_akwm_core_183;
  assign popcount38_akwm_core_251 = ~(input_a[14] & input_a[13]);
  assign popcount38_akwm_core_253 = input_a[1] ^ input_a[27];
  assign popcount38_akwm_core_254 = ~(input_a[36] & input_a[34]);
  assign popcount38_akwm_core_255 = ~popcount38_akwm_core_192;
  assign popcount38_akwm_core_258_not = ~input_a[1];
  assign popcount38_akwm_core_261 = input_a[25] | input_a[9];
  assign popcount38_akwm_core_262 = popcount38_akwm_core_194 | popcount38_akwm_core_192;
  assign popcount38_akwm_core_263 = input_a[36] & input_a[20];
  assign popcount38_akwm_core_264 = ~(input_a[27] ^ input_a[30]);
  assign popcount38_akwm_core_265 = input_a[8] ^ input_a[4];
  assign popcount38_akwm_core_266 = input_a[0] ^ input_a[2];
  assign popcount38_akwm_core_268 = ~(input_a[19] ^ input_a[17]);
  assign popcount38_akwm_core_269 = ~input_a[36];
  assign popcount38_akwm_core_270 = input_a[23] ^ popcount38_akwm_core_248;
  assign popcount38_akwm_core_271 = input_a[23] & popcount38_akwm_core_248;
  assign popcount38_akwm_core_272 = popcount38_akwm_core_137 ^ popcount38_akwm_core_187;
  assign popcount38_akwm_core_273 = popcount38_akwm_core_137 & popcount38_akwm_core_187;
  assign popcount38_akwm_core_274 = popcount38_akwm_core_272 ^ popcount38_akwm_core_271;
  assign popcount38_akwm_core_275 = popcount38_akwm_core_272 & popcount38_akwm_core_271;
  assign popcount38_akwm_core_276 = popcount38_akwm_core_273 | popcount38_akwm_core_275;
  assign popcount38_akwm_core_277 = popcount38_akwm_core_142 ^ popcount38_akwm_core_255;
  assign popcount38_akwm_core_278 = popcount38_akwm_core_142 & popcount38_akwm_core_255;
  assign popcount38_akwm_core_279 = popcount38_akwm_core_277 ^ popcount38_akwm_core_276;
  assign popcount38_akwm_core_280 = popcount38_akwm_core_277 & popcount38_akwm_core_276;
  assign popcount38_akwm_core_281 = popcount38_akwm_core_278 | popcount38_akwm_core_280;
  assign popcount38_akwm_core_282 = popcount38_akwm_core_147 ^ popcount38_akwm_core_262;
  assign popcount38_akwm_core_283 = popcount38_akwm_core_147 & popcount38_akwm_core_262;
  assign popcount38_akwm_core_284 = popcount38_akwm_core_282 ^ popcount38_akwm_core_281;
  assign popcount38_akwm_core_285 = popcount38_akwm_core_282 & popcount38_akwm_core_281;
  assign popcount38_akwm_core_286 = popcount38_akwm_core_283 | popcount38_akwm_core_285;
  assign popcount38_akwm_core_290 = input_a[21] & input_a[15];
  assign popcount38_akwm_core_291 = ~(input_a[22] & input_a[33]);
  assign popcount38_akwm_core_294 = ~(input_a[35] & input_a[27]);
  assign popcount38_akwm_core_295 = input_a[9] | input_a[10];

  assign popcount38_akwm_out[0] = popcount38_akwm_core_270;
  assign popcount38_akwm_out[1] = popcount38_akwm_core_274;
  assign popcount38_akwm_out[2] = popcount38_akwm_core_279;
  assign popcount38_akwm_out[3] = popcount38_akwm_core_284;
  assign popcount38_akwm_out[4] = popcount38_akwm_core_286;
  assign popcount38_akwm_out[5] = 1'b0;
endmodule