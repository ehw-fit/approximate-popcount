// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.00206
// WCE=19.0
// EP=0.897168%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_mpnk(input [32:0] input_a, output [5:0] popcount33_mpnk_out);
  wire popcount33_mpnk_core_035;
  wire popcount33_mpnk_core_037;
  wire popcount33_mpnk_core_039;
  wire popcount33_mpnk_core_040;
  wire popcount33_mpnk_core_041;
  wire popcount33_mpnk_core_043;
  wire popcount33_mpnk_core_044;
  wire popcount33_mpnk_core_045;
  wire popcount33_mpnk_core_046;
  wire popcount33_mpnk_core_048;
  wire popcount33_mpnk_core_050;
  wire popcount33_mpnk_core_051;
  wire popcount33_mpnk_core_054;
  wire popcount33_mpnk_core_055;
  wire popcount33_mpnk_core_056;
  wire popcount33_mpnk_core_057;
  wire popcount33_mpnk_core_058;
  wire popcount33_mpnk_core_059;
  wire popcount33_mpnk_core_060;
  wire popcount33_mpnk_core_061;
  wire popcount33_mpnk_core_064;
  wire popcount33_mpnk_core_066;
  wire popcount33_mpnk_core_070;
  wire popcount33_mpnk_core_071;
  wire popcount33_mpnk_core_074;
  wire popcount33_mpnk_core_075;
  wire popcount33_mpnk_core_077;
  wire popcount33_mpnk_core_078;
  wire popcount33_mpnk_core_079;
  wire popcount33_mpnk_core_081;
  wire popcount33_mpnk_core_082;
  wire popcount33_mpnk_core_083;
  wire popcount33_mpnk_core_085;
  wire popcount33_mpnk_core_086;
  wire popcount33_mpnk_core_087;
  wire popcount33_mpnk_core_088;
  wire popcount33_mpnk_core_090;
  wire popcount33_mpnk_core_091;
  wire popcount33_mpnk_core_093;
  wire popcount33_mpnk_core_094;
  wire popcount33_mpnk_core_096;
  wire popcount33_mpnk_core_097;
  wire popcount33_mpnk_core_099;
  wire popcount33_mpnk_core_100;
  wire popcount33_mpnk_core_101;
  wire popcount33_mpnk_core_102;
  wire popcount33_mpnk_core_104;
  wire popcount33_mpnk_core_105;
  wire popcount33_mpnk_core_107;
  wire popcount33_mpnk_core_109;
  wire popcount33_mpnk_core_110;
  wire popcount33_mpnk_core_111;
  wire popcount33_mpnk_core_116;
  wire popcount33_mpnk_core_117;
  wire popcount33_mpnk_core_118;
  wire popcount33_mpnk_core_119;
  wire popcount33_mpnk_core_120;
  wire popcount33_mpnk_core_121;
  wire popcount33_mpnk_core_122;
  wire popcount33_mpnk_core_123_not;
  wire popcount33_mpnk_core_126;
  wire popcount33_mpnk_core_127;
  wire popcount33_mpnk_core_130;
  wire popcount33_mpnk_core_133;
  wire popcount33_mpnk_core_134;
  wire popcount33_mpnk_core_135_not;
  wire popcount33_mpnk_core_136;
  wire popcount33_mpnk_core_138;
  wire popcount33_mpnk_core_139;
  wire popcount33_mpnk_core_141;
  wire popcount33_mpnk_core_143;
  wire popcount33_mpnk_core_144;
  wire popcount33_mpnk_core_146;
  wire popcount33_mpnk_core_150;
  wire popcount33_mpnk_core_152;
  wire popcount33_mpnk_core_153;
  wire popcount33_mpnk_core_154;
  wire popcount33_mpnk_core_155;
  wire popcount33_mpnk_core_158;
  wire popcount33_mpnk_core_159;
  wire popcount33_mpnk_core_160;
  wire popcount33_mpnk_core_161;
  wire popcount33_mpnk_core_162;
  wire popcount33_mpnk_core_163;
  wire popcount33_mpnk_core_165;
  wire popcount33_mpnk_core_167;
  wire popcount33_mpnk_core_168;
  wire popcount33_mpnk_core_169;
  wire popcount33_mpnk_core_170;
  wire popcount33_mpnk_core_172;
  wire popcount33_mpnk_core_173;
  wire popcount33_mpnk_core_174;
  wire popcount33_mpnk_core_175;
  wire popcount33_mpnk_core_177;
  wire popcount33_mpnk_core_179;
  wire popcount33_mpnk_core_181;
  wire popcount33_mpnk_core_182;
  wire popcount33_mpnk_core_183;
  wire popcount33_mpnk_core_184;
  wire popcount33_mpnk_core_186;
  wire popcount33_mpnk_core_189;
  wire popcount33_mpnk_core_191;
  wire popcount33_mpnk_core_193;
  wire popcount33_mpnk_core_194;
  wire popcount33_mpnk_core_196;
  wire popcount33_mpnk_core_197;
  wire popcount33_mpnk_core_199;
  wire popcount33_mpnk_core_201;
  wire popcount33_mpnk_core_203;
  wire popcount33_mpnk_core_204;
  wire popcount33_mpnk_core_205;
  wire popcount33_mpnk_core_207;
  wire popcount33_mpnk_core_208;
  wire popcount33_mpnk_core_209;
  wire popcount33_mpnk_core_210;
  wire popcount33_mpnk_core_211;
  wire popcount33_mpnk_core_213;
  wire popcount33_mpnk_core_214;
  wire popcount33_mpnk_core_215;
  wire popcount33_mpnk_core_216;
  wire popcount33_mpnk_core_218;
  wire popcount33_mpnk_core_219;
  wire popcount33_mpnk_core_220;
  wire popcount33_mpnk_core_226;
  wire popcount33_mpnk_core_227;
  wire popcount33_mpnk_core_228;
  wire popcount33_mpnk_core_229;
  wire popcount33_mpnk_core_231_not;
  wire popcount33_mpnk_core_233;
  wire popcount33_mpnk_core_234;

  assign popcount33_mpnk_core_035 = ~(input_a[30] & input_a[8]);
  assign popcount33_mpnk_core_037 = ~(input_a[32] | input_a[19]);
  assign popcount33_mpnk_core_039 = ~(input_a[18] ^ input_a[10]);
  assign popcount33_mpnk_core_040 = ~(input_a[8] ^ input_a[9]);
  assign popcount33_mpnk_core_041 = ~(input_a[30] | input_a[11]);
  assign popcount33_mpnk_core_043 = ~input_a[26];
  assign popcount33_mpnk_core_044 = ~(input_a[30] & input_a[22]);
  assign popcount33_mpnk_core_045 = ~(input_a[9] ^ input_a[26]);
  assign popcount33_mpnk_core_046 = ~(input_a[7] & input_a[7]);
  assign popcount33_mpnk_core_048 = input_a[22] | input_a[16];
  assign popcount33_mpnk_core_050 = input_a[17] | input_a[16];
  assign popcount33_mpnk_core_051 = input_a[12] | input_a[10];
  assign popcount33_mpnk_core_054 = ~(input_a[24] & input_a[0]);
  assign popcount33_mpnk_core_055 = input_a[23] | input_a[28];
  assign popcount33_mpnk_core_056 = input_a[17] ^ input_a[20];
  assign popcount33_mpnk_core_057 = ~(input_a[22] & input_a[5]);
  assign popcount33_mpnk_core_058 = input_a[20] | input_a[19];
  assign popcount33_mpnk_core_059 = ~input_a[23];
  assign popcount33_mpnk_core_060 = ~input_a[13];
  assign popcount33_mpnk_core_061 = input_a[22] ^ input_a[28];
  assign popcount33_mpnk_core_064 = ~(input_a[1] ^ input_a[0]);
  assign popcount33_mpnk_core_066 = input_a[30] & input_a[7];
  assign popcount33_mpnk_core_070 = input_a[1] & input_a[6];
  assign popcount33_mpnk_core_071 = ~(input_a[0] ^ input_a[25]);
  assign popcount33_mpnk_core_074 = ~input_a[11];
  assign popcount33_mpnk_core_075 = ~input_a[8];
  assign popcount33_mpnk_core_077 = input_a[25] & input_a[25];
  assign popcount33_mpnk_core_078 = input_a[11] | input_a[28];
  assign popcount33_mpnk_core_079 = ~(input_a[1] & input_a[22]);
  assign popcount33_mpnk_core_081 = ~input_a[19];
  assign popcount33_mpnk_core_082 = ~input_a[11];
  assign popcount33_mpnk_core_083 = ~(input_a[25] ^ input_a[31]);
  assign popcount33_mpnk_core_085 = ~(input_a[32] ^ input_a[21]);
  assign popcount33_mpnk_core_086 = input_a[13] & input_a[13];
  assign popcount33_mpnk_core_087 = ~input_a[6];
  assign popcount33_mpnk_core_088 = ~(input_a[27] ^ input_a[23]);
  assign popcount33_mpnk_core_090 = ~(input_a[18] | input_a[16]);
  assign popcount33_mpnk_core_091 = input_a[4] | input_a[15];
  assign popcount33_mpnk_core_093 = ~input_a[29];
  assign popcount33_mpnk_core_094 = ~(input_a[2] ^ input_a[7]);
  assign popcount33_mpnk_core_096 = input_a[0] | input_a[23];
  assign popcount33_mpnk_core_097 = input_a[9] | input_a[28];
  assign popcount33_mpnk_core_099 = ~(input_a[13] ^ input_a[16]);
  assign popcount33_mpnk_core_100 = ~(input_a[29] | input_a[22]);
  assign popcount33_mpnk_core_101 = input_a[27] ^ input_a[25];
  assign popcount33_mpnk_core_102 = input_a[30] & input_a[8];
  assign popcount33_mpnk_core_104 = input_a[3] & input_a[18];
  assign popcount33_mpnk_core_105 = input_a[20] | input_a[10];
  assign popcount33_mpnk_core_107 = ~(input_a[32] & input_a[30]);
  assign popcount33_mpnk_core_109 = ~input_a[28];
  assign popcount33_mpnk_core_110 = ~input_a[8];
  assign popcount33_mpnk_core_111 = ~(input_a[1] & input_a[22]);
  assign popcount33_mpnk_core_116 = input_a[24] ^ input_a[12];
  assign popcount33_mpnk_core_117 = ~(input_a[4] & input_a[19]);
  assign popcount33_mpnk_core_118 = input_a[27] & input_a[1];
  assign popcount33_mpnk_core_119 = input_a[4] | input_a[19];
  assign popcount33_mpnk_core_120 = ~(input_a[24] | input_a[14]);
  assign popcount33_mpnk_core_121 = ~input_a[29];
  assign popcount33_mpnk_core_122 = input_a[7] & input_a[1];
  assign popcount33_mpnk_core_123_not = ~input_a[25];
  assign popcount33_mpnk_core_126 = ~(input_a[23] | input_a[0]);
  assign popcount33_mpnk_core_127 = ~(input_a[23] ^ input_a[22]);
  assign popcount33_mpnk_core_130 = ~(input_a[27] ^ input_a[6]);
  assign popcount33_mpnk_core_133 = ~(input_a[21] | input_a[26]);
  assign popcount33_mpnk_core_134 = input_a[32] | input_a[13];
  assign popcount33_mpnk_core_135_not = ~input_a[14];
  assign popcount33_mpnk_core_136 = ~(input_a[0] ^ input_a[24]);
  assign popcount33_mpnk_core_138 = ~(input_a[18] | input_a[28]);
  assign popcount33_mpnk_core_139 = ~input_a[7];
  assign popcount33_mpnk_core_141 = ~(input_a[2] & input_a[31]);
  assign popcount33_mpnk_core_143 = input_a[16] ^ input_a[25];
  assign popcount33_mpnk_core_144 = ~(input_a[14] | input_a[25]);
  assign popcount33_mpnk_core_146 = ~(input_a[22] ^ input_a[4]);
  assign popcount33_mpnk_core_150 = ~(input_a[26] ^ input_a[5]);
  assign popcount33_mpnk_core_152 = input_a[30] | input_a[6];
  assign popcount33_mpnk_core_153 = input_a[1] | input_a[17];
  assign popcount33_mpnk_core_154 = ~(input_a[27] ^ input_a[28]);
  assign popcount33_mpnk_core_155 = ~(input_a[17] ^ input_a[3]);
  assign popcount33_mpnk_core_158 = input_a[22] | input_a[9];
  assign popcount33_mpnk_core_159 = input_a[27] & input_a[24];
  assign popcount33_mpnk_core_160 = input_a[2] | input_a[16];
  assign popcount33_mpnk_core_161 = input_a[25] & input_a[20];
  assign popcount33_mpnk_core_162 = input_a[31] | input_a[8];
  assign popcount33_mpnk_core_163 = input_a[26] & input_a[12];
  assign popcount33_mpnk_core_165 = ~(input_a[30] ^ input_a[20]);
  assign popcount33_mpnk_core_167 = input_a[22] ^ input_a[28];
  assign popcount33_mpnk_core_168 = input_a[11] ^ input_a[13];
  assign popcount33_mpnk_core_169 = ~(input_a[13] & input_a[10]);
  assign popcount33_mpnk_core_170 = input_a[19] | input_a[23];
  assign popcount33_mpnk_core_172 = ~(input_a[25] & input_a[3]);
  assign popcount33_mpnk_core_173 = ~(input_a[4] | input_a[31]);
  assign popcount33_mpnk_core_174 = ~input_a[8];
  assign popcount33_mpnk_core_175 = input_a[29] & input_a[24];
  assign popcount33_mpnk_core_177 = input_a[25] | input_a[20];
  assign popcount33_mpnk_core_179 = ~(input_a[15] | input_a[32]);
  assign popcount33_mpnk_core_181 = input_a[7] & input_a[3];
  assign popcount33_mpnk_core_182 = ~(input_a[6] & input_a[13]);
  assign popcount33_mpnk_core_183 = input_a[20] ^ input_a[13];
  assign popcount33_mpnk_core_184 = ~(input_a[0] & input_a[10]);
  assign popcount33_mpnk_core_186 = input_a[21] | input_a[19];
  assign popcount33_mpnk_core_189 = ~(input_a[30] | input_a[8]);
  assign popcount33_mpnk_core_191 = ~input_a[31];
  assign popcount33_mpnk_core_193 = ~(input_a[32] & input_a[26]);
  assign popcount33_mpnk_core_194 = ~(input_a[6] ^ input_a[4]);
  assign popcount33_mpnk_core_196 = ~input_a[5];
  assign popcount33_mpnk_core_197 = ~(input_a[5] & input_a[2]);
  assign popcount33_mpnk_core_199 = ~input_a[24];
  assign popcount33_mpnk_core_201 = ~(input_a[21] ^ input_a[11]);
  assign popcount33_mpnk_core_203 = input_a[21] ^ input_a[29];
  assign popcount33_mpnk_core_204 = input_a[23] | input_a[31];
  assign popcount33_mpnk_core_205 = input_a[21] ^ input_a[30];
  assign popcount33_mpnk_core_207 = ~(input_a[8] ^ input_a[5]);
  assign popcount33_mpnk_core_208 = ~input_a[0];
  assign popcount33_mpnk_core_209 = input_a[17] ^ input_a[26];
  assign popcount33_mpnk_core_210 = ~(input_a[17] | input_a[30]);
  assign popcount33_mpnk_core_211 = input_a[27] & input_a[13];
  assign popcount33_mpnk_core_213 = input_a[11] ^ input_a[32];
  assign popcount33_mpnk_core_214 = ~(input_a[3] & input_a[27]);
  assign popcount33_mpnk_core_215 = input_a[5] ^ input_a[16];
  assign popcount33_mpnk_core_216 = ~(input_a[30] ^ input_a[18]);
  assign popcount33_mpnk_core_218 = ~(input_a[30] & input_a[21]);
  assign popcount33_mpnk_core_219 = input_a[9] ^ input_a[29];
  assign popcount33_mpnk_core_220 = input_a[32] | input_a[22];
  assign popcount33_mpnk_core_226 = input_a[6] & input_a[26];
  assign popcount33_mpnk_core_227 = ~(input_a[12] & input_a[23]);
  assign popcount33_mpnk_core_228 = ~(input_a[17] ^ input_a[20]);
  assign popcount33_mpnk_core_229 = input_a[14] | input_a[17];
  assign popcount33_mpnk_core_231_not = ~input_a[29];
  assign popcount33_mpnk_core_233 = input_a[30] ^ input_a[20];
  assign popcount33_mpnk_core_234 = input_a[20] | input_a[25];

  assign popcount33_mpnk_out[0] = input_a[11];
  assign popcount33_mpnk_out[1] = 1'b0;
  assign popcount33_mpnk_out[2] = input_a[1];
  assign popcount33_mpnk_out[3] = 1'b0;
  assign popcount33_mpnk_out[4] = 1'b1;
  assign popcount33_mpnk_out[5] = 1'b0;
endmodule