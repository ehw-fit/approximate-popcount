// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.80172
// WCE=18.0
// EP=0.890175%
// Printed PDK parameters:
//  Area=7320940.0
//  Delay=19521304.0
//  Power=240110.0

module popcount36_pgij(input [35:0] input_a, output [5:0] popcount36_pgij_out);
  wire popcount36_pgij_core_038;
  wire popcount36_pgij_core_039;
  wire popcount36_pgij_core_040;
  wire popcount36_pgij_core_042;
  wire popcount36_pgij_core_043;
  wire popcount36_pgij_core_044;
  wire popcount36_pgij_core_047;
  wire popcount36_pgij_core_048;
  wire popcount36_pgij_core_053;
  wire popcount36_pgij_core_054;
  wire popcount36_pgij_core_055;
  wire popcount36_pgij_core_056;
  wire popcount36_pgij_core_058;
  wire popcount36_pgij_core_059;
  wire popcount36_pgij_core_061;
  wire popcount36_pgij_core_063;
  wire popcount36_pgij_core_065;
  wire popcount36_pgij_core_066;
  wire popcount36_pgij_core_067;
  wire popcount36_pgij_core_071;
  wire popcount36_pgij_core_072;
  wire popcount36_pgij_core_073;
  wire popcount36_pgij_core_078;
  wire popcount36_pgij_core_079;
  wire popcount36_pgij_core_080;
  wire popcount36_pgij_core_082;
  wire popcount36_pgij_core_083;
  wire popcount36_pgij_core_084;
  wire popcount36_pgij_core_085;
  wire popcount36_pgij_core_087;
  wire popcount36_pgij_core_088;
  wire popcount36_pgij_core_089;
  wire popcount36_pgij_core_090;
  wire popcount36_pgij_core_091;
  wire popcount36_pgij_core_092;
  wire popcount36_pgij_core_095;
  wire popcount36_pgij_core_097;
  wire popcount36_pgij_core_098;
  wire popcount36_pgij_core_101;
  wire popcount36_pgij_core_102;
  wire popcount36_pgij_core_103;
  wire popcount36_pgij_core_104;
  wire popcount36_pgij_core_106;
  wire popcount36_pgij_core_107;
  wire popcount36_pgij_core_109;
  wire popcount36_pgij_core_110;
  wire popcount36_pgij_core_112;
  wire popcount36_pgij_core_113;
  wire popcount36_pgij_core_114;
  wire popcount36_pgij_core_115;
  wire popcount36_pgij_core_116;
  wire popcount36_pgij_core_118;
  wire popcount36_pgij_core_120;
  wire popcount36_pgij_core_121;
  wire popcount36_pgij_core_122;
  wire popcount36_pgij_core_123;
  wire popcount36_pgij_core_124;
  wire popcount36_pgij_core_125;
  wire popcount36_pgij_core_127;
  wire popcount36_pgij_core_128;
  wire popcount36_pgij_core_129;
  wire popcount36_pgij_core_130;
  wire popcount36_pgij_core_131;
  wire popcount36_pgij_core_133;
  wire popcount36_pgij_core_134;
  wire popcount36_pgij_core_135;
  wire popcount36_pgij_core_136;
  wire popcount36_pgij_core_137;
  wire popcount36_pgij_core_141;
  wire popcount36_pgij_core_143;
  wire popcount36_pgij_core_144;
  wire popcount36_pgij_core_146;
  wire popcount36_pgij_core_147;
  wire popcount36_pgij_core_148;
  wire popcount36_pgij_core_149;
  wire popcount36_pgij_core_150;
  wire popcount36_pgij_core_153;
  wire popcount36_pgij_core_154;
  wire popcount36_pgij_core_155;
  wire popcount36_pgij_core_156;
  wire popcount36_pgij_core_158;
  wire popcount36_pgij_core_159;
  wire popcount36_pgij_core_160;
  wire popcount36_pgij_core_165;
  wire popcount36_pgij_core_166;
  wire popcount36_pgij_core_167;
  wire popcount36_pgij_core_168;
  wire popcount36_pgij_core_169;
  wire popcount36_pgij_core_170;
  wire popcount36_pgij_core_171;
  wire popcount36_pgij_core_172;
  wire popcount36_pgij_core_173;
  wire popcount36_pgij_core_174;
  wire popcount36_pgij_core_175;
  wire popcount36_pgij_core_178;
  wire popcount36_pgij_core_179;
  wire popcount36_pgij_core_180_not;
  wire popcount36_pgij_core_181;
  wire popcount36_pgij_core_185;
  wire popcount36_pgij_core_186;
  wire popcount36_pgij_core_187;
  wire popcount36_pgij_core_188;
  wire popcount36_pgij_core_189;
  wire popcount36_pgij_core_193_not;
  wire popcount36_pgij_core_194;
  wire popcount36_pgij_core_196;
  wire popcount36_pgij_core_197;
  wire popcount36_pgij_core_198;
  wire popcount36_pgij_core_199;
  wire popcount36_pgij_core_201;
  wire popcount36_pgij_core_202;
  wire popcount36_pgij_core_203;
  wire popcount36_pgij_core_204;
  wire popcount36_pgij_core_205;
  wire popcount36_pgij_core_207;
  wire popcount36_pgij_core_208;
  wire popcount36_pgij_core_209;
  wire popcount36_pgij_core_213;
  wire popcount36_pgij_core_215;
  wire popcount36_pgij_core_216;
  wire popcount36_pgij_core_217;
  wire popcount36_pgij_core_218_not;
  wire popcount36_pgij_core_219;
  wire popcount36_pgij_core_223;
  wire popcount36_pgij_core_225;
  wire popcount36_pgij_core_227;
  wire popcount36_pgij_core_231;
  wire popcount36_pgij_core_232;
  wire popcount36_pgij_core_233;
  wire popcount36_pgij_core_234;
  wire popcount36_pgij_core_235;
  wire popcount36_pgij_core_237;
  wire popcount36_pgij_core_238;
  wire popcount36_pgij_core_239;
  wire popcount36_pgij_core_241;
  wire popcount36_pgij_core_242;
  wire popcount36_pgij_core_243;
  wire popcount36_pgij_core_244;
  wire popcount36_pgij_core_247;
  wire popcount36_pgij_core_249;
  wire popcount36_pgij_core_250;
  wire popcount36_pgij_core_251;
  wire popcount36_pgij_core_252;
  wire popcount36_pgij_core_255;
  wire popcount36_pgij_core_256;
  wire popcount36_pgij_core_257;
  wire popcount36_pgij_core_258;
  wire popcount36_pgij_core_259;
  wire popcount36_pgij_core_260;
  wire popcount36_pgij_core_261;
  wire popcount36_pgij_core_262;
  wire popcount36_pgij_core_264;
  wire popcount36_pgij_core_265;
  wire popcount36_pgij_core_266;
  wire popcount36_pgij_core_267;
  wire popcount36_pgij_core_268;
  wire popcount36_pgij_core_269;
  wire popcount36_pgij_core_270;
  wire popcount36_pgij_core_272;
  wire popcount36_pgij_core_273;
  wire popcount36_pgij_core_274;
  wire popcount36_pgij_core_275;

  assign popcount36_pgij_core_038 = ~(input_a[21] & input_a[30]);
  assign popcount36_pgij_core_039 = input_a[26] | input_a[17];
  assign popcount36_pgij_core_040 = input_a[9] ^ input_a[0];
  assign popcount36_pgij_core_042 = ~(input_a[24] ^ input_a[8]);
  assign popcount36_pgij_core_043 = input_a[0] | input_a[32];
  assign popcount36_pgij_core_044 = ~(input_a[31] ^ input_a[13]);
  assign popcount36_pgij_core_047 = ~input_a[12];
  assign popcount36_pgij_core_048 = input_a[13] ^ input_a[25];
  assign popcount36_pgij_core_053 = ~(input_a[17] | input_a[18]);
  assign popcount36_pgij_core_054 = input_a[26] & input_a[1];
  assign popcount36_pgij_core_055 = input_a[14] ^ input_a[20];
  assign popcount36_pgij_core_056 = ~input_a[0];
  assign popcount36_pgij_core_058 = ~(input_a[1] & input_a[18]);
  assign popcount36_pgij_core_059 = input_a[33] & input_a[15];
  assign popcount36_pgij_core_061 = input_a[2] & input_a[25];
  assign popcount36_pgij_core_063 = input_a[6] ^ input_a[5];
  assign popcount36_pgij_core_065 = input_a[0] & input_a[10];
  assign popcount36_pgij_core_066 = ~(input_a[0] | input_a[3]);
  assign popcount36_pgij_core_067 = ~(input_a[21] | input_a[7]);
  assign popcount36_pgij_core_071 = ~(input_a[35] & input_a[10]);
  assign popcount36_pgij_core_072 = ~(input_a[21] ^ input_a[28]);
  assign popcount36_pgij_core_073 = ~(input_a[3] & input_a[30]);
  assign popcount36_pgij_core_078 = input_a[18] | input_a[26];
  assign popcount36_pgij_core_079 = input_a[28] ^ input_a[19];
  assign popcount36_pgij_core_080 = ~(input_a[34] & input_a[1]);
  assign popcount36_pgij_core_082 = input_a[5] | input_a[19];
  assign popcount36_pgij_core_083 = ~(input_a[3] | input_a[20]);
  assign popcount36_pgij_core_084 = ~(input_a[21] ^ input_a[24]);
  assign popcount36_pgij_core_085 = ~(input_a[12] & input_a[17]);
  assign popcount36_pgij_core_087 = ~(input_a[18] ^ input_a[33]);
  assign popcount36_pgij_core_088 = input_a[30] ^ input_a[19];
  assign popcount36_pgij_core_089 = ~(input_a[31] & input_a[22]);
  assign popcount36_pgij_core_090 = input_a[34] & input_a[29];
  assign popcount36_pgij_core_091 = input_a[25] | input_a[19];
  assign popcount36_pgij_core_092 = ~input_a[6];
  assign popcount36_pgij_core_095 = ~(input_a[8] | input_a[23]);
  assign popcount36_pgij_core_097 = input_a[11] ^ input_a[9];
  assign popcount36_pgij_core_098 = ~(input_a[16] & input_a[10]);
  assign popcount36_pgij_core_101 = ~(input_a[9] ^ input_a[32]);
  assign popcount36_pgij_core_102 = input_a[13] | input_a[12];
  assign popcount36_pgij_core_103 = ~(input_a[23] | input_a[34]);
  assign popcount36_pgij_core_104 = ~(input_a[26] | input_a[4]);
  assign popcount36_pgij_core_106 = ~(input_a[22] ^ input_a[7]);
  assign popcount36_pgij_core_107 = input_a[17] ^ input_a[0];
  assign popcount36_pgij_core_109 = ~(input_a[33] & input_a[17]);
  assign popcount36_pgij_core_110 = ~(input_a[10] ^ input_a[0]);
  assign popcount36_pgij_core_112 = input_a[2] & input_a[26];
  assign popcount36_pgij_core_113 = ~(input_a[23] & input_a[34]);
  assign popcount36_pgij_core_114 = ~(input_a[22] & input_a[13]);
  assign popcount36_pgij_core_115 = ~input_a[14];
  assign popcount36_pgij_core_116 = ~input_a[26];
  assign popcount36_pgij_core_118 = ~(input_a[12] ^ input_a[29]);
  assign popcount36_pgij_core_120 = input_a[26] ^ input_a[10];
  assign popcount36_pgij_core_121 = input_a[34] & input_a[5];
  assign popcount36_pgij_core_122 = input_a[5] ^ input_a[2];
  assign popcount36_pgij_core_123 = input_a[8] | input_a[16];
  assign popcount36_pgij_core_124 = input_a[13] & input_a[7];
  assign popcount36_pgij_core_125 = input_a[2] | input_a[12];
  assign popcount36_pgij_core_127 = input_a[16] | input_a[9];
  assign popcount36_pgij_core_128 = input_a[34] | input_a[22];
  assign popcount36_pgij_core_129 = input_a[16] ^ popcount36_pgij_core_115;
  assign popcount36_pgij_core_130 = input_a[14] ^ input_a[33];
  assign popcount36_pgij_core_131 = ~popcount36_pgij_core_129;
  assign popcount36_pgij_core_133 = input_a[16] | popcount36_pgij_core_129;
  assign popcount36_pgij_core_134 = ~(input_a[21] & input_a[34]);
  assign popcount36_pgij_core_135 = input_a[20] ^ input_a[1];
  assign popcount36_pgij_core_136 = input_a[16] | popcount36_pgij_core_133;
  assign popcount36_pgij_core_137 = ~(input_a[15] | input_a[33]);
  assign popcount36_pgij_core_141 = ~(input_a[1] | input_a[5]);
  assign popcount36_pgij_core_143 = ~(input_a[13] | input_a[32]);
  assign popcount36_pgij_core_144 = ~(input_a[20] ^ input_a[8]);
  assign popcount36_pgij_core_146 = ~(input_a[16] | input_a[28]);
  assign popcount36_pgij_core_147 = input_a[17] & input_a[4];
  assign popcount36_pgij_core_148 = input_a[4] & input_a[28];
  assign popcount36_pgij_core_149 = ~(input_a[26] ^ input_a[32]);
  assign popcount36_pgij_core_150 = ~(input_a[4] ^ input_a[30]);
  assign popcount36_pgij_core_153 = ~(input_a[24] ^ input_a[8]);
  assign popcount36_pgij_core_154 = input_a[10] | input_a[26];
  assign popcount36_pgij_core_155 = ~(input_a[28] | input_a[2]);
  assign popcount36_pgij_core_156 = input_a[27] | input_a[1];
  assign popcount36_pgij_core_158 = ~(input_a[2] & input_a[30]);
  assign popcount36_pgij_core_159 = input_a[4] ^ input_a[30];
  assign popcount36_pgij_core_160 = ~(input_a[18] ^ input_a[7]);
  assign popcount36_pgij_core_165 = input_a[5] ^ input_a[14];
  assign popcount36_pgij_core_166 = ~input_a[17];
  assign popcount36_pgij_core_167 = ~(input_a[15] & input_a[30]);
  assign popcount36_pgij_core_168 = ~(input_a[22] & input_a[15]);
  assign popcount36_pgij_core_169 = ~(input_a[1] & input_a[34]);
  assign popcount36_pgij_core_170 = input_a[7] | input_a[19];
  assign popcount36_pgij_core_171 = input_a[27] & input_a[15];
  assign popcount36_pgij_core_172 = input_a[34] | input_a[13];
  assign popcount36_pgij_core_173 = ~(input_a[12] & input_a[26]);
  assign popcount36_pgij_core_174 = input_a[3] & input_a[26];
  assign popcount36_pgij_core_175 = ~(input_a[10] ^ input_a[9]);
  assign popcount36_pgij_core_178 = input_a[25] & input_a[10];
  assign popcount36_pgij_core_179 = ~input_a[15];
  assign popcount36_pgij_core_180_not = ~input_a[1];
  assign popcount36_pgij_core_181 = ~(input_a[28] ^ input_a[9]);
  assign popcount36_pgij_core_185 = input_a[7] & input_a[35];
  assign popcount36_pgij_core_186 = ~input_a[14];
  assign popcount36_pgij_core_187 = input_a[27] ^ input_a[3];
  assign popcount36_pgij_core_188 = ~input_a[18];
  assign popcount36_pgij_core_189 = ~input_a[1];
  assign popcount36_pgij_core_193_not = ~input_a[14];
  assign popcount36_pgij_core_194 = ~(input_a[35] & input_a[8]);
  assign popcount36_pgij_core_196 = ~input_a[11];
  assign popcount36_pgij_core_197 = input_a[28] ^ input_a[30];
  assign popcount36_pgij_core_198 = ~(input_a[26] ^ input_a[9]);
  assign popcount36_pgij_core_199 = input_a[30] ^ input_a[13];
  assign popcount36_pgij_core_201 = ~(input_a[12] | input_a[5]);
  assign popcount36_pgij_core_202 = ~(input_a[25] | input_a[17]);
  assign popcount36_pgij_core_203 = ~(input_a[10] & input_a[23]);
  assign popcount36_pgij_core_204 = input_a[5] | input_a[9];
  assign popcount36_pgij_core_205 = ~(input_a[33] ^ input_a[18]);
  assign popcount36_pgij_core_207 = ~(input_a[2] | input_a[6]);
  assign popcount36_pgij_core_208 = input_a[8] | input_a[13];
  assign popcount36_pgij_core_209 = ~(input_a[3] ^ input_a[9]);
  assign popcount36_pgij_core_213 = ~(input_a[19] & input_a[26]);
  assign popcount36_pgij_core_215 = ~(input_a[22] & input_a[1]);
  assign popcount36_pgij_core_216 = input_a[16] | input_a[4];
  assign popcount36_pgij_core_217 = ~input_a[17];
  assign popcount36_pgij_core_218_not = ~input_a[28];
  assign popcount36_pgij_core_219 = ~(input_a[20] | input_a[9]);
  assign popcount36_pgij_core_223 = ~input_a[29];
  assign popcount36_pgij_core_225 = input_a[17] & input_a[22];
  assign popcount36_pgij_core_227 = ~(input_a[29] & input_a[12]);
  assign popcount36_pgij_core_231 = ~(input_a[11] | input_a[33]);
  assign popcount36_pgij_core_232 = ~input_a[16];
  assign popcount36_pgij_core_233 = input_a[18] ^ input_a[25];
  assign popcount36_pgij_core_234 = input_a[33] | input_a[25];
  assign popcount36_pgij_core_235 = ~(input_a[15] & input_a[35]);
  assign popcount36_pgij_core_237 = input_a[7] ^ popcount36_pgij_core_234;
  assign popcount36_pgij_core_238 = input_a[7] & popcount36_pgij_core_234;
  assign popcount36_pgij_core_239 = input_a[14] | popcount36_pgij_core_238;
  assign popcount36_pgij_core_241 = input_a[4] ^ input_a[14];
  assign popcount36_pgij_core_242 = input_a[14] | popcount36_pgij_core_239;
  assign popcount36_pgij_core_243 = ~(input_a[20] ^ input_a[18]);
  assign popcount36_pgij_core_244 = input_a[14] & input_a[29];
  assign popcount36_pgij_core_247 = ~(input_a[11] & input_a[7]);
  assign popcount36_pgij_core_249 = ~(input_a[8] & input_a[27]);
  assign popcount36_pgij_core_250 = input_a[5] ^ input_a[32];
  assign popcount36_pgij_core_251 = input_a[11] & input_a[34];
  assign popcount36_pgij_core_252 = ~(input_a[31] | input_a[2]);
  assign popcount36_pgij_core_255 = input_a[9] & popcount36_pgij_core_251;
  assign popcount36_pgij_core_256 = popcount36_pgij_core_232 | popcount36_pgij_core_255;
  assign popcount36_pgij_core_257 = popcount36_pgij_core_131 | popcount36_pgij_core_237;
  assign popcount36_pgij_core_258 = popcount36_pgij_core_131 & popcount36_pgij_core_237;
  assign popcount36_pgij_core_259 = ~(popcount36_pgij_core_257 & popcount36_pgij_core_256);
  assign popcount36_pgij_core_260 = popcount36_pgij_core_257 & popcount36_pgij_core_256;
  assign popcount36_pgij_core_261 = popcount36_pgij_core_258 | popcount36_pgij_core_260;
  assign popcount36_pgij_core_262 = ~(popcount36_pgij_core_136 & popcount36_pgij_core_242);
  assign popcount36_pgij_core_264 = popcount36_pgij_core_262 ^ popcount36_pgij_core_261;
  assign popcount36_pgij_core_265 = popcount36_pgij_core_262 & popcount36_pgij_core_261;
  assign popcount36_pgij_core_266 = input_a[14] | popcount36_pgij_core_265;
  assign popcount36_pgij_core_267 = ~input_a[29];
  assign popcount36_pgij_core_268 = ~(input_a[2] ^ input_a[16]);
  assign popcount36_pgij_core_269 = input_a[7] | popcount36_pgij_core_266;
  assign popcount36_pgij_core_270 = input_a[16] & input_a[34];
  assign popcount36_pgij_core_272 = ~(input_a[32] | input_a[22]);
  assign popcount36_pgij_core_273 = input_a[15] ^ input_a[25];
  assign popcount36_pgij_core_274 = ~(input_a[15] & input_a[22]);
  assign popcount36_pgij_core_275 = ~(input_a[11] ^ input_a[19]);

  assign popcount36_pgij_out[0] = input_a[0];
  assign popcount36_pgij_out[1] = 1'b0;
  assign popcount36_pgij_out[2] = popcount36_pgij_core_259;
  assign popcount36_pgij_out[3] = popcount36_pgij_core_264;
  assign popcount36_pgij_out[4] = popcount36_pgij_core_269;
  assign popcount36_pgij_out[5] = 1'b0;
endmodule