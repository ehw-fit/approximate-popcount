// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.63243
// WCE=19.0
// EP=0.928879%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_ue9l(input [21:0] input_a, output [4:0] popcount22_ue9l_out);
  wire popcount22_ue9l_core_025;
  wire popcount22_ue9l_core_026;
  wire popcount22_ue9l_core_027;
  wire popcount22_ue9l_core_029;
  wire popcount22_ue9l_core_032;
  wire popcount22_ue9l_core_033;
  wire popcount22_ue9l_core_037;
  wire popcount22_ue9l_core_039;
  wire popcount22_ue9l_core_040;
  wire popcount22_ue9l_core_041;
  wire popcount22_ue9l_core_042;
  wire popcount22_ue9l_core_043;
  wire popcount22_ue9l_core_044;
  wire popcount22_ue9l_core_047;
  wire popcount22_ue9l_core_049;
  wire popcount22_ue9l_core_052;
  wire popcount22_ue9l_core_053;
  wire popcount22_ue9l_core_054;
  wire popcount22_ue9l_core_055;
  wire popcount22_ue9l_core_056;
  wire popcount22_ue9l_core_057;
  wire popcount22_ue9l_core_059;
  wire popcount22_ue9l_core_063;
  wire popcount22_ue9l_core_065;
  wire popcount22_ue9l_core_066;
  wire popcount22_ue9l_core_067;
  wire popcount22_ue9l_core_068;
  wire popcount22_ue9l_core_069;
  wire popcount22_ue9l_core_070;
  wire popcount22_ue9l_core_071;
  wire popcount22_ue9l_core_073;
  wire popcount22_ue9l_core_074;
  wire popcount22_ue9l_core_075;
  wire popcount22_ue9l_core_076;
  wire popcount22_ue9l_core_078;
  wire popcount22_ue9l_core_082;
  wire popcount22_ue9l_core_083;
  wire popcount22_ue9l_core_084;
  wire popcount22_ue9l_core_087;
  wire popcount22_ue9l_core_088;
  wire popcount22_ue9l_core_089;
  wire popcount22_ue9l_core_092;
  wire popcount22_ue9l_core_093;
  wire popcount22_ue9l_core_094;
  wire popcount22_ue9l_core_095;
  wire popcount22_ue9l_core_097;
  wire popcount22_ue9l_core_098_not;
  wire popcount22_ue9l_core_099;
  wire popcount22_ue9l_core_102;
  wire popcount22_ue9l_core_103;
  wire popcount22_ue9l_core_104;
  wire popcount22_ue9l_core_105;
  wire popcount22_ue9l_core_107;
  wire popcount22_ue9l_core_108;
  wire popcount22_ue9l_core_109;
  wire popcount22_ue9l_core_110;
  wire popcount22_ue9l_core_111;
  wire popcount22_ue9l_core_113_not;
  wire popcount22_ue9l_core_114;
  wire popcount22_ue9l_core_115;
  wire popcount22_ue9l_core_119;
  wire popcount22_ue9l_core_120;
  wire popcount22_ue9l_core_121;
  wire popcount22_ue9l_core_123;
  wire popcount22_ue9l_core_124;
  wire popcount22_ue9l_core_125;
  wire popcount22_ue9l_core_127;
  wire popcount22_ue9l_core_128;
  wire popcount22_ue9l_core_131;
  wire popcount22_ue9l_core_132;
  wire popcount22_ue9l_core_133;
  wire popcount22_ue9l_core_134;
  wire popcount22_ue9l_core_136;
  wire popcount22_ue9l_core_137;
  wire popcount22_ue9l_core_138;
  wire popcount22_ue9l_core_139;
  wire popcount22_ue9l_core_141;
  wire popcount22_ue9l_core_142;
  wire popcount22_ue9l_core_143;
  wire popcount22_ue9l_core_144;
  wire popcount22_ue9l_core_146;
  wire popcount22_ue9l_core_150;
  wire popcount22_ue9l_core_151;
  wire popcount22_ue9l_core_152;
  wire popcount22_ue9l_core_153;
  wire popcount22_ue9l_core_155;
  wire popcount22_ue9l_core_156;
  wire popcount22_ue9l_core_157;
  wire popcount22_ue9l_core_159;

  assign popcount22_ue9l_core_025 = input_a[2] ^ input_a[3];
  assign popcount22_ue9l_core_026 = input_a[14] ^ input_a[0];
  assign popcount22_ue9l_core_027 = ~(input_a[14] ^ input_a[18]);
  assign popcount22_ue9l_core_029 = input_a[19] | input_a[3];
  assign popcount22_ue9l_core_032 = input_a[14] | input_a[15];
  assign popcount22_ue9l_core_033 = ~(input_a[7] & input_a[9]);
  assign popcount22_ue9l_core_037 = ~(input_a[5] ^ input_a[19]);
  assign popcount22_ue9l_core_039 = input_a[7] | input_a[18];
  assign popcount22_ue9l_core_040 = ~(input_a[20] ^ input_a[19]);
  assign popcount22_ue9l_core_041 = ~(input_a[20] | input_a[12]);
  assign popcount22_ue9l_core_042 = ~(input_a[6] ^ input_a[16]);
  assign popcount22_ue9l_core_043 = ~(input_a[10] ^ input_a[5]);
  assign popcount22_ue9l_core_044 = ~input_a[16];
  assign popcount22_ue9l_core_047 = ~(input_a[6] ^ input_a[3]);
  assign popcount22_ue9l_core_049 = ~input_a[6];
  assign popcount22_ue9l_core_052 = ~(input_a[16] ^ input_a[11]);
  assign popcount22_ue9l_core_053 = ~(input_a[8] ^ input_a[19]);
  assign popcount22_ue9l_core_054 = ~(input_a[0] | input_a[7]);
  assign popcount22_ue9l_core_055 = ~input_a[6];
  assign popcount22_ue9l_core_056 = input_a[8] ^ input_a[1];
  assign popcount22_ue9l_core_057 = ~(input_a[16] | input_a[16]);
  assign popcount22_ue9l_core_059 = input_a[0] & input_a[0];
  assign popcount22_ue9l_core_063 = ~(input_a[3] & input_a[15]);
  assign popcount22_ue9l_core_065 = ~(input_a[14] | input_a[12]);
  assign popcount22_ue9l_core_066 = ~(input_a[6] ^ input_a[16]);
  assign popcount22_ue9l_core_067 = input_a[7] | input_a[6];
  assign popcount22_ue9l_core_068 = ~(input_a[12] ^ input_a[15]);
  assign popcount22_ue9l_core_069 = ~(input_a[10] & input_a[21]);
  assign popcount22_ue9l_core_070 = ~(input_a[9] & input_a[1]);
  assign popcount22_ue9l_core_071 = input_a[18] & input_a[15];
  assign popcount22_ue9l_core_073 = input_a[2] ^ input_a[6];
  assign popcount22_ue9l_core_074 = ~(input_a[2] ^ input_a[13]);
  assign popcount22_ue9l_core_075 = ~input_a[4];
  assign popcount22_ue9l_core_076 = ~(input_a[16] ^ input_a[9]);
  assign popcount22_ue9l_core_078 = ~(input_a[17] & input_a[5]);
  assign popcount22_ue9l_core_082 = ~(input_a[17] ^ input_a[11]);
  assign popcount22_ue9l_core_083 = ~(input_a[10] & input_a[2]);
  assign popcount22_ue9l_core_084 = input_a[18] & input_a[6];
  assign popcount22_ue9l_core_087 = ~(input_a[20] ^ input_a[19]);
  assign popcount22_ue9l_core_088 = input_a[2] & input_a[16];
  assign popcount22_ue9l_core_089 = ~input_a[4];
  assign popcount22_ue9l_core_092 = ~(input_a[11] | input_a[11]);
  assign popcount22_ue9l_core_093 = input_a[18] ^ input_a[2];
  assign popcount22_ue9l_core_094 = ~(input_a[5] & input_a[21]);
  assign popcount22_ue9l_core_095 = input_a[13] ^ input_a[17];
  assign popcount22_ue9l_core_097 = input_a[20] & input_a[17];
  assign popcount22_ue9l_core_098_not = ~input_a[0];
  assign popcount22_ue9l_core_099 = ~(input_a[1] | input_a[0]);
  assign popcount22_ue9l_core_102 = input_a[4] & input_a[21];
  assign popcount22_ue9l_core_103 = ~(input_a[10] ^ input_a[17]);
  assign popcount22_ue9l_core_104 = input_a[1] ^ input_a[16];
  assign popcount22_ue9l_core_105 = input_a[4] | input_a[12];
  assign popcount22_ue9l_core_107 = input_a[19] & input_a[7];
  assign popcount22_ue9l_core_108 = ~input_a[0];
  assign popcount22_ue9l_core_109 = ~(input_a[10] | input_a[11]);
  assign popcount22_ue9l_core_110 = ~(input_a[21] | input_a[2]);
  assign popcount22_ue9l_core_111 = ~(input_a[20] ^ input_a[18]);
  assign popcount22_ue9l_core_113_not = ~input_a[14];
  assign popcount22_ue9l_core_114 = input_a[21] | input_a[12];
  assign popcount22_ue9l_core_115 = ~(input_a[21] ^ input_a[16]);
  assign popcount22_ue9l_core_119 = ~(input_a[4] & input_a[11]);
  assign popcount22_ue9l_core_120 = ~(input_a[18] | input_a[0]);
  assign popcount22_ue9l_core_121 = input_a[4] ^ input_a[16];
  assign popcount22_ue9l_core_123 = ~(input_a[10] ^ input_a[4]);
  assign popcount22_ue9l_core_124 = input_a[19] | input_a[19];
  assign popcount22_ue9l_core_125 = ~input_a[19];
  assign popcount22_ue9l_core_127 = input_a[10] & input_a[16];
  assign popcount22_ue9l_core_128 = input_a[20] | input_a[18];
  assign popcount22_ue9l_core_131 = ~input_a[6];
  assign popcount22_ue9l_core_132 = ~(input_a[3] & input_a[4]);
  assign popcount22_ue9l_core_133 = ~(input_a[21] & input_a[0]);
  assign popcount22_ue9l_core_134 = input_a[1] & input_a[4];
  assign popcount22_ue9l_core_136 = ~(input_a[12] ^ input_a[13]);
  assign popcount22_ue9l_core_137 = ~(input_a[5] ^ input_a[4]);
  assign popcount22_ue9l_core_138 = ~(input_a[0] | input_a[6]);
  assign popcount22_ue9l_core_139 = input_a[14] ^ input_a[3];
  assign popcount22_ue9l_core_141 = ~input_a[19];
  assign popcount22_ue9l_core_142 = input_a[8] | input_a[1];
  assign popcount22_ue9l_core_143 = ~(input_a[2] | input_a[17]);
  assign popcount22_ue9l_core_144 = input_a[19] ^ input_a[17];
  assign popcount22_ue9l_core_146 = input_a[6] | input_a[13];
  assign popcount22_ue9l_core_150 = ~(input_a[19] & input_a[0]);
  assign popcount22_ue9l_core_151 = input_a[9] ^ input_a[0];
  assign popcount22_ue9l_core_152 = ~(input_a[20] ^ input_a[12]);
  assign popcount22_ue9l_core_153 = ~input_a[9];
  assign popcount22_ue9l_core_155 = ~(input_a[3] | input_a[18]);
  assign popcount22_ue9l_core_156 = ~(input_a[0] & input_a[4]);
  assign popcount22_ue9l_core_157 = ~(input_a[7] & input_a[15]);
  assign popcount22_ue9l_core_159 = ~(input_a[7] ^ input_a[3]);

  assign popcount22_ue9l_out[0] = input_a[4];
  assign popcount22_ue9l_out[1] = 1'b0;
  assign popcount22_ue9l_out[2] = input_a[2];
  assign popcount22_ue9l_out[3] = input_a[11];
  assign popcount22_ue9l_out[4] = 1'b0;
endmodule