// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=17.9084
// WCE=58.0
// EP=0.982627%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_fd46(input [38:0] input_a, output [5:0] popcount39_fd46_out);
  wire popcount39_fd46_core_041;
  wire popcount39_fd46_core_042;
  wire popcount39_fd46_core_043;
  wire popcount39_fd46_core_044_not;
  wire popcount39_fd46_core_045;
  wire popcount39_fd46_core_046;
  wire popcount39_fd46_core_047;
  wire popcount39_fd46_core_048;
  wire popcount39_fd46_core_049;
  wire popcount39_fd46_core_051;
  wire popcount39_fd46_core_053;
  wire popcount39_fd46_core_054;
  wire popcount39_fd46_core_055;
  wire popcount39_fd46_core_057;
  wire popcount39_fd46_core_059;
  wire popcount39_fd46_core_063;
  wire popcount39_fd46_core_064;
  wire popcount39_fd46_core_065_not;
  wire popcount39_fd46_core_066;
  wire popcount39_fd46_core_069;
  wire popcount39_fd46_core_070;
  wire popcount39_fd46_core_072;
  wire popcount39_fd46_core_074;
  wire popcount39_fd46_core_075;
  wire popcount39_fd46_core_076;
  wire popcount39_fd46_core_077;
  wire popcount39_fd46_core_078;
  wire popcount39_fd46_core_079;
  wire popcount39_fd46_core_080;
  wire popcount39_fd46_core_081;
  wire popcount39_fd46_core_082;
  wire popcount39_fd46_core_083;
  wire popcount39_fd46_core_084_not;
  wire popcount39_fd46_core_085;
  wire popcount39_fd46_core_089;
  wire popcount39_fd46_core_091;
  wire popcount39_fd46_core_092;
  wire popcount39_fd46_core_093;
  wire popcount39_fd46_core_094;
  wire popcount39_fd46_core_095;
  wire popcount39_fd46_core_096;
  wire popcount39_fd46_core_097;
  wire popcount39_fd46_core_098;
  wire popcount39_fd46_core_099;
  wire popcount39_fd46_core_100;
  wire popcount39_fd46_core_101;
  wire popcount39_fd46_core_102;
  wire popcount39_fd46_core_103;
  wire popcount39_fd46_core_104;
  wire popcount39_fd46_core_106;
  wire popcount39_fd46_core_107_not;
  wire popcount39_fd46_core_109;
  wire popcount39_fd46_core_110;
  wire popcount39_fd46_core_111;
  wire popcount39_fd46_core_113;
  wire popcount39_fd46_core_114;
  wire popcount39_fd46_core_115;
  wire popcount39_fd46_core_116;
  wire popcount39_fd46_core_117;
  wire popcount39_fd46_core_118;
  wire popcount39_fd46_core_119;
  wire popcount39_fd46_core_120;
  wire popcount39_fd46_core_122;
  wire popcount39_fd46_core_123;
  wire popcount39_fd46_core_126;
  wire popcount39_fd46_core_127;
  wire popcount39_fd46_core_128;
  wire popcount39_fd46_core_130;
  wire popcount39_fd46_core_131;
  wire popcount39_fd46_core_133;
  wire popcount39_fd46_core_136;
  wire popcount39_fd46_core_137;
  wire popcount39_fd46_core_139;
  wire popcount39_fd46_core_140;
  wire popcount39_fd46_core_141;
  wire popcount39_fd46_core_142;
  wire popcount39_fd46_core_146;
  wire popcount39_fd46_core_148;
  wire popcount39_fd46_core_149;
  wire popcount39_fd46_core_151;
  wire popcount39_fd46_core_152;
  wire popcount39_fd46_core_154;
  wire popcount39_fd46_core_156;
  wire popcount39_fd46_core_157;
  wire popcount39_fd46_core_159;
  wire popcount39_fd46_core_160;
  wire popcount39_fd46_core_163;
  wire popcount39_fd46_core_165;
  wire popcount39_fd46_core_167;
  wire popcount39_fd46_core_168;
  wire popcount39_fd46_core_170;
  wire popcount39_fd46_core_171;
  wire popcount39_fd46_core_173;
  wire popcount39_fd46_core_174;
  wire popcount39_fd46_core_175;
  wire popcount39_fd46_core_176;
  wire popcount39_fd46_core_180;
  wire popcount39_fd46_core_182;
  wire popcount39_fd46_core_183;
  wire popcount39_fd46_core_184;
  wire popcount39_fd46_core_185;
  wire popcount39_fd46_core_187;
  wire popcount39_fd46_core_189;
  wire popcount39_fd46_core_191;
  wire popcount39_fd46_core_192;
  wire popcount39_fd46_core_194;
  wire popcount39_fd46_core_196;
  wire popcount39_fd46_core_197;
  wire popcount39_fd46_core_198;
  wire popcount39_fd46_core_200;
  wire popcount39_fd46_core_202;
  wire popcount39_fd46_core_203;
  wire popcount39_fd46_core_204;
  wire popcount39_fd46_core_205;
  wire popcount39_fd46_core_206;
  wire popcount39_fd46_core_215;
  wire popcount39_fd46_core_216;
  wire popcount39_fd46_core_217;
  wire popcount39_fd46_core_218;
  wire popcount39_fd46_core_220;
  wire popcount39_fd46_core_221;
  wire popcount39_fd46_core_224;
  wire popcount39_fd46_core_226;
  wire popcount39_fd46_core_227;
  wire popcount39_fd46_core_228;
  wire popcount39_fd46_core_229;
  wire popcount39_fd46_core_231;
  wire popcount39_fd46_core_232;
  wire popcount39_fd46_core_234;
  wire popcount39_fd46_core_235;
  wire popcount39_fd46_core_236;
  wire popcount39_fd46_core_237;
  wire popcount39_fd46_core_239;
  wire popcount39_fd46_core_241;
  wire popcount39_fd46_core_242;
  wire popcount39_fd46_core_243;
  wire popcount39_fd46_core_244;
  wire popcount39_fd46_core_246;
  wire popcount39_fd46_core_247;
  wire popcount39_fd46_core_248_not;
  wire popcount39_fd46_core_250;
  wire popcount39_fd46_core_252;
  wire popcount39_fd46_core_253;
  wire popcount39_fd46_core_254;
  wire popcount39_fd46_core_255;
  wire popcount39_fd46_core_259;
  wire popcount39_fd46_core_261;
  wire popcount39_fd46_core_262;
  wire popcount39_fd46_core_263;
  wire popcount39_fd46_core_264;
  wire popcount39_fd46_core_265;
  wire popcount39_fd46_core_266;
  wire popcount39_fd46_core_268;
  wire popcount39_fd46_core_269;
  wire popcount39_fd46_core_270;
  wire popcount39_fd46_core_271;
  wire popcount39_fd46_core_272;
  wire popcount39_fd46_core_274;
  wire popcount39_fd46_core_279;
  wire popcount39_fd46_core_281;
  wire popcount39_fd46_core_283;
  wire popcount39_fd46_core_285;
  wire popcount39_fd46_core_286;
  wire popcount39_fd46_core_287;
  wire popcount39_fd46_core_290;
  wire popcount39_fd46_core_291;
  wire popcount39_fd46_core_292;
  wire popcount39_fd46_core_293;
  wire popcount39_fd46_core_294;
  wire popcount39_fd46_core_298;
  wire popcount39_fd46_core_300;
  wire popcount39_fd46_core_303;
  wire popcount39_fd46_core_304;
  wire popcount39_fd46_core_305;
  wire popcount39_fd46_core_306;

  assign popcount39_fd46_core_041 = input_a[7] ^ input_a[10];
  assign popcount39_fd46_core_042 = input_a[28] & input_a[4];
  assign popcount39_fd46_core_043 = input_a[35] ^ input_a[0];
  assign popcount39_fd46_core_044_not = ~input_a[29];
  assign popcount39_fd46_core_045 = ~(input_a[31] | input_a[22]);
  assign popcount39_fd46_core_046 = ~(input_a[21] | input_a[18]);
  assign popcount39_fd46_core_047 = input_a[33] | input_a[38];
  assign popcount39_fd46_core_048 = input_a[12] ^ input_a[2];
  assign popcount39_fd46_core_049 = ~(input_a[28] ^ input_a[11]);
  assign popcount39_fd46_core_051 = input_a[34] | input_a[5];
  assign popcount39_fd46_core_053 = ~(input_a[34] & input_a[19]);
  assign popcount39_fd46_core_054 = ~input_a[21];
  assign popcount39_fd46_core_055 = ~(input_a[18] | input_a[12]);
  assign popcount39_fd46_core_057 = ~(input_a[32] & input_a[23]);
  assign popcount39_fd46_core_059 = ~(input_a[36] ^ input_a[27]);
  assign popcount39_fd46_core_063 = input_a[19] ^ input_a[2];
  assign popcount39_fd46_core_064 = input_a[38] | input_a[4];
  assign popcount39_fd46_core_065_not = ~input_a[28];
  assign popcount39_fd46_core_066 = ~(input_a[4] ^ input_a[31]);
  assign popcount39_fd46_core_069 = ~input_a[2];
  assign popcount39_fd46_core_070 = input_a[2] & input_a[8];
  assign popcount39_fd46_core_072 = input_a[37] ^ input_a[11];
  assign popcount39_fd46_core_074 = ~(input_a[5] & input_a[18]);
  assign popcount39_fd46_core_075 = ~input_a[33];
  assign popcount39_fd46_core_076 = ~(input_a[3] & input_a[10]);
  assign popcount39_fd46_core_077 = ~(input_a[26] & input_a[6]);
  assign popcount39_fd46_core_078 = input_a[32] | input_a[22];
  assign popcount39_fd46_core_079 = input_a[18] & input_a[21];
  assign popcount39_fd46_core_080 = input_a[32] | input_a[7];
  assign popcount39_fd46_core_081 = input_a[34] & input_a[18];
  assign popcount39_fd46_core_082 = ~(input_a[13] | input_a[32]);
  assign popcount39_fd46_core_083 = ~(input_a[16] & input_a[18]);
  assign popcount39_fd46_core_084_not = ~input_a[19];
  assign popcount39_fd46_core_085 = input_a[19] | input_a[1];
  assign popcount39_fd46_core_089 = ~(input_a[10] & input_a[3]);
  assign popcount39_fd46_core_091 = input_a[19] ^ input_a[22];
  assign popcount39_fd46_core_092 = ~(input_a[23] & input_a[10]);
  assign popcount39_fd46_core_093 = input_a[10] ^ input_a[18];
  assign popcount39_fd46_core_094 = ~(input_a[2] | input_a[10]);
  assign popcount39_fd46_core_095 = input_a[3] & input_a[7];
  assign popcount39_fd46_core_096 = input_a[38] | input_a[28];
  assign popcount39_fd46_core_097 = ~(input_a[0] & input_a[36]);
  assign popcount39_fd46_core_098 = input_a[24] | input_a[1];
  assign popcount39_fd46_core_099 = input_a[10] ^ input_a[20];
  assign popcount39_fd46_core_100 = ~input_a[3];
  assign popcount39_fd46_core_101 = ~(input_a[27] | input_a[5]);
  assign popcount39_fd46_core_102 = input_a[18] & input_a[17];
  assign popcount39_fd46_core_103 = ~(input_a[33] | input_a[0]);
  assign popcount39_fd46_core_104 = input_a[5] & input_a[5];
  assign popcount39_fd46_core_106 = ~(input_a[30] ^ input_a[9]);
  assign popcount39_fd46_core_107_not = ~input_a[7];
  assign popcount39_fd46_core_109 = ~(input_a[3] | input_a[6]);
  assign popcount39_fd46_core_110 = ~input_a[9];
  assign popcount39_fd46_core_111 = input_a[21] & input_a[11];
  assign popcount39_fd46_core_113 = input_a[11] & input_a[17];
  assign popcount39_fd46_core_114 = ~input_a[34];
  assign popcount39_fd46_core_115 = input_a[6] ^ input_a[38];
  assign popcount39_fd46_core_116 = input_a[19] & input_a[26];
  assign popcount39_fd46_core_117 = input_a[28] | input_a[4];
  assign popcount39_fd46_core_118 = ~(input_a[12] & input_a[24]);
  assign popcount39_fd46_core_119 = ~(input_a[3] | input_a[15]);
  assign popcount39_fd46_core_120 = ~(input_a[0] ^ input_a[29]);
  assign popcount39_fd46_core_122 = input_a[2] | input_a[24];
  assign popcount39_fd46_core_123 = ~input_a[38];
  assign popcount39_fd46_core_126 = input_a[7] | input_a[23];
  assign popcount39_fd46_core_127 = ~(input_a[11] & input_a[32]);
  assign popcount39_fd46_core_128 = input_a[12] | input_a[2];
  assign popcount39_fd46_core_130 = input_a[31] | input_a[18];
  assign popcount39_fd46_core_131 = ~(input_a[22] | input_a[1]);
  assign popcount39_fd46_core_133 = ~input_a[38];
  assign popcount39_fd46_core_136 = input_a[32] | input_a[9];
  assign popcount39_fd46_core_137 = ~(input_a[27] ^ input_a[0]);
  assign popcount39_fd46_core_139 = ~(input_a[2] | input_a[20]);
  assign popcount39_fd46_core_140 = ~(input_a[8] & input_a[27]);
  assign popcount39_fd46_core_141 = ~input_a[14];
  assign popcount39_fd46_core_142 = input_a[9] ^ input_a[8];
  assign popcount39_fd46_core_146 = input_a[28] & input_a[21];
  assign popcount39_fd46_core_148 = input_a[33] | input_a[4];
  assign popcount39_fd46_core_149 = ~input_a[34];
  assign popcount39_fd46_core_151 = ~(input_a[4] | input_a[31]);
  assign popcount39_fd46_core_152 = ~(input_a[16] ^ input_a[0]);
  assign popcount39_fd46_core_154 = input_a[29] ^ input_a[34];
  assign popcount39_fd46_core_156 = ~(input_a[33] & input_a[16]);
  assign popcount39_fd46_core_157 = ~input_a[35];
  assign popcount39_fd46_core_159 = input_a[26] & input_a[25];
  assign popcount39_fd46_core_160 = ~(input_a[33] & input_a[24]);
  assign popcount39_fd46_core_163 = ~(input_a[30] | input_a[7]);
  assign popcount39_fd46_core_165 = ~(input_a[20] & input_a[19]);
  assign popcount39_fd46_core_167 = ~(input_a[36] | input_a[31]);
  assign popcount39_fd46_core_168 = ~(input_a[4] ^ input_a[13]);
  assign popcount39_fd46_core_170 = input_a[3] & input_a[10];
  assign popcount39_fd46_core_171 = ~(input_a[2] & input_a[34]);
  assign popcount39_fd46_core_173 = ~(input_a[8] | input_a[16]);
  assign popcount39_fd46_core_174 = ~(input_a[38] & input_a[22]);
  assign popcount39_fd46_core_175 = input_a[18] & input_a[37];
  assign popcount39_fd46_core_176 = input_a[2] | input_a[32];
  assign popcount39_fd46_core_180 = ~(input_a[23] & input_a[21]);
  assign popcount39_fd46_core_182 = ~input_a[34];
  assign popcount39_fd46_core_183 = ~(input_a[16] ^ input_a[26]);
  assign popcount39_fd46_core_184 = input_a[16] | input_a[19];
  assign popcount39_fd46_core_185 = input_a[14] | input_a[11];
  assign popcount39_fd46_core_187 = ~(input_a[22] | input_a[8]);
  assign popcount39_fd46_core_189 = input_a[31] | input_a[8];
  assign popcount39_fd46_core_191 = input_a[28] | input_a[27];
  assign popcount39_fd46_core_192 = ~(input_a[17] | input_a[7]);
  assign popcount39_fd46_core_194 = ~(input_a[5] ^ input_a[8]);
  assign popcount39_fd46_core_196 = input_a[7] ^ input_a[27];
  assign popcount39_fd46_core_197 = ~(input_a[16] & input_a[31]);
  assign popcount39_fd46_core_198 = ~input_a[0];
  assign popcount39_fd46_core_200 = ~(input_a[10] | input_a[31]);
  assign popcount39_fd46_core_202 = input_a[27] ^ input_a[21];
  assign popcount39_fd46_core_203 = input_a[16] | input_a[35];
  assign popcount39_fd46_core_204 = ~(input_a[31] | input_a[38]);
  assign popcount39_fd46_core_205 = ~input_a[13];
  assign popcount39_fd46_core_206 = input_a[33] | input_a[28];
  assign popcount39_fd46_core_215 = input_a[21] | input_a[7];
  assign popcount39_fd46_core_216 = ~input_a[5];
  assign popcount39_fd46_core_217 = ~input_a[35];
  assign popcount39_fd46_core_218 = input_a[0] & input_a[36];
  assign popcount39_fd46_core_220 = input_a[20] ^ input_a[38];
  assign popcount39_fd46_core_221 = input_a[15] | input_a[5];
  assign popcount39_fd46_core_224 = ~(input_a[9] | input_a[19]);
  assign popcount39_fd46_core_226 = input_a[12] & input_a[13];
  assign popcount39_fd46_core_227 = ~(input_a[37] | input_a[11]);
  assign popcount39_fd46_core_228 = ~(input_a[38] & input_a[20]);
  assign popcount39_fd46_core_229 = ~(input_a[14] | input_a[19]);
  assign popcount39_fd46_core_231 = input_a[8] | input_a[28];
  assign popcount39_fd46_core_232 = ~(input_a[2] & input_a[4]);
  assign popcount39_fd46_core_234 = ~(input_a[15] & input_a[29]);
  assign popcount39_fd46_core_235 = input_a[18] & input_a[29];
  assign popcount39_fd46_core_236 = ~(input_a[37] ^ input_a[8]);
  assign popcount39_fd46_core_237 = ~(input_a[19] | input_a[1]);
  assign popcount39_fd46_core_239 = ~(input_a[6] ^ input_a[21]);
  assign popcount39_fd46_core_241 = input_a[6] & input_a[8];
  assign popcount39_fd46_core_242 = input_a[19] ^ input_a[29];
  assign popcount39_fd46_core_243 = ~(input_a[28] & input_a[7]);
  assign popcount39_fd46_core_244 = ~(input_a[3] | input_a[28]);
  assign popcount39_fd46_core_246 = ~(input_a[37] & input_a[27]);
  assign popcount39_fd46_core_247 = ~(input_a[19] & input_a[31]);
  assign popcount39_fd46_core_248_not = ~input_a[7];
  assign popcount39_fd46_core_250 = input_a[27] ^ input_a[23];
  assign popcount39_fd46_core_252 = ~(input_a[36] | input_a[36]);
  assign popcount39_fd46_core_253 = ~(input_a[14] ^ input_a[32]);
  assign popcount39_fd46_core_254 = input_a[13] ^ input_a[22];
  assign popcount39_fd46_core_255 = ~(input_a[15] & input_a[23]);
  assign popcount39_fd46_core_259 = ~input_a[24];
  assign popcount39_fd46_core_261 = input_a[19] | input_a[1];
  assign popcount39_fd46_core_262 = ~(input_a[7] | input_a[3]);
  assign popcount39_fd46_core_263 = ~(input_a[28] ^ input_a[27]);
  assign popcount39_fd46_core_264 = ~(input_a[25] ^ input_a[1]);
  assign popcount39_fd46_core_265 = ~(input_a[23] ^ input_a[38]);
  assign popcount39_fd46_core_266 = ~(input_a[36] & input_a[36]);
  assign popcount39_fd46_core_268 = ~(input_a[1] & input_a[3]);
  assign popcount39_fd46_core_269 = ~input_a[13];
  assign popcount39_fd46_core_270 = ~(input_a[22] ^ input_a[3]);
  assign popcount39_fd46_core_271 = ~(input_a[29] | input_a[12]);
  assign popcount39_fd46_core_272 = ~(input_a[4] ^ input_a[10]);
  assign popcount39_fd46_core_274 = ~(input_a[8] & input_a[6]);
  assign popcount39_fd46_core_279 = input_a[10] & input_a[19];
  assign popcount39_fd46_core_281 = ~(input_a[32] ^ input_a[16]);
  assign popcount39_fd46_core_283 = ~input_a[15];
  assign popcount39_fd46_core_285 = input_a[36] ^ input_a[10];
  assign popcount39_fd46_core_286 = ~input_a[2];
  assign popcount39_fd46_core_287 = input_a[10] ^ input_a[8];
  assign popcount39_fd46_core_290 = ~input_a[29];
  assign popcount39_fd46_core_291 = ~(input_a[21] ^ input_a[17]);
  assign popcount39_fd46_core_292 = input_a[37] ^ input_a[10];
  assign popcount39_fd46_core_293 = ~(input_a[17] & input_a[4]);
  assign popcount39_fd46_core_294 = input_a[15] & input_a[23];
  assign popcount39_fd46_core_298 = ~(input_a[13] & input_a[35]);
  assign popcount39_fd46_core_300 = input_a[8] ^ input_a[2];
  assign popcount39_fd46_core_303 = ~(input_a[34] | input_a[28]);
  assign popcount39_fd46_core_304 = input_a[21] | input_a[38];
  assign popcount39_fd46_core_305 = ~(input_a[25] & input_a[23]);
  assign popcount39_fd46_core_306 = input_a[11] ^ input_a[2];

  assign popcount39_fd46_out[0] = 1'b1;
  assign popcount39_fd46_out[1] = 1'b0;
  assign popcount39_fd46_out[2] = input_a[37];
  assign popcount39_fd46_out[3] = input_a[0];
  assign popcount39_fd46_out[4] = input_a[1];
  assign popcount39_fd46_out[5] = 1'b0;
endmodule