// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.81602
// WCE=21.0
// EP=0.888866%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_ia07(input [38:0] input_a, output [5:0] popcount39_ia07_out);
  wire popcount39_ia07_core_041;
  wire popcount39_ia07_core_042;
  wire popcount39_ia07_core_043;
  wire popcount39_ia07_core_044;
  wire popcount39_ia07_core_046;
  wire popcount39_ia07_core_047;
  wire popcount39_ia07_core_048;
  wire popcount39_ia07_core_049;
  wire popcount39_ia07_core_050;
  wire popcount39_ia07_core_051;
  wire popcount39_ia07_core_052;
  wire popcount39_ia07_core_054;
  wire popcount39_ia07_core_055;
  wire popcount39_ia07_core_056;
  wire popcount39_ia07_core_057;
  wire popcount39_ia07_core_058;
  wire popcount39_ia07_core_059;
  wire popcount39_ia07_core_060_not;
  wire popcount39_ia07_core_061;
  wire popcount39_ia07_core_062;
  wire popcount39_ia07_core_063;
  wire popcount39_ia07_core_064;
  wire popcount39_ia07_core_065;
  wire popcount39_ia07_core_066;
  wire popcount39_ia07_core_068;
  wire popcount39_ia07_core_069;
  wire popcount39_ia07_core_070;
  wire popcount39_ia07_core_072;
  wire popcount39_ia07_core_074;
  wire popcount39_ia07_core_075;
  wire popcount39_ia07_core_076;
  wire popcount39_ia07_core_077;
  wire popcount39_ia07_core_078;
  wire popcount39_ia07_core_079;
  wire popcount39_ia07_core_080;
  wire popcount39_ia07_core_081;
  wire popcount39_ia07_core_084;
  wire popcount39_ia07_core_085;
  wire popcount39_ia07_core_086;
  wire popcount39_ia07_core_087;
  wire popcount39_ia07_core_088;
  wire popcount39_ia07_core_091;
  wire popcount39_ia07_core_093;
  wire popcount39_ia07_core_094;
  wire popcount39_ia07_core_097;
  wire popcount39_ia07_core_098;
  wire popcount39_ia07_core_100;
  wire popcount39_ia07_core_101;
  wire popcount39_ia07_core_102;
  wire popcount39_ia07_core_105;
  wire popcount39_ia07_core_106;
  wire popcount39_ia07_core_108;
  wire popcount39_ia07_core_110;
  wire popcount39_ia07_core_111;
  wire popcount39_ia07_core_112;
  wire popcount39_ia07_core_113;
  wire popcount39_ia07_core_114;
  wire popcount39_ia07_core_116;
  wire popcount39_ia07_core_117;
  wire popcount39_ia07_core_118;
  wire popcount39_ia07_core_119;
  wire popcount39_ia07_core_120;
  wire popcount39_ia07_core_121;
  wire popcount39_ia07_core_123;
  wire popcount39_ia07_core_124;
  wire popcount39_ia07_core_128;
  wire popcount39_ia07_core_129;
  wire popcount39_ia07_core_130;
  wire popcount39_ia07_core_131;
  wire popcount39_ia07_core_132;
  wire popcount39_ia07_core_133;
  wire popcount39_ia07_core_134;
  wire popcount39_ia07_core_135;
  wire popcount39_ia07_core_136;
  wire popcount39_ia07_core_137;
  wire popcount39_ia07_core_140;
  wire popcount39_ia07_core_142;
  wire popcount39_ia07_core_143;
  wire popcount39_ia07_core_144;
  wire popcount39_ia07_core_145;
  wire popcount39_ia07_core_146;
  wire popcount39_ia07_core_147;
  wire popcount39_ia07_core_149;
  wire popcount39_ia07_core_150;
  wire popcount39_ia07_core_151;
  wire popcount39_ia07_core_152;
  wire popcount39_ia07_core_154;
  wire popcount39_ia07_core_157;
  wire popcount39_ia07_core_160_not;
  wire popcount39_ia07_core_161;
  wire popcount39_ia07_core_165;
  wire popcount39_ia07_core_166;
  wire popcount39_ia07_core_168;
  wire popcount39_ia07_core_170;
  wire popcount39_ia07_core_171;
  wire popcount39_ia07_core_176;
  wire popcount39_ia07_core_177;
  wire popcount39_ia07_core_178;
  wire popcount39_ia07_core_182;
  wire popcount39_ia07_core_183;
  wire popcount39_ia07_core_185;
  wire popcount39_ia07_core_186;
  wire popcount39_ia07_core_187;
  wire popcount39_ia07_core_188;
  wire popcount39_ia07_core_191;
  wire popcount39_ia07_core_192_not;
  wire popcount39_ia07_core_195;
  wire popcount39_ia07_core_196;
  wire popcount39_ia07_core_198;
  wire popcount39_ia07_core_199;
  wire popcount39_ia07_core_201;
  wire popcount39_ia07_core_202;
  wire popcount39_ia07_core_204;
  wire popcount39_ia07_core_205;
  wire popcount39_ia07_core_206;
  wire popcount39_ia07_core_209;
  wire popcount39_ia07_core_210;
  wire popcount39_ia07_core_211;
  wire popcount39_ia07_core_213;
  wire popcount39_ia07_core_217;
  wire popcount39_ia07_core_218;
  wire popcount39_ia07_core_219;
  wire popcount39_ia07_core_220;
  wire popcount39_ia07_core_221;
  wire popcount39_ia07_core_225;
  wire popcount39_ia07_core_226;
  wire popcount39_ia07_core_227;
  wire popcount39_ia07_core_234;
  wire popcount39_ia07_core_235;
  wire popcount39_ia07_core_236;
  wire popcount39_ia07_core_237;
  wire popcount39_ia07_core_239;
  wire popcount39_ia07_core_242;
  wire popcount39_ia07_core_243;
  wire popcount39_ia07_core_244;
  wire popcount39_ia07_core_245;
  wire popcount39_ia07_core_246;
  wire popcount39_ia07_core_247;
  wire popcount39_ia07_core_248;
  wire popcount39_ia07_core_250;
  wire popcount39_ia07_core_251;
  wire popcount39_ia07_core_252;
  wire popcount39_ia07_core_255;
  wire popcount39_ia07_core_257;
  wire popcount39_ia07_core_260;
  wire popcount39_ia07_core_262;
  wire popcount39_ia07_core_263;
  wire popcount39_ia07_core_264;
  wire popcount39_ia07_core_267;
  wire popcount39_ia07_core_269;
  wire popcount39_ia07_core_273;
  wire popcount39_ia07_core_274;
  wire popcount39_ia07_core_275;
  wire popcount39_ia07_core_276;
  wire popcount39_ia07_core_277;
  wire popcount39_ia07_core_280;
  wire popcount39_ia07_core_282;
  wire popcount39_ia07_core_284;
  wire popcount39_ia07_core_288_not;
  wire popcount39_ia07_core_291;
  wire popcount39_ia07_core_293;
  wire popcount39_ia07_core_295;
  wire popcount39_ia07_core_296;
  wire popcount39_ia07_core_298;
  wire popcount39_ia07_core_301;
  wire popcount39_ia07_core_302;

  assign popcount39_ia07_core_041 = input_a[13] & input_a[2];
  assign popcount39_ia07_core_042 = input_a[20] | input_a[3];
  assign popcount39_ia07_core_043 = input_a[19] | input_a[7];
  assign popcount39_ia07_core_044 = input_a[27] & input_a[25];
  assign popcount39_ia07_core_046 = ~(input_a[18] & input_a[14]);
  assign popcount39_ia07_core_047 = input_a[30] | input_a[22];
  assign popcount39_ia07_core_048 = input_a[5] ^ input_a[20];
  assign popcount39_ia07_core_049 = input_a[37] ^ input_a[2];
  assign popcount39_ia07_core_050 = ~(input_a[15] | input_a[24]);
  assign popcount39_ia07_core_051 = input_a[33] & input_a[12];
  assign popcount39_ia07_core_052 = ~input_a[36];
  assign popcount39_ia07_core_054 = input_a[0] | input_a[25];
  assign popcount39_ia07_core_055 = ~input_a[26];
  assign popcount39_ia07_core_056 = input_a[32] | input_a[3];
  assign popcount39_ia07_core_057 = input_a[5] & input_a[15];
  assign popcount39_ia07_core_058 = input_a[17] ^ input_a[1];
  assign popcount39_ia07_core_059 = ~input_a[9];
  assign popcount39_ia07_core_060_not = ~input_a[5];
  assign popcount39_ia07_core_061 = input_a[21] ^ input_a[19];
  assign popcount39_ia07_core_062 = input_a[38] | input_a[7];
  assign popcount39_ia07_core_063 = input_a[33] & input_a[23];
  assign popcount39_ia07_core_064 = ~(input_a[29] ^ input_a[38]);
  assign popcount39_ia07_core_065 = input_a[11] | input_a[34];
  assign popcount39_ia07_core_066 = input_a[24] ^ input_a[18];
  assign popcount39_ia07_core_068 = ~(input_a[17] & input_a[36]);
  assign popcount39_ia07_core_069 = input_a[5] | input_a[32];
  assign popcount39_ia07_core_070 = input_a[1] ^ input_a[25];
  assign popcount39_ia07_core_072 = ~(input_a[27] | input_a[29]);
  assign popcount39_ia07_core_074 = input_a[8] ^ input_a[18];
  assign popcount39_ia07_core_075 = ~(input_a[37] & input_a[2]);
  assign popcount39_ia07_core_076 = input_a[26] | input_a[12];
  assign popcount39_ia07_core_077 = input_a[3] & input_a[38];
  assign popcount39_ia07_core_078 = ~(input_a[24] & input_a[18]);
  assign popcount39_ia07_core_079 = ~(input_a[29] | input_a[11]);
  assign popcount39_ia07_core_080 = input_a[38] ^ input_a[18];
  assign popcount39_ia07_core_081 = input_a[25] & input_a[19];
  assign popcount39_ia07_core_084 = ~input_a[2];
  assign popcount39_ia07_core_085 = input_a[31] & input_a[7];
  assign popcount39_ia07_core_086 = ~(input_a[0] ^ input_a[13]);
  assign popcount39_ia07_core_087 = input_a[7] | input_a[1];
  assign popcount39_ia07_core_088 = ~input_a[11];
  assign popcount39_ia07_core_091 = ~(input_a[10] | input_a[25]);
  assign popcount39_ia07_core_093 = ~(input_a[9] ^ input_a[24]);
  assign popcount39_ia07_core_094 = ~(input_a[9] | input_a[20]);
  assign popcount39_ia07_core_097 = input_a[23] | input_a[29];
  assign popcount39_ia07_core_098 = input_a[33] ^ input_a[33];
  assign popcount39_ia07_core_100 = ~(input_a[31] & input_a[24]);
  assign popcount39_ia07_core_101 = ~(input_a[37] & input_a[18]);
  assign popcount39_ia07_core_102 = input_a[2] ^ input_a[25];
  assign popcount39_ia07_core_105 = input_a[22] ^ input_a[6];
  assign popcount39_ia07_core_106 = ~(input_a[7] | input_a[12]);
  assign popcount39_ia07_core_108 = input_a[15] | input_a[9];
  assign popcount39_ia07_core_110 = ~(input_a[9] | input_a[16]);
  assign popcount39_ia07_core_111 = ~input_a[14];
  assign popcount39_ia07_core_112 = ~(input_a[36] ^ input_a[35]);
  assign popcount39_ia07_core_113 = ~input_a[25];
  assign popcount39_ia07_core_114 = ~(input_a[2] ^ input_a[37]);
  assign popcount39_ia07_core_116 = input_a[24] | input_a[29];
  assign popcount39_ia07_core_117 = ~(input_a[4] | input_a[27]);
  assign popcount39_ia07_core_118 = input_a[12] & input_a[19];
  assign popcount39_ia07_core_119 = input_a[6] ^ input_a[12];
  assign popcount39_ia07_core_120 = ~input_a[29];
  assign popcount39_ia07_core_121 = ~(input_a[20] | input_a[13]);
  assign popcount39_ia07_core_123 = ~input_a[21];
  assign popcount39_ia07_core_124 = ~input_a[36];
  assign popcount39_ia07_core_128 = ~(input_a[27] ^ input_a[4]);
  assign popcount39_ia07_core_129 = input_a[35] ^ input_a[2];
  assign popcount39_ia07_core_130 = input_a[18] & input_a[31];
  assign popcount39_ia07_core_131 = ~(input_a[11] ^ input_a[6]);
  assign popcount39_ia07_core_132 = ~(input_a[11] ^ input_a[24]);
  assign popcount39_ia07_core_133 = ~(input_a[3] & input_a[4]);
  assign popcount39_ia07_core_134 = ~(input_a[25] & input_a[33]);
  assign popcount39_ia07_core_135 = ~(input_a[29] & input_a[32]);
  assign popcount39_ia07_core_136 = input_a[2] & input_a[12];
  assign popcount39_ia07_core_137 = ~(input_a[13] & input_a[23]);
  assign popcount39_ia07_core_140 = ~(input_a[36] ^ input_a[31]);
  assign popcount39_ia07_core_142 = input_a[2] | input_a[2];
  assign popcount39_ia07_core_143 = input_a[10] ^ input_a[1];
  assign popcount39_ia07_core_144 = ~(input_a[2] | input_a[30]);
  assign popcount39_ia07_core_145 = input_a[22] & input_a[21];
  assign popcount39_ia07_core_146 = ~(input_a[28] | input_a[2]);
  assign popcount39_ia07_core_147 = input_a[37] & input_a[28];
  assign popcount39_ia07_core_149 = input_a[36] & input_a[23];
  assign popcount39_ia07_core_150 = input_a[15] ^ input_a[1];
  assign popcount39_ia07_core_151 = input_a[1] | input_a[34];
  assign popcount39_ia07_core_152 = ~(input_a[25] | input_a[8]);
  assign popcount39_ia07_core_154 = ~input_a[21];
  assign popcount39_ia07_core_157 = input_a[28] ^ input_a[6];
  assign popcount39_ia07_core_160_not = ~input_a[32];
  assign popcount39_ia07_core_161 = ~(input_a[9] & input_a[3]);
  assign popcount39_ia07_core_165 = ~(input_a[15] & input_a[35]);
  assign popcount39_ia07_core_166 = ~input_a[21];
  assign popcount39_ia07_core_168 = ~(input_a[12] & input_a[24]);
  assign popcount39_ia07_core_170 = input_a[21] | input_a[27];
  assign popcount39_ia07_core_171 = input_a[28] ^ input_a[9];
  assign popcount39_ia07_core_176 = ~(input_a[4] ^ input_a[12]);
  assign popcount39_ia07_core_177 = ~(input_a[35] | input_a[36]);
  assign popcount39_ia07_core_178 = ~(input_a[34] & input_a[8]);
  assign popcount39_ia07_core_182 = input_a[1] & input_a[27];
  assign popcount39_ia07_core_183 = ~(input_a[21] | input_a[30]);
  assign popcount39_ia07_core_185 = ~input_a[21];
  assign popcount39_ia07_core_186 = ~(input_a[11] & input_a[38]);
  assign popcount39_ia07_core_187 = ~(input_a[8] | input_a[30]);
  assign popcount39_ia07_core_188 = ~input_a[22];
  assign popcount39_ia07_core_191 = input_a[24] & input_a[20];
  assign popcount39_ia07_core_192_not = ~input_a[1];
  assign popcount39_ia07_core_195 = ~(input_a[16] | input_a[21]);
  assign popcount39_ia07_core_196 = ~(input_a[6] | input_a[27]);
  assign popcount39_ia07_core_198 = ~(input_a[6] | input_a[16]);
  assign popcount39_ia07_core_199 = input_a[19] & input_a[26];
  assign popcount39_ia07_core_201 = input_a[3] | input_a[25];
  assign popcount39_ia07_core_202 = ~input_a[8];
  assign popcount39_ia07_core_204 = ~(input_a[16] | input_a[12]);
  assign popcount39_ia07_core_205 = input_a[37] | input_a[25];
  assign popcount39_ia07_core_206 = ~(input_a[14] & input_a[20]);
  assign popcount39_ia07_core_209 = input_a[4] & input_a[27];
  assign popcount39_ia07_core_210 = input_a[10] ^ input_a[2];
  assign popcount39_ia07_core_211 = input_a[21] | input_a[38];
  assign popcount39_ia07_core_213 = ~(input_a[21] ^ input_a[0]);
  assign popcount39_ia07_core_217 = ~input_a[6];
  assign popcount39_ia07_core_218 = ~input_a[6];
  assign popcount39_ia07_core_219 = ~input_a[14];
  assign popcount39_ia07_core_220 = ~(input_a[1] | input_a[11]);
  assign popcount39_ia07_core_221 = input_a[2] & input_a[20];
  assign popcount39_ia07_core_225 = ~input_a[20];
  assign popcount39_ia07_core_226 = ~(input_a[13] | input_a[38]);
  assign popcount39_ia07_core_227 = input_a[34] | input_a[27];
  assign popcount39_ia07_core_234 = ~(input_a[36] ^ input_a[36]);
  assign popcount39_ia07_core_235 = ~input_a[14];
  assign popcount39_ia07_core_236 = ~(input_a[36] | input_a[35]);
  assign popcount39_ia07_core_237 = input_a[9] & input_a[24];
  assign popcount39_ia07_core_239 = input_a[20] ^ input_a[27];
  assign popcount39_ia07_core_242 = ~(input_a[17] & input_a[38]);
  assign popcount39_ia07_core_243 = input_a[28] ^ input_a[37];
  assign popcount39_ia07_core_244 = input_a[25] & input_a[12];
  assign popcount39_ia07_core_245 = ~(input_a[32] | input_a[28]);
  assign popcount39_ia07_core_246 = ~(input_a[36] ^ input_a[15]);
  assign popcount39_ia07_core_247 = ~input_a[22];
  assign popcount39_ia07_core_248 = input_a[9] | input_a[18];
  assign popcount39_ia07_core_250 = ~(input_a[23] | input_a[22]);
  assign popcount39_ia07_core_251 = ~(input_a[22] | input_a[9]);
  assign popcount39_ia07_core_252 = input_a[20] | input_a[4];
  assign popcount39_ia07_core_255 = input_a[25] | input_a[16];
  assign popcount39_ia07_core_257 = input_a[30] ^ input_a[9];
  assign popcount39_ia07_core_260 = ~(input_a[31] ^ input_a[9]);
  assign popcount39_ia07_core_262 = input_a[34] ^ input_a[14];
  assign popcount39_ia07_core_263 = input_a[25] | input_a[23];
  assign popcount39_ia07_core_264 = input_a[37] ^ input_a[28];
  assign popcount39_ia07_core_267 = ~(input_a[9] | input_a[4]);
  assign popcount39_ia07_core_269 = ~(input_a[9] & input_a[16]);
  assign popcount39_ia07_core_273 = ~(input_a[5] & input_a[38]);
  assign popcount39_ia07_core_274 = input_a[6] & input_a[4];
  assign popcount39_ia07_core_275 = ~(input_a[37] | input_a[19]);
  assign popcount39_ia07_core_276 = input_a[10] & input_a[14];
  assign popcount39_ia07_core_277 = ~(input_a[14] & input_a[31]);
  assign popcount39_ia07_core_280 = input_a[35] & input_a[9];
  assign popcount39_ia07_core_282 = ~input_a[1];
  assign popcount39_ia07_core_284 = input_a[23] ^ input_a[5];
  assign popcount39_ia07_core_288_not = ~input_a[29];
  assign popcount39_ia07_core_291 = ~(input_a[2] & input_a[9]);
  assign popcount39_ia07_core_293 = input_a[17] ^ input_a[24];
  assign popcount39_ia07_core_295 = ~(input_a[17] | input_a[3]);
  assign popcount39_ia07_core_296 = input_a[8] | input_a[37];
  assign popcount39_ia07_core_298 = input_a[4] | input_a[26];
  assign popcount39_ia07_core_301 = ~(input_a[12] | input_a[29]);
  assign popcount39_ia07_core_302 = ~(input_a[17] & input_a[38]);

  assign popcount39_ia07_out[0] = input_a[23];
  assign popcount39_ia07_out[1] = 1'b1;
  assign popcount39_ia07_out[2] = input_a[28];
  assign popcount39_ia07_out[3] = 1'b0;
  assign popcount39_ia07_out[4] = 1'b1;
  assign popcount39_ia07_out[5] = 1'b0;
endmodule