// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=11.7369
// WCE=42.0
// EP=0.969712%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount45_dcjf(input [44:0] input_a, output [5:0] popcount45_dcjf_out);
  wire popcount45_dcjf_core_047;
  wire popcount45_dcjf_core_049;
  wire popcount45_dcjf_core_050;
  wire popcount45_dcjf_core_054;
  wire popcount45_dcjf_core_055;
  wire popcount45_dcjf_core_057;
  wire popcount45_dcjf_core_058;
  wire popcount45_dcjf_core_060;
  wire popcount45_dcjf_core_061;
  wire popcount45_dcjf_core_062;
  wire popcount45_dcjf_core_063;
  wire popcount45_dcjf_core_064;
  wire popcount45_dcjf_core_065;
  wire popcount45_dcjf_core_067;
  wire popcount45_dcjf_core_068;
  wire popcount45_dcjf_core_069;
  wire popcount45_dcjf_core_072;
  wire popcount45_dcjf_core_073;
  wire popcount45_dcjf_core_074;
  wire popcount45_dcjf_core_075;
  wire popcount45_dcjf_core_077;
  wire popcount45_dcjf_core_078;
  wire popcount45_dcjf_core_080;
  wire popcount45_dcjf_core_081;
  wire popcount45_dcjf_core_083;
  wire popcount45_dcjf_core_086;
  wire popcount45_dcjf_core_087;
  wire popcount45_dcjf_core_091;
  wire popcount45_dcjf_core_093;
  wire popcount45_dcjf_core_094;
  wire popcount45_dcjf_core_095;
  wire popcount45_dcjf_core_099;
  wire popcount45_dcjf_core_100;
  wire popcount45_dcjf_core_101;
  wire popcount45_dcjf_core_102;
  wire popcount45_dcjf_core_103;
  wire popcount45_dcjf_core_104;
  wire popcount45_dcjf_core_105;
  wire popcount45_dcjf_core_106;
  wire popcount45_dcjf_core_109;
  wire popcount45_dcjf_core_110;
  wire popcount45_dcjf_core_111;
  wire popcount45_dcjf_core_113;
  wire popcount45_dcjf_core_114;
  wire popcount45_dcjf_core_116;
  wire popcount45_dcjf_core_117;
  wire popcount45_dcjf_core_118;
  wire popcount45_dcjf_core_119;
  wire popcount45_dcjf_core_121;
  wire popcount45_dcjf_core_123;
  wire popcount45_dcjf_core_124;
  wire popcount45_dcjf_core_125;
  wire popcount45_dcjf_core_126;
  wire popcount45_dcjf_core_127;
  wire popcount45_dcjf_core_129;
  wire popcount45_dcjf_core_130;
  wire popcount45_dcjf_core_133;
  wire popcount45_dcjf_core_135;
  wire popcount45_dcjf_core_139;
  wire popcount45_dcjf_core_141;
  wire popcount45_dcjf_core_142;
  wire popcount45_dcjf_core_143;
  wire popcount45_dcjf_core_144;
  wire popcount45_dcjf_core_145;
  wire popcount45_dcjf_core_146;
  wire popcount45_dcjf_core_150;
  wire popcount45_dcjf_core_152;
  wire popcount45_dcjf_core_153;
  wire popcount45_dcjf_core_155;
  wire popcount45_dcjf_core_156;
  wire popcount45_dcjf_core_157;
  wire popcount45_dcjf_core_159;
  wire popcount45_dcjf_core_160;
  wire popcount45_dcjf_core_161;
  wire popcount45_dcjf_core_162;
  wire popcount45_dcjf_core_163;
  wire popcount45_dcjf_core_164;
  wire popcount45_dcjf_core_165;
  wire popcount45_dcjf_core_167;
  wire popcount45_dcjf_core_168;
  wire popcount45_dcjf_core_169;
  wire popcount45_dcjf_core_172;
  wire popcount45_dcjf_core_173;
  wire popcount45_dcjf_core_174;
  wire popcount45_dcjf_core_176;
  wire popcount45_dcjf_core_177;
  wire popcount45_dcjf_core_180;
  wire popcount45_dcjf_core_181;
  wire popcount45_dcjf_core_182;
  wire popcount45_dcjf_core_183;
  wire popcount45_dcjf_core_185;
  wire popcount45_dcjf_core_186;
  wire popcount45_dcjf_core_187;
  wire popcount45_dcjf_core_188;
  wire popcount45_dcjf_core_191;
  wire popcount45_dcjf_core_195;
  wire popcount45_dcjf_core_197;
  wire popcount45_dcjf_core_198;
  wire popcount45_dcjf_core_199;
  wire popcount45_dcjf_core_200;
  wire popcount45_dcjf_core_201;
  wire popcount45_dcjf_core_202;
  wire popcount45_dcjf_core_203;
  wire popcount45_dcjf_core_204;
  wire popcount45_dcjf_core_205;
  wire popcount45_dcjf_core_206;
  wire popcount45_dcjf_core_207;
  wire popcount45_dcjf_core_208;
  wire popcount45_dcjf_core_211;
  wire popcount45_dcjf_core_212;
  wire popcount45_dcjf_core_214;
  wire popcount45_dcjf_core_216;
  wire popcount45_dcjf_core_217;
  wire popcount45_dcjf_core_220;
  wire popcount45_dcjf_core_221;
  wire popcount45_dcjf_core_222;
  wire popcount45_dcjf_core_225;
  wire popcount45_dcjf_core_226;
  wire popcount45_dcjf_core_227;
  wire popcount45_dcjf_core_229;
  wire popcount45_dcjf_core_230;
  wire popcount45_dcjf_core_231;
  wire popcount45_dcjf_core_232;
  wire popcount45_dcjf_core_234;
  wire popcount45_dcjf_core_236;
  wire popcount45_dcjf_core_238;
  wire popcount45_dcjf_core_240;
  wire popcount45_dcjf_core_242;
  wire popcount45_dcjf_core_248;
  wire popcount45_dcjf_core_249;
  wire popcount45_dcjf_core_250;
  wire popcount45_dcjf_core_252;
  wire popcount45_dcjf_core_254_not;
  wire popcount45_dcjf_core_255;
  wire popcount45_dcjf_core_256;
  wire popcount45_dcjf_core_258;
  wire popcount45_dcjf_core_259;
  wire popcount45_dcjf_core_260;
  wire popcount45_dcjf_core_262;
  wire popcount45_dcjf_core_264;
  wire popcount45_dcjf_core_265;
  wire popcount45_dcjf_core_266;
  wire popcount45_dcjf_core_267;
  wire popcount45_dcjf_core_268;
  wire popcount45_dcjf_core_270;
  wire popcount45_dcjf_core_272;
  wire popcount45_dcjf_core_273;
  wire popcount45_dcjf_core_274;
  wire popcount45_dcjf_core_275;
  wire popcount45_dcjf_core_276;
  wire popcount45_dcjf_core_277;
  wire popcount45_dcjf_core_278;
  wire popcount45_dcjf_core_279;
  wire popcount45_dcjf_core_280;
  wire popcount45_dcjf_core_282;
  wire popcount45_dcjf_core_283;
  wire popcount45_dcjf_core_285;
  wire popcount45_dcjf_core_286;
  wire popcount45_dcjf_core_288;
  wire popcount45_dcjf_core_289;
  wire popcount45_dcjf_core_292;
  wire popcount45_dcjf_core_294;
  wire popcount45_dcjf_core_299;
  wire popcount45_dcjf_core_300;
  wire popcount45_dcjf_core_301;
  wire popcount45_dcjf_core_303;
  wire popcount45_dcjf_core_305;
  wire popcount45_dcjf_core_306;
  wire popcount45_dcjf_core_307_not;
  wire popcount45_dcjf_core_308;
  wire popcount45_dcjf_core_309;
  wire popcount45_dcjf_core_311_not;
  wire popcount45_dcjf_core_312;
  wire popcount45_dcjf_core_313;
  wire popcount45_dcjf_core_315;
  wire popcount45_dcjf_core_320;
  wire popcount45_dcjf_core_322;
  wire popcount45_dcjf_core_323;
  wire popcount45_dcjf_core_324;
  wire popcount45_dcjf_core_325;
  wire popcount45_dcjf_core_326;
  wire popcount45_dcjf_core_327;
  wire popcount45_dcjf_core_329;
  wire popcount45_dcjf_core_331;
  wire popcount45_dcjf_core_333;
  wire popcount45_dcjf_core_334;
  wire popcount45_dcjf_core_335;
  wire popcount45_dcjf_core_336;
  wire popcount45_dcjf_core_338;
  wire popcount45_dcjf_core_339;
  wire popcount45_dcjf_core_340;
  wire popcount45_dcjf_core_341;
  wire popcount45_dcjf_core_342;
  wire popcount45_dcjf_core_343;
  wire popcount45_dcjf_core_344;
  wire popcount45_dcjf_core_345;
  wire popcount45_dcjf_core_346;
  wire popcount45_dcjf_core_348;
  wire popcount45_dcjf_core_349;
  wire popcount45_dcjf_core_350;
  wire popcount45_dcjf_core_352;
  wire popcount45_dcjf_core_354;
  wire popcount45_dcjf_core_355;

  assign popcount45_dcjf_core_047 = ~(input_a[33] & input_a[30]);
  assign popcount45_dcjf_core_049 = input_a[17] ^ input_a[5];
  assign popcount45_dcjf_core_050 = input_a[0] | input_a[5];
  assign popcount45_dcjf_core_054 = ~(input_a[35] | input_a[7]);
  assign popcount45_dcjf_core_055 = ~(input_a[3] | input_a[5]);
  assign popcount45_dcjf_core_057 = ~input_a[40];
  assign popcount45_dcjf_core_058 = ~(input_a[14] & input_a[35]);
  assign popcount45_dcjf_core_060 = ~(input_a[4] ^ input_a[22]);
  assign popcount45_dcjf_core_061 = input_a[13] ^ input_a[40];
  assign popcount45_dcjf_core_062 = input_a[20] | input_a[20];
  assign popcount45_dcjf_core_063 = ~(input_a[17] | input_a[41]);
  assign popcount45_dcjf_core_064 = ~input_a[20];
  assign popcount45_dcjf_core_065 = input_a[23] | input_a[19];
  assign popcount45_dcjf_core_067 = ~(input_a[19] ^ input_a[13]);
  assign popcount45_dcjf_core_068 = input_a[5] | input_a[9];
  assign popcount45_dcjf_core_069 = ~(input_a[6] & input_a[24]);
  assign popcount45_dcjf_core_072 = input_a[16] & input_a[21];
  assign popcount45_dcjf_core_073 = ~(input_a[37] | input_a[21]);
  assign popcount45_dcjf_core_074 = ~(input_a[36] | input_a[24]);
  assign popcount45_dcjf_core_075 = ~(input_a[19] ^ input_a[35]);
  assign popcount45_dcjf_core_077 = input_a[43] & input_a[1];
  assign popcount45_dcjf_core_078 = input_a[39] ^ input_a[26];
  assign popcount45_dcjf_core_080 = ~input_a[3];
  assign popcount45_dcjf_core_081 = input_a[13] ^ input_a[43];
  assign popcount45_dcjf_core_083 = ~input_a[40];
  assign popcount45_dcjf_core_086 = input_a[41] | input_a[0];
  assign popcount45_dcjf_core_087 = ~input_a[36];
  assign popcount45_dcjf_core_091 = input_a[20] & input_a[16];
  assign popcount45_dcjf_core_093 = ~input_a[38];
  assign popcount45_dcjf_core_094 = ~(input_a[31] | input_a[41]);
  assign popcount45_dcjf_core_095 = ~(input_a[18] | input_a[18]);
  assign popcount45_dcjf_core_099 = input_a[1] | input_a[43];
  assign popcount45_dcjf_core_100 = ~(input_a[34] ^ input_a[29]);
  assign popcount45_dcjf_core_101 = ~input_a[30];
  assign popcount45_dcjf_core_102 = input_a[13] ^ input_a[7];
  assign popcount45_dcjf_core_103 = ~input_a[1];
  assign popcount45_dcjf_core_104 = input_a[43] ^ input_a[9];
  assign popcount45_dcjf_core_105 = ~(input_a[5] | input_a[36]);
  assign popcount45_dcjf_core_106 = ~(input_a[43] | input_a[15]);
  assign popcount45_dcjf_core_109 = ~(input_a[1] | input_a[12]);
  assign popcount45_dcjf_core_110 = input_a[36] ^ input_a[31];
  assign popcount45_dcjf_core_111 = ~(input_a[14] & input_a[29]);
  assign popcount45_dcjf_core_113 = input_a[25] & input_a[14];
  assign popcount45_dcjf_core_114 = input_a[22] | input_a[33];
  assign popcount45_dcjf_core_116 = ~(input_a[3] ^ input_a[42]);
  assign popcount45_dcjf_core_117 = ~(input_a[12] ^ input_a[20]);
  assign popcount45_dcjf_core_118 = ~(input_a[22] ^ input_a[1]);
  assign popcount45_dcjf_core_119 = input_a[42] ^ input_a[6];
  assign popcount45_dcjf_core_121 = input_a[14] & input_a[23];
  assign popcount45_dcjf_core_123 = ~(input_a[24] | input_a[8]);
  assign popcount45_dcjf_core_124 = ~input_a[40];
  assign popcount45_dcjf_core_125 = input_a[21] & input_a[10];
  assign popcount45_dcjf_core_126 = input_a[23] | input_a[30];
  assign popcount45_dcjf_core_127 = ~(input_a[16] & input_a[6]);
  assign popcount45_dcjf_core_129 = ~(input_a[8] | input_a[14]);
  assign popcount45_dcjf_core_130 = ~(input_a[29] | input_a[41]);
  assign popcount45_dcjf_core_133 = ~input_a[36];
  assign popcount45_dcjf_core_135 = input_a[18] ^ input_a[19];
  assign popcount45_dcjf_core_139 = ~(input_a[26] ^ input_a[36]);
  assign popcount45_dcjf_core_141 = ~(input_a[44] & input_a[20]);
  assign popcount45_dcjf_core_142 = ~(input_a[43] | input_a[20]);
  assign popcount45_dcjf_core_143 = input_a[39] ^ input_a[16];
  assign popcount45_dcjf_core_144 = input_a[34] & input_a[41];
  assign popcount45_dcjf_core_145 = ~input_a[2];
  assign popcount45_dcjf_core_146 = ~(input_a[14] ^ input_a[17]);
  assign popcount45_dcjf_core_150 = input_a[16] | input_a[32];
  assign popcount45_dcjf_core_152 = input_a[16] ^ input_a[34];
  assign popcount45_dcjf_core_153 = ~(input_a[18] ^ input_a[14]);
  assign popcount45_dcjf_core_155 = ~(input_a[39] | input_a[38]);
  assign popcount45_dcjf_core_156 = ~(input_a[34] ^ input_a[2]);
  assign popcount45_dcjf_core_157 = ~input_a[25];
  assign popcount45_dcjf_core_159 = ~(input_a[24] | input_a[40]);
  assign popcount45_dcjf_core_160 = ~(input_a[33] | input_a[17]);
  assign popcount45_dcjf_core_161 = input_a[10] | input_a[38];
  assign popcount45_dcjf_core_162 = input_a[5] ^ input_a[44];
  assign popcount45_dcjf_core_163 = ~(input_a[2] ^ input_a[10]);
  assign popcount45_dcjf_core_164 = input_a[42] & input_a[29];
  assign popcount45_dcjf_core_165 = input_a[33] & input_a[14];
  assign popcount45_dcjf_core_167 = ~(input_a[36] ^ input_a[35]);
  assign popcount45_dcjf_core_168 = input_a[43] ^ input_a[14];
  assign popcount45_dcjf_core_169 = ~(input_a[18] & input_a[21]);
  assign popcount45_dcjf_core_172 = input_a[14] & input_a[41];
  assign popcount45_dcjf_core_173 = ~(input_a[32] & input_a[12]);
  assign popcount45_dcjf_core_174 = ~input_a[30];
  assign popcount45_dcjf_core_176 = ~(input_a[14] ^ input_a[39]);
  assign popcount45_dcjf_core_177 = input_a[21] ^ input_a[20];
  assign popcount45_dcjf_core_180 = ~(input_a[32] | input_a[35]);
  assign popcount45_dcjf_core_181 = input_a[5] & input_a[25];
  assign popcount45_dcjf_core_182 = input_a[1] ^ input_a[9];
  assign popcount45_dcjf_core_183 = input_a[0] | input_a[20];
  assign popcount45_dcjf_core_185 = ~(input_a[42] ^ input_a[27]);
  assign popcount45_dcjf_core_186 = ~input_a[20];
  assign popcount45_dcjf_core_187 = input_a[12] | input_a[23];
  assign popcount45_dcjf_core_188 = ~input_a[31];
  assign popcount45_dcjf_core_191 = ~(input_a[4] | input_a[5]);
  assign popcount45_dcjf_core_195 = ~input_a[36];
  assign popcount45_dcjf_core_197 = input_a[10] | input_a[33];
  assign popcount45_dcjf_core_198 = input_a[31] | input_a[44];
  assign popcount45_dcjf_core_199 = input_a[8] & input_a[32];
  assign popcount45_dcjf_core_200 = input_a[5] & input_a[30];
  assign popcount45_dcjf_core_201 = ~(input_a[41] ^ input_a[1]);
  assign popcount45_dcjf_core_202 = ~(input_a[10] & input_a[34]);
  assign popcount45_dcjf_core_203 = ~input_a[6];
  assign popcount45_dcjf_core_204 = ~input_a[44];
  assign popcount45_dcjf_core_205 = input_a[32] ^ input_a[2];
  assign popcount45_dcjf_core_206 = ~(input_a[19] ^ input_a[42]);
  assign popcount45_dcjf_core_207 = input_a[20] | input_a[12];
  assign popcount45_dcjf_core_208 = ~(input_a[26] & input_a[13]);
  assign popcount45_dcjf_core_211 = ~(input_a[31] | input_a[35]);
  assign popcount45_dcjf_core_212 = input_a[40] & input_a[10];
  assign popcount45_dcjf_core_214 = ~input_a[0];
  assign popcount45_dcjf_core_216 = input_a[22] & input_a[38];
  assign popcount45_dcjf_core_217 = ~(input_a[33] ^ input_a[24]);
  assign popcount45_dcjf_core_220 = ~(input_a[40] ^ input_a[41]);
  assign popcount45_dcjf_core_221 = ~(input_a[24] | input_a[40]);
  assign popcount45_dcjf_core_222 = input_a[26] | input_a[32];
  assign popcount45_dcjf_core_225 = ~input_a[3];
  assign popcount45_dcjf_core_226 = input_a[31] | input_a[8];
  assign popcount45_dcjf_core_227 = ~(input_a[12] ^ input_a[11]);
  assign popcount45_dcjf_core_229 = ~(input_a[4] | input_a[29]);
  assign popcount45_dcjf_core_230 = ~(input_a[33] | input_a[21]);
  assign popcount45_dcjf_core_231 = input_a[32] & input_a[19];
  assign popcount45_dcjf_core_232 = ~(input_a[16] & input_a[36]);
  assign popcount45_dcjf_core_234 = ~(input_a[14] | input_a[34]);
  assign popcount45_dcjf_core_236 = input_a[36] | input_a[2];
  assign popcount45_dcjf_core_238 = ~input_a[25];
  assign popcount45_dcjf_core_240 = ~(input_a[5] | input_a[12]);
  assign popcount45_dcjf_core_242 = ~(input_a[12] | input_a[3]);
  assign popcount45_dcjf_core_248 = ~(input_a[31] ^ input_a[14]);
  assign popcount45_dcjf_core_249 = ~(input_a[18] ^ input_a[42]);
  assign popcount45_dcjf_core_250 = ~input_a[2];
  assign popcount45_dcjf_core_252 = input_a[28] & input_a[31];
  assign popcount45_dcjf_core_254_not = ~input_a[40];
  assign popcount45_dcjf_core_255 = ~(input_a[15] | input_a[27]);
  assign popcount45_dcjf_core_256 = input_a[20] | input_a[25];
  assign popcount45_dcjf_core_258 = input_a[9] | input_a[1];
  assign popcount45_dcjf_core_259 = input_a[41] & input_a[37];
  assign popcount45_dcjf_core_260 = ~(input_a[32] | input_a[10]);
  assign popcount45_dcjf_core_262 = ~(input_a[17] ^ input_a[18]);
  assign popcount45_dcjf_core_264 = ~(input_a[14] ^ input_a[15]);
  assign popcount45_dcjf_core_265 = input_a[38] | input_a[14];
  assign popcount45_dcjf_core_266 = input_a[20] ^ input_a[17];
  assign popcount45_dcjf_core_267 = input_a[17] | input_a[31];
  assign popcount45_dcjf_core_268 = ~(input_a[41] & input_a[37]);
  assign popcount45_dcjf_core_270 = ~(input_a[10] | input_a[43]);
  assign popcount45_dcjf_core_272 = ~(input_a[16] ^ input_a[0]);
  assign popcount45_dcjf_core_273 = ~(input_a[8] & input_a[43]);
  assign popcount45_dcjf_core_274 = ~(input_a[44] & input_a[35]);
  assign popcount45_dcjf_core_275 = ~(input_a[21] ^ input_a[22]);
  assign popcount45_dcjf_core_276 = ~(input_a[0] & input_a[9]);
  assign popcount45_dcjf_core_277 = ~(input_a[36] & input_a[23]);
  assign popcount45_dcjf_core_278 = input_a[27] & input_a[14];
  assign popcount45_dcjf_core_279 = ~(input_a[1] ^ input_a[39]);
  assign popcount45_dcjf_core_280 = ~(input_a[35] | input_a[31]);
  assign popcount45_dcjf_core_282 = ~(input_a[9] & input_a[9]);
  assign popcount45_dcjf_core_283 = ~(input_a[1] ^ input_a[28]);
  assign popcount45_dcjf_core_285 = ~(input_a[43] & input_a[19]);
  assign popcount45_dcjf_core_286 = input_a[27] ^ input_a[6];
  assign popcount45_dcjf_core_288 = ~input_a[19];
  assign popcount45_dcjf_core_289 = ~(input_a[32] | input_a[25]);
  assign popcount45_dcjf_core_292 = input_a[27] ^ input_a[19];
  assign popcount45_dcjf_core_294 = ~input_a[12];
  assign popcount45_dcjf_core_299 = ~(input_a[9] | input_a[31]);
  assign popcount45_dcjf_core_300 = ~(input_a[17] ^ input_a[28]);
  assign popcount45_dcjf_core_301 = input_a[14] | input_a[5];
  assign popcount45_dcjf_core_303 = input_a[36] | input_a[40];
  assign popcount45_dcjf_core_305 = ~(input_a[24] ^ input_a[41]);
  assign popcount45_dcjf_core_306 = ~(input_a[38] | input_a[34]);
  assign popcount45_dcjf_core_307_not = ~input_a[13];
  assign popcount45_dcjf_core_308 = ~input_a[23];
  assign popcount45_dcjf_core_309 = input_a[8] ^ input_a[3];
  assign popcount45_dcjf_core_311_not = ~input_a[10];
  assign popcount45_dcjf_core_312 = ~(input_a[43] ^ input_a[2]);
  assign popcount45_dcjf_core_313 = ~(input_a[42] | input_a[39]);
  assign popcount45_dcjf_core_315 = ~input_a[40];
  assign popcount45_dcjf_core_320 = input_a[38] & input_a[13];
  assign popcount45_dcjf_core_322 = ~(input_a[20] ^ input_a[5]);
  assign popcount45_dcjf_core_323 = ~input_a[18];
  assign popcount45_dcjf_core_324 = input_a[14] | input_a[11];
  assign popcount45_dcjf_core_325 = ~input_a[11];
  assign popcount45_dcjf_core_326 = input_a[33] | input_a[31];
  assign popcount45_dcjf_core_327 = ~(input_a[14] | input_a[21]);
  assign popcount45_dcjf_core_329 = ~(input_a[25] & input_a[3]);
  assign popcount45_dcjf_core_331 = ~(input_a[32] | input_a[34]);
  assign popcount45_dcjf_core_333 = ~(input_a[35] ^ input_a[44]);
  assign popcount45_dcjf_core_334 = ~(input_a[0] | input_a[18]);
  assign popcount45_dcjf_core_335 = input_a[14] | input_a[4];
  assign popcount45_dcjf_core_336 = input_a[11] & input_a[42];
  assign popcount45_dcjf_core_338 = ~input_a[20];
  assign popcount45_dcjf_core_339 = ~(input_a[31] | input_a[19]);
  assign popcount45_dcjf_core_340 = ~input_a[27];
  assign popcount45_dcjf_core_341 = ~(input_a[8] & input_a[44]);
  assign popcount45_dcjf_core_342 = input_a[24] & input_a[4];
  assign popcount45_dcjf_core_343 = input_a[16] & input_a[12];
  assign popcount45_dcjf_core_344 = input_a[26] ^ input_a[0];
  assign popcount45_dcjf_core_345 = input_a[0] ^ input_a[27];
  assign popcount45_dcjf_core_346 = ~(input_a[31] | input_a[43]);
  assign popcount45_dcjf_core_348 = ~(input_a[33] ^ input_a[29]);
  assign popcount45_dcjf_core_349 = input_a[37] | input_a[13];
  assign popcount45_dcjf_core_350 = input_a[32] | input_a[42];
  assign popcount45_dcjf_core_352 = ~(input_a[27] | input_a[15]);
  assign popcount45_dcjf_core_354 = ~input_a[19];
  assign popcount45_dcjf_core_355 = ~(input_a[39] & input_a[22]);

  assign popcount45_dcjf_out[0] = 1'b1;
  assign popcount45_dcjf_out[1] = 1'b0;
  assign popcount45_dcjf_out[2] = input_a[44];
  assign popcount45_dcjf_out[3] = input_a[4];
  assign popcount45_dcjf_out[4] = input_a[4];
  assign popcount45_dcjf_out[5] = 1'b0;
endmodule