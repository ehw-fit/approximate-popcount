// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.11436
// WCE=11.0
// EP=0.855839%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount20_028g(input [19:0] input_a, output [4:0] popcount20_028g_out);
  wire popcount20_028g_core_022;
  wire popcount20_028g_core_023;
  wire popcount20_028g_core_027;
  wire popcount20_028g_core_028;
  wire popcount20_028g_core_029;
  wire popcount20_028g_core_030;
  wire popcount20_028g_core_031;
  wire popcount20_028g_core_035;
  wire popcount20_028g_core_037;
  wire popcount20_028g_core_038;
  wire popcount20_028g_core_039;
  wire popcount20_028g_core_044;
  wire popcount20_028g_core_046;
  wire popcount20_028g_core_049_not;
  wire popcount20_028g_core_053;
  wire popcount20_028g_core_054;
  wire popcount20_028g_core_055;
  wire popcount20_028g_core_059;
  wire popcount20_028g_core_060;
  wire popcount20_028g_core_061;
  wire popcount20_028g_core_062;
  wire popcount20_028g_core_063;
  wire popcount20_028g_core_064;
  wire popcount20_028g_core_065;
  wire popcount20_028g_core_066;
  wire popcount20_028g_core_067;
  wire popcount20_028g_core_068;
  wire popcount20_028g_core_071;
  wire popcount20_028g_core_072_not;
  wire popcount20_028g_core_074;
  wire popcount20_028g_core_075;
  wire popcount20_028g_core_077;
  wire popcount20_028g_core_079;
  wire popcount20_028g_core_080;
  wire popcount20_028g_core_083;
  wire popcount20_028g_core_084;
  wire popcount20_028g_core_085;
  wire popcount20_028g_core_087_not;
  wire popcount20_028g_core_088;
  wire popcount20_028g_core_089;
  wire popcount20_028g_core_090;
  wire popcount20_028g_core_091;
  wire popcount20_028g_core_094;
  wire popcount20_028g_core_095;
  wire popcount20_028g_core_096_not;
  wire popcount20_028g_core_098;
  wire popcount20_028g_core_100;
  wire popcount20_028g_core_102;
  wire popcount20_028g_core_103;
  wire popcount20_028g_core_104;
  wire popcount20_028g_core_106;
  wire popcount20_028g_core_107;
  wire popcount20_028g_core_109;
  wire popcount20_028g_core_110;
  wire popcount20_028g_core_111;
  wire popcount20_028g_core_112;
  wire popcount20_028g_core_119;
  wire popcount20_028g_core_120;
  wire popcount20_028g_core_123;
  wire popcount20_028g_core_124;
  wire popcount20_028g_core_125;
  wire popcount20_028g_core_126;
  wire popcount20_028g_core_128;
  wire popcount20_028g_core_129;
  wire popcount20_028g_core_130;
  wire popcount20_028g_core_132;
  wire popcount20_028g_core_133;
  wire popcount20_028g_core_136;
  wire popcount20_028g_core_137_not;
  wire popcount20_028g_core_139;
  wire popcount20_028g_core_140_not;
  wire popcount20_028g_core_141;
  wire popcount20_028g_core_142;
  wire popcount20_028g_core_143;
  wire popcount20_028g_core_144;

  assign popcount20_028g_core_022 = ~input_a[1];
  assign popcount20_028g_core_023 = input_a[12] ^ input_a[4];
  assign popcount20_028g_core_027 = ~(input_a[19] | input_a[3]);
  assign popcount20_028g_core_028 = ~(input_a[11] | input_a[19]);
  assign popcount20_028g_core_029 = input_a[1] & input_a[2];
  assign popcount20_028g_core_030 = ~input_a[19];
  assign popcount20_028g_core_031 = input_a[3] | input_a[6];
  assign popcount20_028g_core_035 = input_a[4] ^ input_a[16];
  assign popcount20_028g_core_037 = ~(input_a[9] | input_a[9]);
  assign popcount20_028g_core_038 = ~(input_a[13] | input_a[19]);
  assign popcount20_028g_core_039 = input_a[16] & input_a[2];
  assign popcount20_028g_core_044 = input_a[1] & input_a[4];
  assign popcount20_028g_core_046 = input_a[5] & input_a[7];
  assign popcount20_028g_core_049_not = ~input_a[2];
  assign popcount20_028g_core_053 = input_a[10] & input_a[19];
  assign popcount20_028g_core_054 = input_a[14] ^ input_a[1];
  assign popcount20_028g_core_055 = input_a[18] | input_a[17];
  assign popcount20_028g_core_059 = ~(input_a[15] & input_a[18]);
  assign popcount20_028g_core_060 = ~(input_a[14] | input_a[14]);
  assign popcount20_028g_core_061 = input_a[7] | input_a[2];
  assign popcount20_028g_core_062 = ~input_a[16];
  assign popcount20_028g_core_063 = ~input_a[2];
  assign popcount20_028g_core_064 = ~(input_a[6] & input_a[13]);
  assign popcount20_028g_core_065 = ~input_a[3];
  assign popcount20_028g_core_066 = input_a[4] & input_a[4];
  assign popcount20_028g_core_067 = input_a[7] | input_a[18];
  assign popcount20_028g_core_068 = input_a[16] & input_a[0];
  assign popcount20_028g_core_071 = input_a[17] & input_a[13];
  assign popcount20_028g_core_072_not = ~input_a[11];
  assign popcount20_028g_core_074 = input_a[1] & input_a[6];
  assign popcount20_028g_core_075 = ~(input_a[13] | input_a[19]);
  assign popcount20_028g_core_077 = ~input_a[4];
  assign popcount20_028g_core_079 = ~(input_a[7] ^ input_a[10]);
  assign popcount20_028g_core_080 = ~input_a[3];
  assign popcount20_028g_core_083 = ~(input_a[5] | input_a[8]);
  assign popcount20_028g_core_084 = input_a[9] ^ input_a[7];
  assign popcount20_028g_core_085 = input_a[1] ^ input_a[19];
  assign popcount20_028g_core_087_not = ~input_a[13];
  assign popcount20_028g_core_088 = ~input_a[14];
  assign popcount20_028g_core_089 = ~input_a[3];
  assign popcount20_028g_core_090 = ~(input_a[10] & input_a[5]);
  assign popcount20_028g_core_091 = input_a[18] & input_a[13];
  assign popcount20_028g_core_094 = ~(input_a[12] | input_a[1]);
  assign popcount20_028g_core_095 = input_a[2] ^ input_a[4];
  assign popcount20_028g_core_096_not = ~input_a[7];
  assign popcount20_028g_core_098 = ~(input_a[13] & input_a[12]);
  assign popcount20_028g_core_100 = ~(input_a[12] | input_a[11]);
  assign popcount20_028g_core_102 = input_a[9] ^ input_a[0];
  assign popcount20_028g_core_103 = input_a[16] & input_a[10];
  assign popcount20_028g_core_104 = input_a[4] | input_a[0];
  assign popcount20_028g_core_106 = input_a[0] | input_a[5];
  assign popcount20_028g_core_107 = ~(input_a[14] ^ input_a[14]);
  assign popcount20_028g_core_109 = ~input_a[18];
  assign popcount20_028g_core_110 = input_a[13] & input_a[10];
  assign popcount20_028g_core_111 = ~input_a[11];
  assign popcount20_028g_core_112 = ~input_a[1];
  assign popcount20_028g_core_119 = ~(input_a[13] ^ input_a[9]);
  assign popcount20_028g_core_120 = ~(input_a[15] | input_a[4]);
  assign popcount20_028g_core_123 = ~(input_a[13] & input_a[8]);
  assign popcount20_028g_core_124 = ~input_a[12];
  assign popcount20_028g_core_125 = ~(input_a[9] & input_a[0]);
  assign popcount20_028g_core_126 = ~(input_a[17] & input_a[2]);
  assign popcount20_028g_core_128 = ~input_a[6];
  assign popcount20_028g_core_129 = ~(input_a[5] ^ input_a[3]);
  assign popcount20_028g_core_130 = input_a[4] | input_a[11];
  assign popcount20_028g_core_132 = ~(input_a[12] & input_a[1]);
  assign popcount20_028g_core_133 = ~input_a[9];
  assign popcount20_028g_core_136 = ~input_a[18];
  assign popcount20_028g_core_137_not = ~input_a[19];
  assign popcount20_028g_core_139 = ~(input_a[18] & input_a[4]);
  assign popcount20_028g_core_140_not = ~input_a[13];
  assign popcount20_028g_core_141 = ~(input_a[14] & input_a[16]);
  assign popcount20_028g_core_142 = ~input_a[10];
  assign popcount20_028g_core_143 = ~(input_a[2] ^ input_a[8]);
  assign popcount20_028g_core_144 = input_a[14] & input_a[3];

  assign popcount20_028g_out[0] = input_a[13];
  assign popcount20_028g_out[1] = 1'b0;
  assign popcount20_028g_out[2] = 1'b0;
  assign popcount20_028g_out[3] = 1'b1;
  assign popcount20_028g_out[4] = 1'b0;
endmodule