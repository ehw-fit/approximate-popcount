// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=9.42559
// WCE=28.0
// EP=0.951022%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_43n0(input [21:0] input_a, output [4:0] popcount22_43n0_out);
  wire popcount22_43n0_core_024;
  wire popcount22_43n0_core_027;
  wire popcount22_43n0_core_028_not;
  wire popcount22_43n0_core_030;
  wire popcount22_43n0_core_031;
  wire popcount22_43n0_core_032;
  wire popcount22_43n0_core_033;
  wire popcount22_43n0_core_034;
  wire popcount22_43n0_core_036;
  wire popcount22_43n0_core_039;
  wire popcount22_43n0_core_042;
  wire popcount22_43n0_core_043;
  wire popcount22_43n0_core_044;
  wire popcount22_43n0_core_045;
  wire popcount22_43n0_core_046;
  wire popcount22_43n0_core_047;
  wire popcount22_43n0_core_048;
  wire popcount22_43n0_core_050;
  wire popcount22_43n0_core_053;
  wire popcount22_43n0_core_054;
  wire popcount22_43n0_core_055;
  wire popcount22_43n0_core_057;
  wire popcount22_43n0_core_058;
  wire popcount22_43n0_core_060;
  wire popcount22_43n0_core_061;
  wire popcount22_43n0_core_062;
  wire popcount22_43n0_core_064;
  wire popcount22_43n0_core_065;
  wire popcount22_43n0_core_068;
  wire popcount22_43n0_core_069;
  wire popcount22_43n0_core_071;
  wire popcount22_43n0_core_073;
  wire popcount22_43n0_core_074_not;
  wire popcount22_43n0_core_075;
  wire popcount22_43n0_core_077;
  wire popcount22_43n0_core_078;
  wire popcount22_43n0_core_079;
  wire popcount22_43n0_core_080;
  wire popcount22_43n0_core_081;
  wire popcount22_43n0_core_082;
  wire popcount22_43n0_core_085;
  wire popcount22_43n0_core_090;
  wire popcount22_43n0_core_092;
  wire popcount22_43n0_core_093;
  wire popcount22_43n0_core_094;
  wire popcount22_43n0_core_096;
  wire popcount22_43n0_core_097;
  wire popcount22_43n0_core_098;
  wire popcount22_43n0_core_100;
  wire popcount22_43n0_core_101;
  wire popcount22_43n0_core_102;
  wire popcount22_43n0_core_105;
  wire popcount22_43n0_core_107;
  wire popcount22_43n0_core_108;
  wire popcount22_43n0_core_109;
  wire popcount22_43n0_core_110;
  wire popcount22_43n0_core_113;
  wire popcount22_43n0_core_115;
  wire popcount22_43n0_core_116;
  wire popcount22_43n0_core_117_not;
  wire popcount22_43n0_core_118;
  wire popcount22_43n0_core_119;
  wire popcount22_43n0_core_124;
  wire popcount22_43n0_core_126;
  wire popcount22_43n0_core_130;
  wire popcount22_43n0_core_133;
  wire popcount22_43n0_core_134;
  wire popcount22_43n0_core_135;
  wire popcount22_43n0_core_137;
  wire popcount22_43n0_core_138;
  wire popcount22_43n0_core_139;
  wire popcount22_43n0_core_140;
  wire popcount22_43n0_core_141;
  wire popcount22_43n0_core_143;
  wire popcount22_43n0_core_144;
  wire popcount22_43n0_core_146;
  wire popcount22_43n0_core_147;
  wire popcount22_43n0_core_149;
  wire popcount22_43n0_core_152;
  wire popcount22_43n0_core_153;
  wire popcount22_43n0_core_156;
  wire popcount22_43n0_core_157;
  wire popcount22_43n0_core_159;
  wire popcount22_43n0_core_160;

  assign popcount22_43n0_core_024 = input_a[4] | input_a[20];
  assign popcount22_43n0_core_027 = input_a[2] | input_a[3];
  assign popcount22_43n0_core_028_not = ~input_a[7];
  assign popcount22_43n0_core_030 = input_a[17] ^ input_a[12];
  assign popcount22_43n0_core_031 = ~(input_a[6] & input_a[1]);
  assign popcount22_43n0_core_032 = input_a[13] | input_a[13];
  assign popcount22_43n0_core_033 = ~(input_a[11] & input_a[20]);
  assign popcount22_43n0_core_034 = input_a[12] & input_a[16];
  assign popcount22_43n0_core_036 = ~(input_a[8] & input_a[8]);
  assign popcount22_43n0_core_039 = input_a[14] & input_a[20];
  assign popcount22_43n0_core_042 = input_a[17] | input_a[18];
  assign popcount22_43n0_core_043 = ~(input_a[12] ^ input_a[6]);
  assign popcount22_43n0_core_044 = input_a[2] ^ input_a[14];
  assign popcount22_43n0_core_045 = ~(input_a[21] ^ input_a[14]);
  assign popcount22_43n0_core_046 = ~(input_a[4] & input_a[17]);
  assign popcount22_43n0_core_047 = ~(input_a[11] & input_a[18]);
  assign popcount22_43n0_core_048 = ~input_a[5];
  assign popcount22_43n0_core_050 = input_a[8] | input_a[3];
  assign popcount22_43n0_core_053 = ~(input_a[10] & input_a[1]);
  assign popcount22_43n0_core_054 = ~(input_a[17] | input_a[13]);
  assign popcount22_43n0_core_055 = input_a[21] | input_a[2];
  assign popcount22_43n0_core_057 = input_a[17] | input_a[0];
  assign popcount22_43n0_core_058 = input_a[10] ^ input_a[6];
  assign popcount22_43n0_core_060 = input_a[0] ^ input_a[7];
  assign popcount22_43n0_core_061 = input_a[12] ^ input_a[9];
  assign popcount22_43n0_core_062 = input_a[11] ^ input_a[12];
  assign popcount22_43n0_core_064 = ~(input_a[0] | input_a[7]);
  assign popcount22_43n0_core_065 = input_a[6] ^ input_a[6];
  assign popcount22_43n0_core_068 = ~input_a[11];
  assign popcount22_43n0_core_069 = ~(input_a[13] ^ input_a[18]);
  assign popcount22_43n0_core_071 = ~input_a[16];
  assign popcount22_43n0_core_073 = ~input_a[1];
  assign popcount22_43n0_core_074_not = ~input_a[16];
  assign popcount22_43n0_core_075 = input_a[15] ^ input_a[7];
  assign popcount22_43n0_core_077 = ~input_a[1];
  assign popcount22_43n0_core_078 = ~(input_a[14] ^ input_a[13]);
  assign popcount22_43n0_core_079 = input_a[4] ^ input_a[14];
  assign popcount22_43n0_core_080 = input_a[20] & input_a[1];
  assign popcount22_43n0_core_081 = ~(input_a[14] & input_a[20]);
  assign popcount22_43n0_core_082 = input_a[11] | input_a[19];
  assign popcount22_43n0_core_085 = ~(input_a[11] ^ input_a[15]);
  assign popcount22_43n0_core_090 = ~(input_a[11] | input_a[13]);
  assign popcount22_43n0_core_092 = input_a[9] | input_a[15];
  assign popcount22_43n0_core_093 = input_a[10] & input_a[0];
  assign popcount22_43n0_core_094 = input_a[8] & input_a[6];
  assign popcount22_43n0_core_096 = ~(input_a[17] | input_a[16]);
  assign popcount22_43n0_core_097 = ~(input_a[14] ^ input_a[5]);
  assign popcount22_43n0_core_098 = ~(input_a[11] & input_a[5]);
  assign popcount22_43n0_core_100 = ~(input_a[10] | input_a[20]);
  assign popcount22_43n0_core_101 = ~input_a[18];
  assign popcount22_43n0_core_102 = ~(input_a[14] | input_a[2]);
  assign popcount22_43n0_core_105 = input_a[3] | input_a[19];
  assign popcount22_43n0_core_107 = input_a[5] & input_a[5];
  assign popcount22_43n0_core_108 = ~(input_a[6] | input_a[2]);
  assign popcount22_43n0_core_109 = ~(input_a[10] & input_a[20]);
  assign popcount22_43n0_core_110 = ~(input_a[4] & input_a[18]);
  assign popcount22_43n0_core_113 = ~(input_a[5] ^ input_a[15]);
  assign popcount22_43n0_core_115 = input_a[3] | input_a[6];
  assign popcount22_43n0_core_116 = input_a[17] | input_a[5];
  assign popcount22_43n0_core_117_not = ~input_a[13];
  assign popcount22_43n0_core_118 = ~(input_a[18] & input_a[6]);
  assign popcount22_43n0_core_119 = input_a[0] ^ input_a[20];
  assign popcount22_43n0_core_124 = ~input_a[20];
  assign popcount22_43n0_core_126 = input_a[14] | input_a[7];
  assign popcount22_43n0_core_130 = input_a[14] & input_a[10];
  assign popcount22_43n0_core_133 = ~input_a[18];
  assign popcount22_43n0_core_134 = input_a[12] ^ input_a[3];
  assign popcount22_43n0_core_135 = input_a[15] & input_a[16];
  assign popcount22_43n0_core_137 = input_a[17] ^ input_a[6];
  assign popcount22_43n0_core_138 = input_a[15] | input_a[4];
  assign popcount22_43n0_core_139 = ~(input_a[17] ^ input_a[4]);
  assign popcount22_43n0_core_140 = ~input_a[16];
  assign popcount22_43n0_core_141 = ~(input_a[10] ^ input_a[6]);
  assign popcount22_43n0_core_143 = ~(input_a[10] & input_a[8]);
  assign popcount22_43n0_core_144 = input_a[14] & input_a[14];
  assign popcount22_43n0_core_146 = ~(input_a[12] & input_a[13]);
  assign popcount22_43n0_core_147 = ~(input_a[20] | input_a[11]);
  assign popcount22_43n0_core_149 = ~input_a[19];
  assign popcount22_43n0_core_152 = input_a[14] ^ input_a[17];
  assign popcount22_43n0_core_153 = ~input_a[12];
  assign popcount22_43n0_core_156 = ~(input_a[17] ^ input_a[6]);
  assign popcount22_43n0_core_157 = ~(input_a[20] | input_a[11]);
  assign popcount22_43n0_core_159 = ~(input_a[18] ^ input_a[21]);
  assign popcount22_43n0_core_160 = ~input_a[2];

  assign popcount22_43n0_out[0] = input_a[8];
  assign popcount22_43n0_out[1] = input_a[1];
  assign popcount22_43n0_out[2] = input_a[1];
  assign popcount22_43n0_out[3] = 1'b1;
  assign popcount22_43n0_out[4] = input_a[5];
endmodule