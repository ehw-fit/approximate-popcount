// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.85007
// WCE=11.0
// EP=0.831812%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_409n(input [21:0] input_a, output [4:0] popcount22_409n_out);
  wire popcount22_409n_core_024;
  wire popcount22_409n_core_026;
  wire popcount22_409n_core_027;
  wire popcount22_409n_core_028;
  wire popcount22_409n_core_029;
  wire popcount22_409n_core_031;
  wire popcount22_409n_core_034;
  wire popcount22_409n_core_036;
  wire popcount22_409n_core_039;
  wire popcount22_409n_core_040;
  wire popcount22_409n_core_041_not;
  wire popcount22_409n_core_042;
  wire popcount22_409n_core_043;
  wire popcount22_409n_core_045;
  wire popcount22_409n_core_046;
  wire popcount22_409n_core_047;
  wire popcount22_409n_core_052;
  wire popcount22_409n_core_053;
  wire popcount22_409n_core_054;
  wire popcount22_409n_core_055;
  wire popcount22_409n_core_056;
  wire popcount22_409n_core_061;
  wire popcount22_409n_core_063;
  wire popcount22_409n_core_064;
  wire popcount22_409n_core_067;
  wire popcount22_409n_core_068_not;
  wire popcount22_409n_core_069_not;
  wire popcount22_409n_core_070;
  wire popcount22_409n_core_071;
  wire popcount22_409n_core_072;
  wire popcount22_409n_core_074;
  wire popcount22_409n_core_076;
  wire popcount22_409n_core_078;
  wire popcount22_409n_core_079;
  wire popcount22_409n_core_081;
  wire popcount22_409n_core_084;
  wire popcount22_409n_core_086;
  wire popcount22_409n_core_087;
  wire popcount22_409n_core_088;
  wire popcount22_409n_core_089;
  wire popcount22_409n_core_093;
  wire popcount22_409n_core_094;
  wire popcount22_409n_core_095;
  wire popcount22_409n_core_097;
  wire popcount22_409n_core_098;
  wire popcount22_409n_core_099;
  wire popcount22_409n_core_100_not;
  wire popcount22_409n_core_101;
  wire popcount22_409n_core_104;
  wire popcount22_409n_core_106;
  wire popcount22_409n_core_111;
  wire popcount22_409n_core_112;
  wire popcount22_409n_core_113;
  wire popcount22_409n_core_114;
  wire popcount22_409n_core_116;
  wire popcount22_409n_core_117;
  wire popcount22_409n_core_118;
  wire popcount22_409n_core_123;
  wire popcount22_409n_core_124;
  wire popcount22_409n_core_125;
  wire popcount22_409n_core_126;
  wire popcount22_409n_core_130;
  wire popcount22_409n_core_132;
  wire popcount22_409n_core_133;
  wire popcount22_409n_core_134;
  wire popcount22_409n_core_135;
  wire popcount22_409n_core_138;
  wire popcount22_409n_core_139;
  wire popcount22_409n_core_140;
  wire popcount22_409n_core_142;
  wire popcount22_409n_core_143;
  wire popcount22_409n_core_146;
  wire popcount22_409n_core_147;
  wire popcount22_409n_core_148;
  wire popcount22_409n_core_149;
  wire popcount22_409n_core_150;
  wire popcount22_409n_core_151;
  wire popcount22_409n_core_152;
  wire popcount22_409n_core_153;
  wire popcount22_409n_core_154;
  wire popcount22_409n_core_158;
  wire popcount22_409n_core_159_not;
  wire popcount22_409n_core_160;
  wire popcount22_409n_core_161;

  assign popcount22_409n_core_024 = input_a[14] ^ input_a[7];
  assign popcount22_409n_core_026 = input_a[13] & input_a[12];
  assign popcount22_409n_core_027 = ~(input_a[1] ^ input_a[4]);
  assign popcount22_409n_core_028 = input_a[0] ^ input_a[21];
  assign popcount22_409n_core_029 = ~(input_a[21] & input_a[14]);
  assign popcount22_409n_core_031 = ~(input_a[2] & input_a[13]);
  assign popcount22_409n_core_034 = input_a[15] ^ input_a[14];
  assign popcount22_409n_core_036 = input_a[1] | input_a[18];
  assign popcount22_409n_core_039 = ~(input_a[13] ^ input_a[11]);
  assign popcount22_409n_core_040 = ~(input_a[2] | input_a[17]);
  assign popcount22_409n_core_041_not = ~input_a[21];
  assign popcount22_409n_core_042 = ~(input_a[12] ^ input_a[17]);
  assign popcount22_409n_core_043 = input_a[7] ^ input_a[14];
  assign popcount22_409n_core_045 = ~(input_a[5] | input_a[4]);
  assign popcount22_409n_core_046 = ~(input_a[8] | input_a[0]);
  assign popcount22_409n_core_047 = ~(input_a[14] ^ input_a[0]);
  assign popcount22_409n_core_052 = input_a[13] | input_a[4];
  assign popcount22_409n_core_053 = ~input_a[12];
  assign popcount22_409n_core_054 = input_a[14] | input_a[6];
  assign popcount22_409n_core_055 = ~(input_a[7] ^ input_a[10]);
  assign popcount22_409n_core_056 = ~(input_a[0] | input_a[8]);
  assign popcount22_409n_core_061 = ~(input_a[13] | input_a[3]);
  assign popcount22_409n_core_063 = ~(input_a[9] | input_a[13]);
  assign popcount22_409n_core_064 = ~(input_a[6] | input_a[21]);
  assign popcount22_409n_core_067 = input_a[16] ^ input_a[0];
  assign popcount22_409n_core_068_not = ~input_a[2];
  assign popcount22_409n_core_069_not = ~input_a[10];
  assign popcount22_409n_core_070 = ~input_a[8];
  assign popcount22_409n_core_071 = input_a[11] ^ input_a[14];
  assign popcount22_409n_core_072 = ~(input_a[13] | input_a[9]);
  assign popcount22_409n_core_074 = ~input_a[0];
  assign popcount22_409n_core_076 = input_a[1] | input_a[6];
  assign popcount22_409n_core_078 = ~(input_a[11] | input_a[21]);
  assign popcount22_409n_core_079 = ~(input_a[19] | input_a[16]);
  assign popcount22_409n_core_081 = ~(input_a[5] & input_a[4]);
  assign popcount22_409n_core_084 = input_a[10] | input_a[21];
  assign popcount22_409n_core_086 = input_a[16] | input_a[18];
  assign popcount22_409n_core_087 = ~(input_a[18] & input_a[14]);
  assign popcount22_409n_core_088 = ~input_a[2];
  assign popcount22_409n_core_089 = ~input_a[20];
  assign popcount22_409n_core_093 = input_a[1] | input_a[17];
  assign popcount22_409n_core_094 = ~(input_a[20] | input_a[10]);
  assign popcount22_409n_core_095 = ~(input_a[13] ^ input_a[13]);
  assign popcount22_409n_core_097 = ~(input_a[4] | input_a[12]);
  assign popcount22_409n_core_098 = ~(input_a[13] & input_a[0]);
  assign popcount22_409n_core_099 = ~(input_a[21] | input_a[7]);
  assign popcount22_409n_core_100_not = ~input_a[13];
  assign popcount22_409n_core_101 = ~(input_a[14] | input_a[6]);
  assign popcount22_409n_core_104 = ~(input_a[16] & input_a[0]);
  assign popcount22_409n_core_106 = input_a[21] | input_a[2];
  assign popcount22_409n_core_111 = ~input_a[9];
  assign popcount22_409n_core_112 = ~input_a[6];
  assign popcount22_409n_core_113 = ~(input_a[14] & input_a[1]);
  assign popcount22_409n_core_114 = input_a[5] & input_a[16];
  assign popcount22_409n_core_116 = ~(input_a[13] ^ input_a[12]);
  assign popcount22_409n_core_117 = ~(input_a[13] ^ input_a[21]);
  assign popcount22_409n_core_118 = ~input_a[7];
  assign popcount22_409n_core_123 = input_a[11] ^ input_a[15];
  assign popcount22_409n_core_124 = ~(input_a[1] & input_a[18]);
  assign popcount22_409n_core_125 = ~(input_a[6] & input_a[16]);
  assign popcount22_409n_core_126 = ~input_a[8];
  assign popcount22_409n_core_130 = input_a[20] & input_a[8];
  assign popcount22_409n_core_132 = input_a[13] & input_a[18];
  assign popcount22_409n_core_133 = ~input_a[16];
  assign popcount22_409n_core_134 = input_a[10] & input_a[12];
  assign popcount22_409n_core_135 = input_a[0] ^ input_a[18];
  assign popcount22_409n_core_138 = ~input_a[6];
  assign popcount22_409n_core_139 = ~input_a[13];
  assign popcount22_409n_core_140 = input_a[10] & input_a[12];
  assign popcount22_409n_core_142 = ~(input_a[9] & input_a[15]);
  assign popcount22_409n_core_143 = input_a[14] | input_a[7];
  assign popcount22_409n_core_146 = ~(input_a[16] & input_a[5]);
  assign popcount22_409n_core_147 = ~input_a[17];
  assign popcount22_409n_core_148 = input_a[6] ^ input_a[21];
  assign popcount22_409n_core_149 = input_a[0] & input_a[16];
  assign popcount22_409n_core_150 = ~(input_a[15] & input_a[0]);
  assign popcount22_409n_core_151 = ~(input_a[17] ^ input_a[8]);
  assign popcount22_409n_core_152 = ~input_a[17];
  assign popcount22_409n_core_153 = ~(input_a[17] | input_a[9]);
  assign popcount22_409n_core_154 = input_a[19] & input_a[1];
  assign popcount22_409n_core_158 = input_a[8] & input_a[18];
  assign popcount22_409n_core_159_not = ~input_a[6];
  assign popcount22_409n_core_160 = ~(input_a[19] & input_a[11]);
  assign popcount22_409n_core_161 = ~input_a[14];

  assign popcount22_409n_out[0] = 1'b1;
  assign popcount22_409n_out[1] = 1'b1;
  assign popcount22_409n_out[2] = 1'b0;
  assign popcount22_409n_out[3] = 1'b1;
  assign popcount22_409n_out[4] = 1'b0;
endmodule