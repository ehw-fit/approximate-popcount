// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.69209
// WCE=27.0
// EP=0.943799%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_un7b(input [35:0] input_a, output [5:0] popcount36_un7b_out);
  wire popcount36_un7b_core_038;
  wire popcount36_un7b_core_039;
  wire popcount36_un7b_core_040;
  wire popcount36_un7b_core_042;
  wire popcount36_un7b_core_043;
  wire popcount36_un7b_core_044;
  wire popcount36_un7b_core_045;
  wire popcount36_un7b_core_047;
  wire popcount36_un7b_core_049;
  wire popcount36_un7b_core_050;
  wire popcount36_un7b_core_051;
  wire popcount36_un7b_core_052;
  wire popcount36_un7b_core_054;
  wire popcount36_un7b_core_055;
  wire popcount36_un7b_core_056;
  wire popcount36_un7b_core_058;
  wire popcount36_un7b_core_059;
  wire popcount36_un7b_core_060;
  wire popcount36_un7b_core_062;
  wire popcount36_un7b_core_063;
  wire popcount36_un7b_core_064;
  wire popcount36_un7b_core_065;
  wire popcount36_un7b_core_068;
  wire popcount36_un7b_core_069;
  wire popcount36_un7b_core_070;
  wire popcount36_un7b_core_071;
  wire popcount36_un7b_core_072;
  wire popcount36_un7b_core_074;
  wire popcount36_un7b_core_075;
  wire popcount36_un7b_core_076;
  wire popcount36_un7b_core_077;
  wire popcount36_un7b_core_081;
  wire popcount36_un7b_core_083;
  wire popcount36_un7b_core_084;
  wire popcount36_un7b_core_087;
  wire popcount36_un7b_core_089;
  wire popcount36_un7b_core_090;
  wire popcount36_un7b_core_092;
  wire popcount36_un7b_core_093;
  wire popcount36_un7b_core_094;
  wire popcount36_un7b_core_095;
  wire popcount36_un7b_core_097;
  wire popcount36_un7b_core_100;
  wire popcount36_un7b_core_103;
  wire popcount36_un7b_core_104_not;
  wire popcount36_un7b_core_107;
  wire popcount36_un7b_core_108;
  wire popcount36_un7b_core_110;
  wire popcount36_un7b_core_111;
  wire popcount36_un7b_core_118;
  wire popcount36_un7b_core_119;
  wire popcount36_un7b_core_121;
  wire popcount36_un7b_core_124;
  wire popcount36_un7b_core_126;
  wire popcount36_un7b_core_127;
  wire popcount36_un7b_core_128;
  wire popcount36_un7b_core_130;
  wire popcount36_un7b_core_131;
  wire popcount36_un7b_core_133;
  wire popcount36_un7b_core_134;
  wire popcount36_un7b_core_135;
  wire popcount36_un7b_core_136;
  wire popcount36_un7b_core_137;
  wire popcount36_un7b_core_138_not;
  wire popcount36_un7b_core_139;
  wire popcount36_un7b_core_144;
  wire popcount36_un7b_core_145;
  wire popcount36_un7b_core_146;
  wire popcount36_un7b_core_149;
  wire popcount36_un7b_core_150;
  wire popcount36_un7b_core_151;
  wire popcount36_un7b_core_153;
  wire popcount36_un7b_core_154;
  wire popcount36_un7b_core_155;
  wire popcount36_un7b_core_157;
  wire popcount36_un7b_core_158;
  wire popcount36_un7b_core_159;
  wire popcount36_un7b_core_160;
  wire popcount36_un7b_core_162;
  wire popcount36_un7b_core_163;
  wire popcount36_un7b_core_166;
  wire popcount36_un7b_core_169;
  wire popcount36_un7b_core_170;
  wire popcount36_un7b_core_172;
  wire popcount36_un7b_core_173;
  wire popcount36_un7b_core_174;
  wire popcount36_un7b_core_177;
  wire popcount36_un7b_core_178;
  wire popcount36_un7b_core_179;
  wire popcount36_un7b_core_181;
  wire popcount36_un7b_core_183;
  wire popcount36_un7b_core_184;
  wire popcount36_un7b_core_186;
  wire popcount36_un7b_core_187;
  wire popcount36_un7b_core_189;
  wire popcount36_un7b_core_191;
  wire popcount36_un7b_core_196;
  wire popcount36_un7b_core_198;
  wire popcount36_un7b_core_199;
  wire popcount36_un7b_core_200;
  wire popcount36_un7b_core_201;
  wire popcount36_un7b_core_202;
  wire popcount36_un7b_core_204;
  wire popcount36_un7b_core_206;
  wire popcount36_un7b_core_207;
  wire popcount36_un7b_core_208;
  wire popcount36_un7b_core_209;
  wire popcount36_un7b_core_210;
  wire popcount36_un7b_core_211;
  wire popcount36_un7b_core_213;
  wire popcount36_un7b_core_215;
  wire popcount36_un7b_core_216;
  wire popcount36_un7b_core_217;
  wire popcount36_un7b_core_218;
  wire popcount36_un7b_core_219;
  wire popcount36_un7b_core_220;
  wire popcount36_un7b_core_221;
  wire popcount36_un7b_core_222;
  wire popcount36_un7b_core_225;
  wire popcount36_un7b_core_228;
  wire popcount36_un7b_core_229;
  wire popcount36_un7b_core_230;
  wire popcount36_un7b_core_232;
  wire popcount36_un7b_core_233;
  wire popcount36_un7b_core_234;
  wire popcount36_un7b_core_235;
  wire popcount36_un7b_core_238;
  wire popcount36_un7b_core_239;
  wire popcount36_un7b_core_240;
  wire popcount36_un7b_core_244;
  wire popcount36_un7b_core_245;
  wire popcount36_un7b_core_246;
  wire popcount36_un7b_core_248;
  wire popcount36_un7b_core_249;
  wire popcount36_un7b_core_250;
  wire popcount36_un7b_core_251;
  wire popcount36_un7b_core_253;
  wire popcount36_un7b_core_254;
  wire popcount36_un7b_core_255;
  wire popcount36_un7b_core_257;
  wire popcount36_un7b_core_258;
  wire popcount36_un7b_core_259;
  wire popcount36_un7b_core_260;
  wire popcount36_un7b_core_261;
  wire popcount36_un7b_core_262;
  wire popcount36_un7b_core_263;
  wire popcount36_un7b_core_265;
  wire popcount36_un7b_core_267;
  wire popcount36_un7b_core_269;
  wire popcount36_un7b_core_270;
  wire popcount36_un7b_core_272;
  wire popcount36_un7b_core_274;
  wire popcount36_un7b_core_275;
  wire popcount36_un7b_core_276;

  assign popcount36_un7b_core_038 = input_a[33] ^ input_a[10];
  assign popcount36_un7b_core_039 = ~(input_a[16] ^ input_a[29]);
  assign popcount36_un7b_core_040 = ~(input_a[12] & input_a[2]);
  assign popcount36_un7b_core_042 = ~(input_a[3] ^ input_a[34]);
  assign popcount36_un7b_core_043 = ~(input_a[20] & input_a[7]);
  assign popcount36_un7b_core_044 = input_a[22] & input_a[34];
  assign popcount36_un7b_core_045 = ~(input_a[19] ^ input_a[5]);
  assign popcount36_un7b_core_047 = ~input_a[10];
  assign popcount36_un7b_core_049 = ~input_a[25];
  assign popcount36_un7b_core_050 = ~input_a[32];
  assign popcount36_un7b_core_051 = input_a[1] & input_a[8];
  assign popcount36_un7b_core_052 = input_a[19] | input_a[13];
  assign popcount36_un7b_core_054 = input_a[0] & input_a[11];
  assign popcount36_un7b_core_055 = ~input_a[5];
  assign popcount36_un7b_core_056 = ~(input_a[22] | input_a[27]);
  assign popcount36_un7b_core_058 = input_a[15] & input_a[31];
  assign popcount36_un7b_core_059 = ~(input_a[25] ^ input_a[1]);
  assign popcount36_un7b_core_060 = ~(input_a[32] | input_a[29]);
  assign popcount36_un7b_core_062 = input_a[1] & input_a[7];
  assign popcount36_un7b_core_063 = input_a[18] ^ input_a[13];
  assign popcount36_un7b_core_064 = ~(input_a[17] ^ input_a[30]);
  assign popcount36_un7b_core_065 = ~(input_a[15] | input_a[20]);
  assign popcount36_un7b_core_068 = ~(input_a[29] & input_a[23]);
  assign popcount36_un7b_core_069 = ~(input_a[22] & input_a[25]);
  assign popcount36_un7b_core_070 = ~(input_a[21] & input_a[12]);
  assign popcount36_un7b_core_071 = ~(input_a[23] | input_a[6]);
  assign popcount36_un7b_core_072 = ~(input_a[18] & input_a[4]);
  assign popcount36_un7b_core_074 = input_a[31] & input_a[1];
  assign popcount36_un7b_core_075 = ~input_a[25];
  assign popcount36_un7b_core_076 = input_a[12] & input_a[19];
  assign popcount36_un7b_core_077 = ~(input_a[25] ^ input_a[1]);
  assign popcount36_un7b_core_081 = ~(input_a[27] ^ input_a[6]);
  assign popcount36_un7b_core_083 = ~(input_a[16] | input_a[10]);
  assign popcount36_un7b_core_084 = ~input_a[13];
  assign popcount36_un7b_core_087 = input_a[19] | input_a[9];
  assign popcount36_un7b_core_089 = input_a[21] | input_a[27];
  assign popcount36_un7b_core_090 = ~(input_a[9] ^ input_a[3]);
  assign popcount36_un7b_core_092 = input_a[25] ^ input_a[1];
  assign popcount36_un7b_core_093 = input_a[33] ^ input_a[33];
  assign popcount36_un7b_core_094 = ~(input_a[3] | input_a[10]);
  assign popcount36_un7b_core_095 = input_a[12] & input_a[19];
  assign popcount36_un7b_core_097 = ~(input_a[17] ^ input_a[28]);
  assign popcount36_un7b_core_100 = input_a[1] & input_a[3];
  assign popcount36_un7b_core_103 = ~input_a[19];
  assign popcount36_un7b_core_104_not = ~input_a[21];
  assign popcount36_un7b_core_107 = ~(input_a[23] | input_a[29]);
  assign popcount36_un7b_core_108 = input_a[20] & input_a[5];
  assign popcount36_un7b_core_110 = ~input_a[27];
  assign popcount36_un7b_core_111 = ~(input_a[19] & input_a[6]);
  assign popcount36_un7b_core_118 = input_a[8] & input_a[24];
  assign popcount36_un7b_core_119 = input_a[21] & input_a[19];
  assign popcount36_un7b_core_121 = ~(input_a[31] & input_a[12]);
  assign popcount36_un7b_core_124 = input_a[5] | input_a[22];
  assign popcount36_un7b_core_126 = input_a[31] ^ input_a[16];
  assign popcount36_un7b_core_127 = ~(input_a[35] ^ input_a[4]);
  assign popcount36_un7b_core_128 = input_a[17] ^ input_a[28];
  assign popcount36_un7b_core_130 = input_a[33] ^ input_a[20];
  assign popcount36_un7b_core_131 = input_a[31] | input_a[21];
  assign popcount36_un7b_core_133 = ~(input_a[13] ^ input_a[14]);
  assign popcount36_un7b_core_134 = input_a[8] | input_a[31];
  assign popcount36_un7b_core_135 = input_a[24] | input_a[16];
  assign popcount36_un7b_core_136 = ~(input_a[8] | input_a[0]);
  assign popcount36_un7b_core_137 = ~(input_a[5] ^ input_a[8]);
  assign popcount36_un7b_core_138_not = ~input_a[22];
  assign popcount36_un7b_core_139 = input_a[15] ^ input_a[18];
  assign popcount36_un7b_core_144 = input_a[34] | input_a[4];
  assign popcount36_un7b_core_145 = ~(input_a[26] ^ input_a[23]);
  assign popcount36_un7b_core_146 = input_a[4] & input_a[16];
  assign popcount36_un7b_core_149 = input_a[28] ^ input_a[1];
  assign popcount36_un7b_core_150 = ~(input_a[34] ^ input_a[26]);
  assign popcount36_un7b_core_151 = ~(input_a[5] & input_a[0]);
  assign popcount36_un7b_core_153 = input_a[26] ^ input_a[13];
  assign popcount36_un7b_core_154 = ~(input_a[25] ^ input_a[24]);
  assign popcount36_un7b_core_155 = input_a[29] ^ input_a[19];
  assign popcount36_un7b_core_157 = ~input_a[13];
  assign popcount36_un7b_core_158 = ~(input_a[24] & input_a[3]);
  assign popcount36_un7b_core_159 = ~(input_a[5] | input_a[31]);
  assign popcount36_un7b_core_160 = input_a[28] ^ input_a[4];
  assign popcount36_un7b_core_162 = ~input_a[32];
  assign popcount36_un7b_core_163 = input_a[22] ^ input_a[33];
  assign popcount36_un7b_core_166 = ~input_a[27];
  assign popcount36_un7b_core_169 = ~(input_a[22] & input_a[5]);
  assign popcount36_un7b_core_170 = input_a[19] ^ input_a[34];
  assign popcount36_un7b_core_172 = input_a[2] ^ input_a[32];
  assign popcount36_un7b_core_173 = ~(input_a[25] ^ input_a[21]);
  assign popcount36_un7b_core_174 = ~input_a[1];
  assign popcount36_un7b_core_177 = ~input_a[13];
  assign popcount36_un7b_core_178 = ~(input_a[30] & input_a[29]);
  assign popcount36_un7b_core_179 = ~(input_a[8] & input_a[20]);
  assign popcount36_un7b_core_181 = ~(input_a[14] & input_a[19]);
  assign popcount36_un7b_core_183 = ~(input_a[29] ^ input_a[22]);
  assign popcount36_un7b_core_184 = input_a[30] | input_a[33];
  assign popcount36_un7b_core_186 = input_a[34] ^ input_a[16];
  assign popcount36_un7b_core_187 = ~(input_a[3] | input_a[2]);
  assign popcount36_un7b_core_189 = ~(input_a[9] | input_a[0]);
  assign popcount36_un7b_core_191 = input_a[20] & input_a[29];
  assign popcount36_un7b_core_196 = ~(input_a[8] & input_a[24]);
  assign popcount36_un7b_core_198 = ~(input_a[20] & input_a[0]);
  assign popcount36_un7b_core_199 = input_a[27] ^ input_a[25];
  assign popcount36_un7b_core_200 = ~(input_a[26] ^ input_a[22]);
  assign popcount36_un7b_core_201 = input_a[34] & input_a[27];
  assign popcount36_un7b_core_202 = ~input_a[34];
  assign popcount36_un7b_core_204 = ~input_a[3];
  assign popcount36_un7b_core_206 = input_a[23] & input_a[18];
  assign popcount36_un7b_core_207 = ~input_a[15];
  assign popcount36_un7b_core_208 = ~(input_a[13] | input_a[29]);
  assign popcount36_un7b_core_209 = ~input_a[11];
  assign popcount36_un7b_core_210 = input_a[13] & input_a[0];
  assign popcount36_un7b_core_211 = input_a[6] & input_a[22];
  assign popcount36_un7b_core_213 = input_a[30] & input_a[24];
  assign popcount36_un7b_core_215 = ~input_a[14];
  assign popcount36_un7b_core_216 = input_a[9] | input_a[13];
  assign popcount36_un7b_core_217 = input_a[22] ^ input_a[6];
  assign popcount36_un7b_core_218 = ~(input_a[26] & input_a[17]);
  assign popcount36_un7b_core_219 = ~(input_a[35] & input_a[11]);
  assign popcount36_un7b_core_220 = ~input_a[15];
  assign popcount36_un7b_core_221 = input_a[28] | input_a[2];
  assign popcount36_un7b_core_222 = input_a[19] | input_a[22];
  assign popcount36_un7b_core_225 = ~(input_a[17] & input_a[18]);
  assign popcount36_un7b_core_228 = input_a[13] | input_a[1];
  assign popcount36_un7b_core_229 = ~(input_a[33] ^ input_a[8]);
  assign popcount36_un7b_core_230 = input_a[23] ^ input_a[11];
  assign popcount36_un7b_core_232 = ~(input_a[1] | input_a[17]);
  assign popcount36_un7b_core_233 = input_a[30] ^ input_a[23];
  assign popcount36_un7b_core_234 = ~(input_a[15] | input_a[5]);
  assign popcount36_un7b_core_235 = ~(input_a[2] & input_a[16]);
  assign popcount36_un7b_core_238 = ~(input_a[26] | input_a[17]);
  assign popcount36_un7b_core_239 = input_a[14] ^ input_a[34];
  assign popcount36_un7b_core_240 = ~input_a[24];
  assign popcount36_un7b_core_244 = ~(input_a[29] ^ input_a[10]);
  assign popcount36_un7b_core_245 = ~(input_a[23] ^ input_a[8]);
  assign popcount36_un7b_core_246 = input_a[30] & input_a[28];
  assign popcount36_un7b_core_248 = ~input_a[23];
  assign popcount36_un7b_core_249 = ~input_a[4];
  assign popcount36_un7b_core_250 = ~input_a[11];
  assign popcount36_un7b_core_251 = input_a[5] & input_a[35];
  assign popcount36_un7b_core_253 = ~input_a[33];
  assign popcount36_un7b_core_254 = input_a[8] ^ input_a[30];
  assign popcount36_un7b_core_255 = input_a[28] & input_a[14];
  assign popcount36_un7b_core_257 = ~input_a[0];
  assign popcount36_un7b_core_258 = ~input_a[34];
  assign popcount36_un7b_core_259 = ~(input_a[35] | input_a[28]);
  assign popcount36_un7b_core_260 = ~(input_a[25] ^ input_a[20]);
  assign popcount36_un7b_core_261 = ~(input_a[10] ^ input_a[17]);
  assign popcount36_un7b_core_262 = ~(input_a[19] ^ input_a[5]);
  assign popcount36_un7b_core_263 = ~(input_a[6] ^ input_a[16]);
  assign popcount36_un7b_core_265 = ~(input_a[9] & input_a[20]);
  assign popcount36_un7b_core_267 = ~input_a[21];
  assign popcount36_un7b_core_269 = ~input_a[9];
  assign popcount36_un7b_core_270 = input_a[13] & input_a[3];
  assign popcount36_un7b_core_272 = ~input_a[11];
  assign popcount36_un7b_core_274 = ~(input_a[16] | input_a[13]);
  assign popcount36_un7b_core_275 = input_a[13] | input_a[28];
  assign popcount36_un7b_core_276 = ~(input_a[19] & input_a[3]);

  assign popcount36_un7b_out[0] = 1'b0;
  assign popcount36_un7b_out[1] = input_a[0];
  assign popcount36_un7b_out[2] = input_a[21];
  assign popcount36_un7b_out[3] = input_a[19];
  assign popcount36_un7b_out[4] = 1'b1;
  assign popcount36_un7b_out[5] = 1'b0;
endmodule