// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=9.91731
// WCE=28.0
// EP=0.953631%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_39ti(input [20:0] input_a, output [4:0] popcount21_39ti_out);
  wire popcount21_39ti_core_023;
  wire popcount21_39ti_core_025;
  wire popcount21_39ti_core_031;
  wire popcount21_39ti_core_032;
  wire popcount21_39ti_core_033;
  wire popcount21_39ti_core_034;
  wire popcount21_39ti_core_036;
  wire popcount21_39ti_core_037_not;
  wire popcount21_39ti_core_038;
  wire popcount21_39ti_core_040;
  wire popcount21_39ti_core_043;
  wire popcount21_39ti_core_045;
  wire popcount21_39ti_core_048;
  wire popcount21_39ti_core_049;
  wire popcount21_39ti_core_051;
  wire popcount21_39ti_core_052;
  wire popcount21_39ti_core_055_not;
  wire popcount21_39ti_core_056;
  wire popcount21_39ti_core_057;
  wire popcount21_39ti_core_059;
  wire popcount21_39ti_core_063;
  wire popcount21_39ti_core_066;
  wire popcount21_39ti_core_067;
  wire popcount21_39ti_core_068_not;
  wire popcount21_39ti_core_069;
  wire popcount21_39ti_core_072;
  wire popcount21_39ti_core_075_not;
  wire popcount21_39ti_core_077;
  wire popcount21_39ti_core_079;
  wire popcount21_39ti_core_080;
  wire popcount21_39ti_core_081;
  wire popcount21_39ti_core_083;
  wire popcount21_39ti_core_085;
  wire popcount21_39ti_core_087;
  wire popcount21_39ti_core_088;
  wire popcount21_39ti_core_093;
  wire popcount21_39ti_core_094;
  wire popcount21_39ti_core_095;
  wire popcount21_39ti_core_096;
  wire popcount21_39ti_core_098;
  wire popcount21_39ti_core_100;
  wire popcount21_39ti_core_103;
  wire popcount21_39ti_core_106;
  wire popcount21_39ti_core_107;
  wire popcount21_39ti_core_108;
  wire popcount21_39ti_core_109;
  wire popcount21_39ti_core_110;
  wire popcount21_39ti_core_114;
  wire popcount21_39ti_core_116;
  wire popcount21_39ti_core_117;
  wire popcount21_39ti_core_120;
  wire popcount21_39ti_core_121;
  wire popcount21_39ti_core_123;
  wire popcount21_39ti_core_124;
  wire popcount21_39ti_core_125;
  wire popcount21_39ti_core_126_not;
  wire popcount21_39ti_core_127;
  wire popcount21_39ti_core_128;
  wire popcount21_39ti_core_129;
  wire popcount21_39ti_core_130;
  wire popcount21_39ti_core_131;
  wire popcount21_39ti_core_132;
  wire popcount21_39ti_core_133;
  wire popcount21_39ti_core_135;
  wire popcount21_39ti_core_136;
  wire popcount21_39ti_core_137;
  wire popcount21_39ti_core_138;
  wire popcount21_39ti_core_139;
  wire popcount21_39ti_core_140;
  wire popcount21_39ti_core_142;
  wire popcount21_39ti_core_143;
  wire popcount21_39ti_core_145_not;
  wire popcount21_39ti_core_149;
  wire popcount21_39ti_core_151;
  wire popcount21_39ti_core_152;
  wire popcount21_39ti_core_153;

  assign popcount21_39ti_core_023 = input_a[8] | input_a[12];
  assign popcount21_39ti_core_025 = ~(input_a[0] & input_a[6]);
  assign popcount21_39ti_core_031 = ~input_a[15];
  assign popcount21_39ti_core_032 = ~(input_a[5] | input_a[14]);
  assign popcount21_39ti_core_033 = ~(input_a[6] | input_a[20]);
  assign popcount21_39ti_core_034 = input_a[13] ^ input_a[2];
  assign popcount21_39ti_core_036 = ~(input_a[20] & input_a[7]);
  assign popcount21_39ti_core_037_not = ~input_a[2];
  assign popcount21_39ti_core_038 = input_a[5] | input_a[12];
  assign popcount21_39ti_core_040 = ~(input_a[5] ^ input_a[10]);
  assign popcount21_39ti_core_043 = input_a[12] | input_a[2];
  assign popcount21_39ti_core_045 = input_a[15] | input_a[5];
  assign popcount21_39ti_core_048 = input_a[11] | input_a[10];
  assign popcount21_39ti_core_049 = ~(input_a[11] & input_a[19]);
  assign popcount21_39ti_core_051 = ~(input_a[9] | input_a[0]);
  assign popcount21_39ti_core_052 = ~(input_a[4] & input_a[3]);
  assign popcount21_39ti_core_055_not = ~input_a[1];
  assign popcount21_39ti_core_056 = ~input_a[11];
  assign popcount21_39ti_core_057 = ~(input_a[10] & input_a[5]);
  assign popcount21_39ti_core_059 = input_a[14] & input_a[16];
  assign popcount21_39ti_core_063 = ~(input_a[5] & input_a[20]);
  assign popcount21_39ti_core_066 = input_a[5] ^ input_a[9];
  assign popcount21_39ti_core_067 = ~(input_a[6] ^ input_a[13]);
  assign popcount21_39ti_core_068_not = ~input_a[17];
  assign popcount21_39ti_core_069 = ~input_a[12];
  assign popcount21_39ti_core_072 = ~(input_a[7] | input_a[1]);
  assign popcount21_39ti_core_075_not = ~input_a[2];
  assign popcount21_39ti_core_077 = ~input_a[11];
  assign popcount21_39ti_core_079 = ~(input_a[14] & input_a[11]);
  assign popcount21_39ti_core_080 = ~input_a[19];
  assign popcount21_39ti_core_081 = ~(input_a[15] | input_a[10]);
  assign popcount21_39ti_core_083 = ~(input_a[20] & input_a[11]);
  assign popcount21_39ti_core_085 = input_a[4] ^ input_a[13];
  assign popcount21_39ti_core_087 = input_a[13] | input_a[9];
  assign popcount21_39ti_core_088 = input_a[4] ^ input_a[6];
  assign popcount21_39ti_core_093 = input_a[18] ^ input_a[15];
  assign popcount21_39ti_core_094 = ~(input_a[10] & input_a[0]);
  assign popcount21_39ti_core_095 = input_a[13] | input_a[10];
  assign popcount21_39ti_core_096 = input_a[18] | input_a[9];
  assign popcount21_39ti_core_098 = input_a[9] | input_a[8];
  assign popcount21_39ti_core_100 = input_a[1] & input_a[17];
  assign popcount21_39ti_core_103 = input_a[9] | input_a[2];
  assign popcount21_39ti_core_106 = ~input_a[7];
  assign popcount21_39ti_core_107 = ~(input_a[20] ^ input_a[3]);
  assign popcount21_39ti_core_108 = ~input_a[15];
  assign popcount21_39ti_core_109 = ~(input_a[9] & input_a[15]);
  assign popcount21_39ti_core_110 = ~(input_a[9] ^ input_a[18]);
  assign popcount21_39ti_core_114 = ~input_a[2];
  assign popcount21_39ti_core_116 = ~(input_a[4] ^ input_a[19]);
  assign popcount21_39ti_core_117 = ~input_a[19];
  assign popcount21_39ti_core_120 = ~input_a[5];
  assign popcount21_39ti_core_121 = input_a[7] & input_a[11];
  assign popcount21_39ti_core_123 = ~input_a[0];
  assign popcount21_39ti_core_124 = input_a[17] & input_a[15];
  assign popcount21_39ti_core_125 = ~(input_a[0] | input_a[9]);
  assign popcount21_39ti_core_126_not = ~input_a[16];
  assign popcount21_39ti_core_127 = ~(input_a[11] & input_a[8]);
  assign popcount21_39ti_core_128 = ~(input_a[4] ^ input_a[15]);
  assign popcount21_39ti_core_129 = ~(input_a[1] & input_a[2]);
  assign popcount21_39ti_core_130 = ~(input_a[8] & input_a[20]);
  assign popcount21_39ti_core_131 = ~(input_a[6] ^ input_a[20]);
  assign popcount21_39ti_core_132 = input_a[0] ^ input_a[4];
  assign popcount21_39ti_core_133 = input_a[6] ^ input_a[4];
  assign popcount21_39ti_core_135 = input_a[8] & input_a[19];
  assign popcount21_39ti_core_136 = input_a[11] | input_a[5];
  assign popcount21_39ti_core_137 = ~(input_a[13] & input_a[11]);
  assign popcount21_39ti_core_138 = input_a[10] ^ input_a[13];
  assign popcount21_39ti_core_139 = ~(input_a[20] & input_a[1]);
  assign popcount21_39ti_core_140 = ~(input_a[9] | input_a[13]);
  assign popcount21_39ti_core_142 = input_a[12] & input_a[12];
  assign popcount21_39ti_core_143 = input_a[13] ^ input_a[3];
  assign popcount21_39ti_core_145_not = ~input_a[0];
  assign popcount21_39ti_core_149 = input_a[13] ^ input_a[5];
  assign popcount21_39ti_core_151 = input_a[14] | input_a[10];
  assign popcount21_39ti_core_152 = ~(input_a[14] & input_a[0]);
  assign popcount21_39ti_core_153 = ~input_a[1];

  assign popcount21_39ti_out[0] = input_a[10];
  assign popcount21_39ti_out[1] = input_a[9];
  assign popcount21_39ti_out[2] = input_a[19];
  assign popcount21_39ti_out[3] = input_a[9];
  assign popcount21_39ti_out[4] = input_a[19];
endmodule