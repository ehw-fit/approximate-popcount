// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.74951
// WCE=15.0
// EP=0.821869%
// Printed PDK parameters:
//  Area=40012537.0
//  Delay=68833048.0
//  Power=1861800.0

module popcount35_3d5j(input [34:0] input_a, output [5:0] popcount35_3d5j_out);
  wire popcount35_3d5j_core_037;
  wire popcount35_3d5j_core_038;
  wire popcount35_3d5j_core_039;
  wire popcount35_3d5j_core_040;
  wire popcount35_3d5j_core_041;
  wire popcount35_3d5j_core_042;
  wire popcount35_3d5j_core_043;
  wire popcount35_3d5j_core_044;
  wire popcount35_3d5j_core_045;
  wire popcount35_3d5j_core_048;
  wire popcount35_3d5j_core_049;
  wire popcount35_3d5j_core_050;
  wire popcount35_3d5j_core_051;
  wire popcount35_3d5j_core_052;
  wire popcount35_3d5j_core_054;
  wire popcount35_3d5j_core_055;
  wire popcount35_3d5j_core_056;
  wire popcount35_3d5j_core_057;
  wire popcount35_3d5j_core_060;
  wire popcount35_3d5j_core_061;
  wire popcount35_3d5j_core_062;
  wire popcount35_3d5j_core_063;
  wire popcount35_3d5j_core_064;
  wire popcount35_3d5j_core_065;
  wire popcount35_3d5j_core_066;
  wire popcount35_3d5j_core_067;
  wire popcount35_3d5j_core_068;
  wire popcount35_3d5j_core_070;
  wire popcount35_3d5j_core_072;
  wire popcount35_3d5j_core_073;
  wire popcount35_3d5j_core_074;
  wire popcount35_3d5j_core_076;
  wire popcount35_3d5j_core_077;
  wire popcount35_3d5j_core_078;
  wire popcount35_3d5j_core_079;
  wire popcount35_3d5j_core_082;
  wire popcount35_3d5j_core_083;
  wire popcount35_3d5j_core_084;
  wire popcount35_3d5j_core_085;
  wire popcount35_3d5j_core_086;
  wire popcount35_3d5j_core_087;
  wire popcount35_3d5j_core_088;
  wire popcount35_3d5j_core_091;
  wire popcount35_3d5j_core_092;
  wire popcount35_3d5j_core_093;
  wire popcount35_3d5j_core_094;
  wire popcount35_3d5j_core_095;
  wire popcount35_3d5j_core_096;
  wire popcount35_3d5j_core_101;
  wire popcount35_3d5j_core_102;
  wire popcount35_3d5j_core_104;
  wire popcount35_3d5j_core_108;
  wire popcount35_3d5j_core_109;
  wire popcount35_3d5j_core_111;
  wire popcount35_3d5j_core_114;
  wire popcount35_3d5j_core_115;
  wire popcount35_3d5j_core_116;
  wire popcount35_3d5j_core_117;
  wire popcount35_3d5j_core_118;
  wire popcount35_3d5j_core_119;
  wire popcount35_3d5j_core_120;
  wire popcount35_3d5j_core_121;
  wire popcount35_3d5j_core_122;
  wire popcount35_3d5j_core_123;
  wire popcount35_3d5j_core_124;
  wire popcount35_3d5j_core_128;
  wire popcount35_3d5j_core_129;
  wire popcount35_3d5j_core_130;
  wire popcount35_3d5j_core_131;
  wire popcount35_3d5j_core_132;
  wire popcount35_3d5j_core_134;
  wire popcount35_3d5j_core_137;
  wire popcount35_3d5j_core_139;
  wire popcount35_3d5j_core_140;
  wire popcount35_3d5j_core_142;
  wire popcount35_3d5j_core_143;
  wire popcount35_3d5j_core_144;
  wire popcount35_3d5j_core_146;
  wire popcount35_3d5j_core_148;
  wire popcount35_3d5j_core_149;
  wire popcount35_3d5j_core_150;
  wire popcount35_3d5j_core_151;
  wire popcount35_3d5j_core_152;
  wire popcount35_3d5j_core_155;
  wire popcount35_3d5j_core_156;
  wire popcount35_3d5j_core_157;
  wire popcount35_3d5j_core_158;
  wire popcount35_3d5j_core_159;
  wire popcount35_3d5j_core_162;
  wire popcount35_3d5j_core_163;
  wire popcount35_3d5j_core_164;
  wire popcount35_3d5j_core_166;
  wire popcount35_3d5j_core_170;
  wire popcount35_3d5j_core_171;
  wire popcount35_3d5j_core_173;
  wire popcount35_3d5j_core_174;
  wire popcount35_3d5j_core_175;
  wire popcount35_3d5j_core_176;
  wire popcount35_3d5j_core_177_not;
  wire popcount35_3d5j_core_178;
  wire popcount35_3d5j_core_179;
  wire popcount35_3d5j_core_180;
  wire popcount35_3d5j_core_182;
  wire popcount35_3d5j_core_184;
  wire popcount35_3d5j_core_185;
  wire popcount35_3d5j_core_188;
  wire popcount35_3d5j_core_190;
  wire popcount35_3d5j_core_192;
  wire popcount35_3d5j_core_193;
  wire popcount35_3d5j_core_194;
  wire popcount35_3d5j_core_195;
  wire popcount35_3d5j_core_197;
  wire popcount35_3d5j_core_198;
  wire popcount35_3d5j_core_200;
  wire popcount35_3d5j_core_201;
  wire popcount35_3d5j_core_203;
  wire popcount35_3d5j_core_204;
  wire popcount35_3d5j_core_205;
  wire popcount35_3d5j_core_206;
  wire popcount35_3d5j_core_207;
  wire popcount35_3d5j_core_209;
  wire popcount35_3d5j_core_211;
  wire popcount35_3d5j_core_212;
  wire popcount35_3d5j_core_213;
  wire popcount35_3d5j_core_214;
  wire popcount35_3d5j_core_215;
  wire popcount35_3d5j_core_217;
  wire popcount35_3d5j_core_218;
  wire popcount35_3d5j_core_219;
  wire popcount35_3d5j_core_220;
  wire popcount35_3d5j_core_222;
  wire popcount35_3d5j_core_223;
  wire popcount35_3d5j_core_225;
  wire popcount35_3d5j_core_227;
  wire popcount35_3d5j_core_229;
  wire popcount35_3d5j_core_230;
  wire popcount35_3d5j_core_234;
  wire popcount35_3d5j_core_235;
  wire popcount35_3d5j_core_236;
  wire popcount35_3d5j_core_238;
  wire popcount35_3d5j_core_240;
  wire popcount35_3d5j_core_241;
  wire popcount35_3d5j_core_242;
  wire popcount35_3d5j_core_243;
  wire popcount35_3d5j_core_244;
  wire popcount35_3d5j_core_247;
  wire popcount35_3d5j_core_248;
  wire popcount35_3d5j_core_250;
  wire popcount35_3d5j_core_252;
  wire popcount35_3d5j_core_253;
  wire popcount35_3d5j_core_254;
  wire popcount35_3d5j_core_255;
  wire popcount35_3d5j_core_256;
  wire popcount35_3d5j_core_257;
  wire popcount35_3d5j_core_258_not;
  wire popcount35_3d5j_core_259;
  wire popcount35_3d5j_core_260;
  wire popcount35_3d5j_core_261;
  wire popcount35_3d5j_core_262;
  wire popcount35_3d5j_core_264;

  assign popcount35_3d5j_core_037 = input_a[0] ^ input_a[1];
  assign popcount35_3d5j_core_038 = input_a[0] & input_a[1];
  assign popcount35_3d5j_core_039 = input_a[2] ^ input_a[3];
  assign popcount35_3d5j_core_040 = input_a[2] & input_a[3];
  assign popcount35_3d5j_core_041 = popcount35_3d5j_core_037 ^ popcount35_3d5j_core_039;
  assign popcount35_3d5j_core_042 = popcount35_3d5j_core_037 & popcount35_3d5j_core_039;
  assign popcount35_3d5j_core_043 = popcount35_3d5j_core_038 ^ popcount35_3d5j_core_040;
  assign popcount35_3d5j_core_044 = popcount35_3d5j_core_038 & input_a[2];
  assign popcount35_3d5j_core_045 = popcount35_3d5j_core_043 | popcount35_3d5j_core_042;
  assign popcount35_3d5j_core_048 = input_a[13] ^ input_a[12];
  assign popcount35_3d5j_core_049 = input_a[6] & input_a[12];
  assign popcount35_3d5j_core_050 = ~(input_a[6] & input_a[7]);
  assign popcount35_3d5j_core_051 = input_a[6] & input_a[7];
  assign popcount35_3d5j_core_052 = popcount35_3d5j_core_048 ^ popcount35_3d5j_core_050;
  assign popcount35_3d5j_core_054 = input_a[12] ^ popcount35_3d5j_core_051;
  assign popcount35_3d5j_core_055 = popcount35_3d5j_core_049 & input_a[13];
  assign popcount35_3d5j_core_056 = popcount35_3d5j_core_054 | popcount35_3d5j_core_048;
  assign popcount35_3d5j_core_057 = ~(input_a[19] & input_a[25]);
  assign popcount35_3d5j_core_060 = popcount35_3d5j_core_041 & popcount35_3d5j_core_052;
  assign popcount35_3d5j_core_061 = popcount35_3d5j_core_045 ^ popcount35_3d5j_core_056;
  assign popcount35_3d5j_core_062 = popcount35_3d5j_core_045 & popcount35_3d5j_core_056;
  assign popcount35_3d5j_core_063 = popcount35_3d5j_core_061 ^ popcount35_3d5j_core_060;
  assign popcount35_3d5j_core_064 = popcount35_3d5j_core_061 & popcount35_3d5j_core_060;
  assign popcount35_3d5j_core_065 = popcount35_3d5j_core_062 | popcount35_3d5j_core_064;
  assign popcount35_3d5j_core_066 = popcount35_3d5j_core_044 | popcount35_3d5j_core_055;
  assign popcount35_3d5j_core_067 = input_a[24] | input_a[8];
  assign popcount35_3d5j_core_068 = popcount35_3d5j_core_066 | popcount35_3d5j_core_065;
  assign popcount35_3d5j_core_070 = input_a[24] | input_a[23];
  assign popcount35_3d5j_core_072 = input_a[24] & input_a[28];
  assign popcount35_3d5j_core_073 = input_a[33] ^ input_a[29];
  assign popcount35_3d5j_core_074 = input_a[23] & input_a[15];
  assign popcount35_3d5j_core_076 = input_a[29] & input_a[4];
  assign popcount35_3d5j_core_077 = popcount35_3d5j_core_072 | popcount35_3d5j_core_074;
  assign popcount35_3d5j_core_078 = ~(input_a[22] ^ input_a[20]);
  assign popcount35_3d5j_core_079 = popcount35_3d5j_core_077 | popcount35_3d5j_core_076;
  assign popcount35_3d5j_core_082 = ~(input_a[5] & input_a[20]);
  assign popcount35_3d5j_core_083 = input_a[30] & input_a[17];
  assign popcount35_3d5j_core_084 = input_a[1] & input_a[6];
  assign popcount35_3d5j_core_085 = input_a[9] & input_a[33];
  assign popcount35_3d5j_core_086 = ~input_a[31];
  assign popcount35_3d5j_core_087 = input_a[22] & input_a[16];
  assign popcount35_3d5j_core_088 = popcount35_3d5j_core_085 | popcount35_3d5j_core_087;
  assign popcount35_3d5j_core_091 = input_a[27] & input_a[25];
  assign popcount35_3d5j_core_092 = popcount35_3d5j_core_083 ^ popcount35_3d5j_core_088;
  assign popcount35_3d5j_core_093 = popcount35_3d5j_core_083 & popcount35_3d5j_core_088;
  assign popcount35_3d5j_core_094 = popcount35_3d5j_core_092 ^ popcount35_3d5j_core_091;
  assign popcount35_3d5j_core_095 = popcount35_3d5j_core_092 & popcount35_3d5j_core_091;
  assign popcount35_3d5j_core_096 = popcount35_3d5j_core_093 | popcount35_3d5j_core_095;
  assign popcount35_3d5j_core_101 = popcount35_3d5j_core_079 ^ popcount35_3d5j_core_094;
  assign popcount35_3d5j_core_102 = popcount35_3d5j_core_079 & popcount35_3d5j_core_094;
  assign popcount35_3d5j_core_104 = input_a[15] ^ input_a[8];
  assign popcount35_3d5j_core_108 = popcount35_3d5j_core_096 | popcount35_3d5j_core_102;
  assign popcount35_3d5j_core_109 = ~(input_a[27] | input_a[4]);
  assign popcount35_3d5j_core_111 = input_a[30] ^ input_a[30];
  assign popcount35_3d5j_core_114 = input_a[34] & input_a[31];
  assign popcount35_3d5j_core_115 = popcount35_3d5j_core_063 ^ popcount35_3d5j_core_101;
  assign popcount35_3d5j_core_116 = popcount35_3d5j_core_063 & popcount35_3d5j_core_101;
  assign popcount35_3d5j_core_117 = popcount35_3d5j_core_115 ^ popcount35_3d5j_core_114;
  assign popcount35_3d5j_core_118 = popcount35_3d5j_core_115 & popcount35_3d5j_core_114;
  assign popcount35_3d5j_core_119 = popcount35_3d5j_core_116 | popcount35_3d5j_core_118;
  assign popcount35_3d5j_core_120 = popcount35_3d5j_core_068 ^ popcount35_3d5j_core_108;
  assign popcount35_3d5j_core_121 = popcount35_3d5j_core_068 & popcount35_3d5j_core_108;
  assign popcount35_3d5j_core_122 = popcount35_3d5j_core_120 ^ popcount35_3d5j_core_119;
  assign popcount35_3d5j_core_123 = popcount35_3d5j_core_120 & popcount35_3d5j_core_119;
  assign popcount35_3d5j_core_124 = popcount35_3d5j_core_121 | popcount35_3d5j_core_123;
  assign popcount35_3d5j_core_128 = input_a[25] ^ input_a[9];
  assign popcount35_3d5j_core_129 = ~input_a[11];
  assign popcount35_3d5j_core_130 = ~(input_a[12] ^ input_a[27]);
  assign popcount35_3d5j_core_131 = ~(input_a[2] ^ input_a[32]);
  assign popcount35_3d5j_core_132 = input_a[6] & input_a[32];
  assign popcount35_3d5j_core_134 = ~(input_a[20] ^ input_a[31]);
  assign popcount35_3d5j_core_137 = ~(input_a[27] & input_a[14]);
  assign popcount35_3d5j_core_139 = input_a[30] | input_a[2];
  assign popcount35_3d5j_core_140 = ~input_a[13];
  assign popcount35_3d5j_core_142 = ~(input_a[20] ^ input_a[31]);
  assign popcount35_3d5j_core_143 = ~(input_a[2] ^ input_a[20]);
  assign popcount35_3d5j_core_144 = ~(input_a[24] & input_a[10]);
  assign popcount35_3d5j_core_146 = ~input_a[3];
  assign popcount35_3d5j_core_148 = input_a[33] ^ input_a[11];
  assign popcount35_3d5j_core_149 = ~input_a[27];
  assign popcount35_3d5j_core_150 = ~(input_a[1] & input_a[27]);
  assign popcount35_3d5j_core_151 = input_a[3] | input_a[22];
  assign popcount35_3d5j_core_152 = ~(input_a[26] | input_a[10]);
  assign popcount35_3d5j_core_155 = input_a[12] ^ input_a[27];
  assign popcount35_3d5j_core_156 = input_a[16] | input_a[3];
  assign popcount35_3d5j_core_157 = input_a[9] | input_a[31];
  assign popcount35_3d5j_core_158 = input_a[24] & input_a[19];
  assign popcount35_3d5j_core_159 = ~(input_a[0] ^ input_a[29]);
  assign popcount35_3d5j_core_162 = ~(input_a[2] ^ input_a[14]);
  assign popcount35_3d5j_core_163 = ~(input_a[24] & input_a[33]);
  assign popcount35_3d5j_core_164 = input_a[20] ^ input_a[25];
  assign popcount35_3d5j_core_166 = ~(input_a[6] & input_a[5]);
  assign popcount35_3d5j_core_170 = input_a[26] | input_a[8];
  assign popcount35_3d5j_core_171 = ~(input_a[3] & input_a[12]);
  assign popcount35_3d5j_core_173 = input_a[10] & input_a[26];
  assign popcount35_3d5j_core_174 = input_a[5] ^ input_a[22];
  assign popcount35_3d5j_core_175 = input_a[31] | input_a[34];
  assign popcount35_3d5j_core_176 = ~(input_a[12] ^ input_a[0]);
  assign popcount35_3d5j_core_177_not = ~input_a[10];
  assign popcount35_3d5j_core_178 = input_a[28] | input_a[5];
  assign popcount35_3d5j_core_179 = ~(input_a[34] ^ input_a[22]);
  assign popcount35_3d5j_core_180 = ~(input_a[2] & input_a[5]);
  assign popcount35_3d5j_core_182 = input_a[6] ^ input_a[15];
  assign popcount35_3d5j_core_184 = ~(input_a[12] & input_a[30]);
  assign popcount35_3d5j_core_185 = ~(input_a[17] ^ input_a[25]);
  assign popcount35_3d5j_core_188 = ~(input_a[22] | input_a[33]);
  assign popcount35_3d5j_core_190 = ~(input_a[9] ^ input_a[12]);
  assign popcount35_3d5j_core_192 = ~(input_a[19] | input_a[20]);
  assign popcount35_3d5j_core_193 = input_a[16] & input_a[13];
  assign popcount35_3d5j_core_194 = ~(input_a[27] ^ input_a[7]);
  assign popcount35_3d5j_core_195 = input_a[19] ^ input_a[1];
  assign popcount35_3d5j_core_197 = ~(input_a[24] & input_a[2]);
  assign popcount35_3d5j_core_198 = input_a[6] | input_a[6];
  assign popcount35_3d5j_core_200 = ~(input_a[16] ^ input_a[29]);
  assign popcount35_3d5j_core_201 = input_a[15] | input_a[6];
  assign popcount35_3d5j_core_203 = ~(input_a[0] & input_a[3]);
  assign popcount35_3d5j_core_204 = ~(input_a[15] | input_a[20]);
  assign popcount35_3d5j_core_205 = ~input_a[13];
  assign popcount35_3d5j_core_206 = ~(input_a[1] | input_a[34]);
  assign popcount35_3d5j_core_207 = input_a[28] | input_a[17];
  assign popcount35_3d5j_core_209 = input_a[29] | input_a[33];
  assign popcount35_3d5j_core_211 = input_a[12] | input_a[8];
  assign popcount35_3d5j_core_212 = input_a[29] | input_a[6];
  assign popcount35_3d5j_core_213 = ~(input_a[10] ^ input_a[28]);
  assign popcount35_3d5j_core_214 = ~input_a[3];
  assign popcount35_3d5j_core_215 = input_a[27] | input_a[4];
  assign popcount35_3d5j_core_217 = input_a[34] ^ input_a[17];
  assign popcount35_3d5j_core_218 = ~(input_a[8] | input_a[18]);
  assign popcount35_3d5j_core_219 = input_a[14] | input_a[33];
  assign popcount35_3d5j_core_220 = input_a[18] & input_a[19];
  assign popcount35_3d5j_core_222 = ~(input_a[0] | input_a[27]);
  assign popcount35_3d5j_core_223 = ~input_a[4];
  assign popcount35_3d5j_core_225 = ~(input_a[6] | input_a[22]);
  assign popcount35_3d5j_core_227 = input_a[6] ^ input_a[33];
  assign popcount35_3d5j_core_229 = ~(input_a[6] ^ input_a[26]);
  assign popcount35_3d5j_core_230 = ~input_a[23];
  assign popcount35_3d5j_core_234 = input_a[25] ^ input_a[33];
  assign popcount35_3d5j_core_235 = ~(input_a[9] | input_a[6]);
  assign popcount35_3d5j_core_236 = ~(input_a[13] & input_a[33]);
  assign popcount35_3d5j_core_238 = ~(input_a[29] & input_a[4]);
  assign popcount35_3d5j_core_240 = popcount35_3d5j_core_117 ^ popcount35_3d5j_core_220;
  assign popcount35_3d5j_core_241 = popcount35_3d5j_core_117 & popcount35_3d5j_core_220;
  assign popcount35_3d5j_core_242 = popcount35_3d5j_core_240 ^ input_a[21];
  assign popcount35_3d5j_core_243 = popcount35_3d5j_core_240 & input_a[21];
  assign popcount35_3d5j_core_244 = popcount35_3d5j_core_241 | popcount35_3d5j_core_243;
  assign popcount35_3d5j_core_247 = popcount35_3d5j_core_122 ^ popcount35_3d5j_core_244;
  assign popcount35_3d5j_core_248 = popcount35_3d5j_core_122 & popcount35_3d5j_core_244;
  assign popcount35_3d5j_core_250 = ~popcount35_3d5j_core_124;
  assign popcount35_3d5j_core_252 = popcount35_3d5j_core_250 ^ popcount35_3d5j_core_248;
  assign popcount35_3d5j_core_253 = popcount35_3d5j_core_250 & popcount35_3d5j_core_248;
  assign popcount35_3d5j_core_254 = popcount35_3d5j_core_124 | popcount35_3d5j_core_253;
  assign popcount35_3d5j_core_255 = ~(input_a[29] ^ input_a[17]);
  assign popcount35_3d5j_core_256 = input_a[10] & input_a[31];
  assign popcount35_3d5j_core_257 = ~(input_a[15] & input_a[34]);
  assign popcount35_3d5j_core_258_not = ~input_a[28];
  assign popcount35_3d5j_core_259 = ~(input_a[5] | input_a[26]);
  assign popcount35_3d5j_core_260 = ~(input_a[29] | input_a[19]);
  assign popcount35_3d5j_core_261 = ~(input_a[27] ^ input_a[25]);
  assign popcount35_3d5j_core_262 = input_a[21] ^ input_a[0];
  assign popcount35_3d5j_core_264 = ~(input_a[4] | input_a[21]);

  assign popcount35_3d5j_out[0] = input_a[5];
  assign popcount35_3d5j_out[1] = popcount35_3d5j_core_242;
  assign popcount35_3d5j_out[2] = popcount35_3d5j_core_247;
  assign popcount35_3d5j_out[3] = popcount35_3d5j_core_252;
  assign popcount35_3d5j_out[4] = popcount35_3d5j_core_254;
  assign popcount35_3d5j_out[5] = 1'b0;
endmodule