// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.35385
// WCE=19.0
// EP=0.892489%
// Printed PDK parameters:
//  Area=78058625.0
//  Delay=88491568.0
//  Power=3812100.0

module popcount38_sjm1(input [37:0] input_a, output [5:0] popcount38_sjm1_out);
  wire popcount38_sjm1_core_040;
  wire popcount38_sjm1_core_041;
  wire popcount38_sjm1_core_046;
  wire popcount38_sjm1_core_047;
  wire popcount38_sjm1_core_049;
  wire popcount38_sjm1_core_051;
  wire popcount38_sjm1_core_052;
  wire popcount38_sjm1_core_053;
  wire popcount38_sjm1_core_055;
  wire popcount38_sjm1_core_056;
  wire popcount38_sjm1_core_057;
  wire popcount38_sjm1_core_059;
  wire popcount38_sjm1_core_060;
  wire popcount38_sjm1_core_061;
  wire popcount38_sjm1_core_062;
  wire popcount38_sjm1_core_063;
  wire popcount38_sjm1_core_064;
  wire popcount38_sjm1_core_068;
  wire popcount38_sjm1_core_069;
  wire popcount38_sjm1_core_070;
  wire popcount38_sjm1_core_071;
  wire popcount38_sjm1_core_072;
  wire popcount38_sjm1_core_073;
  wire popcount38_sjm1_core_074;
  wire popcount38_sjm1_core_075;
  wire popcount38_sjm1_core_076;
  wire popcount38_sjm1_core_077;
  wire popcount38_sjm1_core_078;
  wire popcount38_sjm1_core_079;
  wire popcount38_sjm1_core_081;
  wire popcount38_sjm1_core_082;
  wire popcount38_sjm1_core_083;
  wire popcount38_sjm1_core_084;
  wire popcount38_sjm1_core_085;
  wire popcount38_sjm1_core_086;
  wire popcount38_sjm1_core_087;
  wire popcount38_sjm1_core_088;
  wire popcount38_sjm1_core_089;
  wire popcount38_sjm1_core_090;
  wire popcount38_sjm1_core_091;
  wire popcount38_sjm1_core_092;
  wire popcount38_sjm1_core_093;
  wire popcount38_sjm1_core_094;
  wire popcount38_sjm1_core_095;
  wire popcount38_sjm1_core_096;
  wire popcount38_sjm1_core_097;
  wire popcount38_sjm1_core_099;
  wire popcount38_sjm1_core_105;
  wire popcount38_sjm1_core_107;
  wire popcount38_sjm1_core_108;
  wire popcount38_sjm1_core_109;
  wire popcount38_sjm1_core_110;
  wire popcount38_sjm1_core_112;
  wire popcount38_sjm1_core_113;
  wire popcount38_sjm1_core_116;
  wire popcount38_sjm1_core_117;
  wire popcount38_sjm1_core_118;
  wire popcount38_sjm1_core_119;
  wire popcount38_sjm1_core_120;
  wire popcount38_sjm1_core_121;
  wire popcount38_sjm1_core_122;
  wire popcount38_sjm1_core_125;
  wire popcount38_sjm1_core_126;
  wire popcount38_sjm1_core_131;
  wire popcount38_sjm1_core_133;
  wire popcount38_sjm1_core_134;
  wire popcount38_sjm1_core_135;
  wire popcount38_sjm1_core_136;
  wire popcount38_sjm1_core_137;
  wire popcount38_sjm1_core_138;
  wire popcount38_sjm1_core_139;
  wire popcount38_sjm1_core_140;
  wire popcount38_sjm1_core_141;
  wire popcount38_sjm1_core_142;
  wire popcount38_sjm1_core_143;
  wire popcount38_sjm1_core_144;
  wire popcount38_sjm1_core_145;
  wire popcount38_sjm1_core_146;
  wire popcount38_sjm1_core_147;
  wire popcount38_sjm1_core_148;
  wire popcount38_sjm1_core_149;
  wire popcount38_sjm1_core_151;
  wire popcount38_sjm1_core_153;
  wire popcount38_sjm1_core_155;
  wire popcount38_sjm1_core_156;
  wire popcount38_sjm1_core_157;
  wire popcount38_sjm1_core_158;
  wire popcount38_sjm1_core_159;
  wire popcount38_sjm1_core_162;
  wire popcount38_sjm1_core_167;
  wire popcount38_sjm1_core_168;
  wire popcount38_sjm1_core_169;
  wire popcount38_sjm1_core_171;
  wire popcount38_sjm1_core_172;
  wire popcount38_sjm1_core_174;
  wire popcount38_sjm1_core_175;
  wire popcount38_sjm1_core_177;
  wire popcount38_sjm1_core_178;
  wire popcount38_sjm1_core_179;
  wire popcount38_sjm1_core_180;
  wire popcount38_sjm1_core_184;
  wire popcount38_sjm1_core_186;
  wire popcount38_sjm1_core_188;
  wire popcount38_sjm1_core_197;
  wire popcount38_sjm1_core_198;
  wire popcount38_sjm1_core_199;
  wire popcount38_sjm1_core_200;
  wire popcount38_sjm1_core_203;
  wire popcount38_sjm1_core_204;
  wire popcount38_sjm1_core_205;
  wire popcount38_sjm1_core_207;
  wire popcount38_sjm1_core_208;
  wire popcount38_sjm1_core_209;
  wire popcount38_sjm1_core_212;
  wire popcount38_sjm1_core_214;
  wire popcount38_sjm1_core_215;
  wire popcount38_sjm1_core_216;
  wire popcount38_sjm1_core_217;
  wire popcount38_sjm1_core_218;
  wire popcount38_sjm1_core_219;
  wire popcount38_sjm1_core_220;
  wire popcount38_sjm1_core_222;
  wire popcount38_sjm1_core_223;
  wire popcount38_sjm1_core_224;
  wire popcount38_sjm1_core_225;
  wire popcount38_sjm1_core_226;
  wire popcount38_sjm1_core_227;
  wire popcount38_sjm1_core_228;
  wire popcount38_sjm1_core_231;
  wire popcount38_sjm1_core_232;
  wire popcount38_sjm1_core_233;
  wire popcount38_sjm1_core_234;
  wire popcount38_sjm1_core_236;
  wire popcount38_sjm1_core_237;
  wire popcount38_sjm1_core_238;
  wire popcount38_sjm1_core_239;
  wire popcount38_sjm1_core_240;
  wire popcount38_sjm1_core_241;
  wire popcount38_sjm1_core_242;
  wire popcount38_sjm1_core_246;
  wire popcount38_sjm1_core_248;
  wire popcount38_sjm1_core_251;
  wire popcount38_sjm1_core_253;
  wire popcount38_sjm1_core_255_not;
  wire popcount38_sjm1_core_256;
  wire popcount38_sjm1_core_257;
  wire popcount38_sjm1_core_260;
  wire popcount38_sjm1_core_261;
  wire popcount38_sjm1_core_262_not;
  wire popcount38_sjm1_core_264;
  wire popcount38_sjm1_core_266;
  wire popcount38_sjm1_core_268;
  wire popcount38_sjm1_core_270;
  wire popcount38_sjm1_core_271;
  wire popcount38_sjm1_core_274;
  wire popcount38_sjm1_core_275;
  wire popcount38_sjm1_core_277;
  wire popcount38_sjm1_core_278;
  wire popcount38_sjm1_core_279;
  wire popcount38_sjm1_core_280;
  wire popcount38_sjm1_core_281;
  wire popcount38_sjm1_core_282;
  wire popcount38_sjm1_core_283;
  wire popcount38_sjm1_core_284;
  wire popcount38_sjm1_core_285;
  wire popcount38_sjm1_core_286;
  wire popcount38_sjm1_core_287;
  wire popcount38_sjm1_core_288;
  wire popcount38_sjm1_core_289;
  wire popcount38_sjm1_core_290;
  wire popcount38_sjm1_core_291;

  assign popcount38_sjm1_core_040 = input_a[0] ^ input_a[1];
  assign popcount38_sjm1_core_041 = input_a[0] & input_a[1];
  assign popcount38_sjm1_core_046 = popcount38_sjm1_core_041 ^ input_a[16];
  assign popcount38_sjm1_core_047 = popcount38_sjm1_core_041 & input_a[16];
  assign popcount38_sjm1_core_049 = ~(input_a[8] & input_a[21]);
  assign popcount38_sjm1_core_051 = input_a[4] ^ input_a[5];
  assign popcount38_sjm1_core_052 = input_a[4] & input_a[5];
  assign popcount38_sjm1_core_053 = input_a[7] ^ input_a[23];
  assign popcount38_sjm1_core_055 = input_a[6] & popcount38_sjm1_core_053;
  assign popcount38_sjm1_core_056 = input_a[6] & popcount38_sjm1_core_053;
  assign popcount38_sjm1_core_057 = input_a[34] ^ popcount38_sjm1_core_056;
  assign popcount38_sjm1_core_059 = popcount38_sjm1_core_051 ^ popcount38_sjm1_core_055;
  assign popcount38_sjm1_core_060 = popcount38_sjm1_core_051 & popcount38_sjm1_core_055;
  assign popcount38_sjm1_core_061 = popcount38_sjm1_core_052 ^ popcount38_sjm1_core_057;
  assign popcount38_sjm1_core_062 = popcount38_sjm1_core_052 & popcount38_sjm1_core_057;
  assign popcount38_sjm1_core_063 = popcount38_sjm1_core_061 ^ popcount38_sjm1_core_060;
  assign popcount38_sjm1_core_064 = ~input_a[36];
  assign popcount38_sjm1_core_068 = input_a[14] ^ popcount38_sjm1_core_059;
  assign popcount38_sjm1_core_069 = input_a[14] & popcount38_sjm1_core_059;
  assign popcount38_sjm1_core_070 = popcount38_sjm1_core_046 ^ popcount38_sjm1_core_063;
  assign popcount38_sjm1_core_071 = popcount38_sjm1_core_046 & popcount38_sjm1_core_063;
  assign popcount38_sjm1_core_072 = popcount38_sjm1_core_070 ^ popcount38_sjm1_core_069;
  assign popcount38_sjm1_core_073 = popcount38_sjm1_core_070 & popcount38_sjm1_core_069;
  assign popcount38_sjm1_core_074 = popcount38_sjm1_core_071 | popcount38_sjm1_core_073;
  assign popcount38_sjm1_core_075 = popcount38_sjm1_core_047 ^ popcount38_sjm1_core_062;
  assign popcount38_sjm1_core_076 = popcount38_sjm1_core_047 & popcount38_sjm1_core_062;
  assign popcount38_sjm1_core_077 = popcount38_sjm1_core_075 ^ popcount38_sjm1_core_074;
  assign popcount38_sjm1_core_078 = popcount38_sjm1_core_075 & popcount38_sjm1_core_074;
  assign popcount38_sjm1_core_079 = popcount38_sjm1_core_076 | popcount38_sjm1_core_078;
  assign popcount38_sjm1_core_081 = ~(input_a[34] | input_a[6]);
  assign popcount38_sjm1_core_082 = input_a[9] ^ input_a[10];
  assign popcount38_sjm1_core_083 = input_a[9] & input_a[10];
  assign popcount38_sjm1_core_084 = input_a[12] ^ input_a[13];
  assign popcount38_sjm1_core_085 = input_a[12] & input_a[13];
  assign popcount38_sjm1_core_086 = input_a[11] ^ popcount38_sjm1_core_084;
  assign popcount38_sjm1_core_087 = input_a[11] & popcount38_sjm1_core_084;
  assign popcount38_sjm1_core_088 = popcount38_sjm1_core_085 ^ popcount38_sjm1_core_087;
  assign popcount38_sjm1_core_089 = popcount38_sjm1_core_085 & popcount38_sjm1_core_087;
  assign popcount38_sjm1_core_090 = popcount38_sjm1_core_082 ^ popcount38_sjm1_core_086;
  assign popcount38_sjm1_core_091 = popcount38_sjm1_core_082 & popcount38_sjm1_core_086;
  assign popcount38_sjm1_core_092 = popcount38_sjm1_core_083 ^ popcount38_sjm1_core_088;
  assign popcount38_sjm1_core_093 = popcount38_sjm1_core_083 & popcount38_sjm1_core_088;
  assign popcount38_sjm1_core_094 = popcount38_sjm1_core_092 ^ popcount38_sjm1_core_091;
  assign popcount38_sjm1_core_095 = popcount38_sjm1_core_092 & popcount38_sjm1_core_091;
  assign popcount38_sjm1_core_096 = popcount38_sjm1_core_093 | popcount38_sjm1_core_095;
  assign popcount38_sjm1_core_097 = popcount38_sjm1_core_089 ^ popcount38_sjm1_core_096;
  assign popcount38_sjm1_core_099 = ~(input_a[33] | input_a[33]);
  assign popcount38_sjm1_core_105 = input_a[11] ^ input_a[37];
  assign popcount38_sjm1_core_107 = ~(popcount38_sjm1_core_099 & input_a[27]);
  assign popcount38_sjm1_core_108 = ~(input_a[18] | input_a[3]);
  assign popcount38_sjm1_core_109 = input_a[4] | input_a[35];
  assign popcount38_sjm1_core_110 = input_a[8] ^ input_a[16];
  assign popcount38_sjm1_core_112 = ~input_a[37];
  assign popcount38_sjm1_core_113 = ~input_a[34];
  assign popcount38_sjm1_core_116 = popcount38_sjm1_core_090 ^ popcount38_sjm1_core_107;
  assign popcount38_sjm1_core_117 = popcount38_sjm1_core_090 & popcount38_sjm1_core_107;
  assign popcount38_sjm1_core_118 = popcount38_sjm1_core_094 ^ input_a[27];
  assign popcount38_sjm1_core_119 = popcount38_sjm1_core_094 & input_a[27];
  assign popcount38_sjm1_core_120 = popcount38_sjm1_core_118 ^ popcount38_sjm1_core_117;
  assign popcount38_sjm1_core_121 = popcount38_sjm1_core_118 & popcount38_sjm1_core_117;
  assign popcount38_sjm1_core_122 = popcount38_sjm1_core_119 | popcount38_sjm1_core_121;
  assign popcount38_sjm1_core_125 = popcount38_sjm1_core_097 ^ popcount38_sjm1_core_122;
  assign popcount38_sjm1_core_126 = popcount38_sjm1_core_097 & popcount38_sjm1_core_122;
  assign popcount38_sjm1_core_131 = input_a[0] | input_a[36];
  assign popcount38_sjm1_core_133 = popcount38_sjm1_core_068 ^ popcount38_sjm1_core_116;
  assign popcount38_sjm1_core_134 = popcount38_sjm1_core_068 & popcount38_sjm1_core_116;
  assign popcount38_sjm1_core_135 = popcount38_sjm1_core_072 ^ popcount38_sjm1_core_120;
  assign popcount38_sjm1_core_136 = popcount38_sjm1_core_072 & popcount38_sjm1_core_120;
  assign popcount38_sjm1_core_137 = popcount38_sjm1_core_135 ^ popcount38_sjm1_core_134;
  assign popcount38_sjm1_core_138 = popcount38_sjm1_core_135 & popcount38_sjm1_core_134;
  assign popcount38_sjm1_core_139 = popcount38_sjm1_core_136 | popcount38_sjm1_core_138;
  assign popcount38_sjm1_core_140 = popcount38_sjm1_core_077 ^ popcount38_sjm1_core_125;
  assign popcount38_sjm1_core_141 = popcount38_sjm1_core_077 & popcount38_sjm1_core_125;
  assign popcount38_sjm1_core_142 = popcount38_sjm1_core_140 ^ popcount38_sjm1_core_139;
  assign popcount38_sjm1_core_143 = popcount38_sjm1_core_140 & popcount38_sjm1_core_139;
  assign popcount38_sjm1_core_144 = popcount38_sjm1_core_141 | popcount38_sjm1_core_143;
  assign popcount38_sjm1_core_145 = popcount38_sjm1_core_079 ^ popcount38_sjm1_core_126;
  assign popcount38_sjm1_core_146 = popcount38_sjm1_core_079 & popcount38_sjm1_core_126;
  assign popcount38_sjm1_core_147 = popcount38_sjm1_core_145 ^ popcount38_sjm1_core_144;
  assign popcount38_sjm1_core_148 = popcount38_sjm1_core_145 & popcount38_sjm1_core_144;
  assign popcount38_sjm1_core_149 = popcount38_sjm1_core_146 | popcount38_sjm1_core_148;
  assign popcount38_sjm1_core_151 = input_a[6] ^ input_a[15];
  assign popcount38_sjm1_core_153 = input_a[14] ^ input_a[30];
  assign popcount38_sjm1_core_155 = ~(input_a[32] ^ input_a[20]);
  assign popcount38_sjm1_core_156 = input_a[19] & input_a[20];
  assign popcount38_sjm1_core_157 = ~(input_a[21] & input_a[22]);
  assign popcount38_sjm1_core_158 = input_a[21] & input_a[22];
  assign popcount38_sjm1_core_159 = input_a[9] ^ input_a[13];
  assign popcount38_sjm1_core_162 = popcount38_sjm1_core_156 & popcount38_sjm1_core_158;
  assign popcount38_sjm1_core_167 = input_a[4] | input_a[13];
  assign popcount38_sjm1_core_168 = ~(input_a[0] ^ input_a[24]);
  assign popcount38_sjm1_core_169 = ~(input_a[16] & input_a[32]);
  assign popcount38_sjm1_core_171 = ~(input_a[21] ^ input_a[5]);
  assign popcount38_sjm1_core_172 = ~input_a[2];
  assign popcount38_sjm1_core_174 = input_a[35] & input_a[16];
  assign popcount38_sjm1_core_175 = input_a[36] | input_a[33];
  assign popcount38_sjm1_core_177 = input_a[9] | input_a[16];
  assign popcount38_sjm1_core_178 = input_a[33] | popcount38_sjm1_core_175;
  assign popcount38_sjm1_core_179 = ~input_a[21];
  assign popcount38_sjm1_core_180 = input_a[30] & input_a[26];
  assign popcount38_sjm1_core_184 = input_a[33] & input_a[30];
  assign popcount38_sjm1_core_186 = input_a[26] ^ input_a[7];
  assign popcount38_sjm1_core_188 = ~(input_a[3] ^ input_a[27]);
  assign popcount38_sjm1_core_197 = input_a[28] ^ input_a[25];
  assign popcount38_sjm1_core_198 = input_a[15] & input_a[29];
  assign popcount38_sjm1_core_199 = input_a[37] & input_a[1];
  assign popcount38_sjm1_core_200 = input_a[31] & input_a[32];
  assign popcount38_sjm1_core_203 = popcount38_sjm1_core_200 ^ input_a[30];
  assign popcount38_sjm1_core_204 = popcount38_sjm1_core_200 & input_a[30];
  assign popcount38_sjm1_core_205 = input_a[35] ^ input_a[10];
  assign popcount38_sjm1_core_207 = popcount38_sjm1_core_198 ^ popcount38_sjm1_core_203;
  assign popcount38_sjm1_core_208 = popcount38_sjm1_core_198 & popcount38_sjm1_core_203;
  assign popcount38_sjm1_core_209 = popcount38_sjm1_core_207 ^ input_a[3];
  assign popcount38_sjm1_core_212 = popcount38_sjm1_core_204 | popcount38_sjm1_core_208;
  assign popcount38_sjm1_core_214 = input_a[33] ^ input_a[34];
  assign popcount38_sjm1_core_215 = ~(input_a[33] | input_a[34]);
  assign popcount38_sjm1_core_216 = input_a[36] ^ input_a[37];
  assign popcount38_sjm1_core_217 = input_a[36] & input_a[37];
  assign popcount38_sjm1_core_218 = input_a[35] ^ popcount38_sjm1_core_216;
  assign popcount38_sjm1_core_219 = input_a[26] & popcount38_sjm1_core_216;
  assign popcount38_sjm1_core_220 = popcount38_sjm1_core_217 ^ popcount38_sjm1_core_219;
  assign popcount38_sjm1_core_222 = ~(popcount38_sjm1_core_214 & input_a[25]);
  assign popcount38_sjm1_core_223 = popcount38_sjm1_core_214 & popcount38_sjm1_core_218;
  assign popcount38_sjm1_core_224 = popcount38_sjm1_core_215 ^ popcount38_sjm1_core_220;
  assign popcount38_sjm1_core_225 = popcount38_sjm1_core_215 & popcount38_sjm1_core_220;
  assign popcount38_sjm1_core_226 = popcount38_sjm1_core_224 ^ popcount38_sjm1_core_223;
  assign popcount38_sjm1_core_227 = popcount38_sjm1_core_224 & popcount38_sjm1_core_223;
  assign popcount38_sjm1_core_228 = popcount38_sjm1_core_225 | popcount38_sjm1_core_227;
  assign popcount38_sjm1_core_231 = input_a[5] | input_a[21];
  assign popcount38_sjm1_core_232 = input_a[23] & input_a[8];
  assign popcount38_sjm1_core_233 = input_a[3] & popcount38_sjm1_core_226;
  assign popcount38_sjm1_core_234 = popcount38_sjm1_core_209 & popcount38_sjm1_core_226;
  assign popcount38_sjm1_core_236 = popcount38_sjm1_core_233 & input_a[33];
  assign popcount38_sjm1_core_237 = popcount38_sjm1_core_234 | popcount38_sjm1_core_236;
  assign popcount38_sjm1_core_238 = popcount38_sjm1_core_212 ^ popcount38_sjm1_core_228;
  assign popcount38_sjm1_core_239 = popcount38_sjm1_core_212 & popcount38_sjm1_core_228;
  assign popcount38_sjm1_core_240 = popcount38_sjm1_core_238 ^ popcount38_sjm1_core_237;
  assign popcount38_sjm1_core_241 = popcount38_sjm1_core_238 & popcount38_sjm1_core_237;
  assign popcount38_sjm1_core_242 = popcount38_sjm1_core_239 | popcount38_sjm1_core_241;
  assign popcount38_sjm1_core_246 = ~input_a[11];
  assign popcount38_sjm1_core_248 = input_a[26] ^ input_a[35];
  assign popcount38_sjm1_core_251 = ~(input_a[20] & input_a[22]);
  assign popcount38_sjm1_core_253 = ~(input_a[23] & input_a[30]);
  assign popcount38_sjm1_core_255_not = ~popcount38_sjm1_core_240;
  assign popcount38_sjm1_core_256 = input_a[12] & input_a[9];
  assign popcount38_sjm1_core_257 = ~popcount38_sjm1_core_255_not;
  assign popcount38_sjm1_core_260 = popcount38_sjm1_core_162 ^ popcount38_sjm1_core_242;
  assign popcount38_sjm1_core_261 = popcount38_sjm1_core_162 & popcount38_sjm1_core_242;
  assign popcount38_sjm1_core_262_not = ~popcount38_sjm1_core_260;
  assign popcount38_sjm1_core_264 = popcount38_sjm1_core_261 | popcount38_sjm1_core_260;
  assign popcount38_sjm1_core_266 = input_a[18] & input_a[21];
  assign popcount38_sjm1_core_268 = input_a[2] & input_a[13];
  assign popcount38_sjm1_core_270 = ~input_a[25];
  assign popcount38_sjm1_core_271 = input_a[2] & popcount38_sjm1_core_248;
  assign popcount38_sjm1_core_274 = popcount38_sjm1_core_137 ^ popcount38_sjm1_core_271;
  assign popcount38_sjm1_core_275 = popcount38_sjm1_core_137 & popcount38_sjm1_core_271;
  assign popcount38_sjm1_core_277 = popcount38_sjm1_core_142 ^ popcount38_sjm1_core_257;
  assign popcount38_sjm1_core_278 = popcount38_sjm1_core_142 & popcount38_sjm1_core_257;
  assign popcount38_sjm1_core_279 = popcount38_sjm1_core_277 ^ popcount38_sjm1_core_275;
  assign popcount38_sjm1_core_280 = popcount38_sjm1_core_277 & popcount38_sjm1_core_275;
  assign popcount38_sjm1_core_281 = popcount38_sjm1_core_278 | popcount38_sjm1_core_280;
  assign popcount38_sjm1_core_282 = popcount38_sjm1_core_147 ^ popcount38_sjm1_core_262_not;
  assign popcount38_sjm1_core_283 = popcount38_sjm1_core_147 & popcount38_sjm1_core_262_not;
  assign popcount38_sjm1_core_284 = input_a[33] ^ input_a[14];
  assign popcount38_sjm1_core_285 = popcount38_sjm1_core_282 & popcount38_sjm1_core_281;
  assign popcount38_sjm1_core_286 = popcount38_sjm1_core_283 | popcount38_sjm1_core_285;
  assign popcount38_sjm1_core_287 = popcount38_sjm1_core_149 ^ popcount38_sjm1_core_264;
  assign popcount38_sjm1_core_288 = popcount38_sjm1_core_149 & popcount38_sjm1_core_264;
  assign popcount38_sjm1_core_289 = popcount38_sjm1_core_287 ^ popcount38_sjm1_core_286;
  assign popcount38_sjm1_core_290 = popcount38_sjm1_core_287 & popcount38_sjm1_core_286;
  assign popcount38_sjm1_core_291 = popcount38_sjm1_core_288 | popcount38_sjm1_core_290;

  assign popcount38_sjm1_out[0] = popcount38_sjm1_core_040;
  assign popcount38_sjm1_out[1] = popcount38_sjm1_core_274;
  assign popcount38_sjm1_out[2] = popcount38_sjm1_core_279;
  assign popcount38_sjm1_out[3] = 1'b0;
  assign popcount38_sjm1_out[4] = popcount38_sjm1_core_289;
  assign popcount38_sjm1_out[5] = popcount38_sjm1_core_291;
endmodule