// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.12771
// WCE=50.0
// EP=0.964124%
// Printed PDK parameters:
//  Area=61865092.0
//  Delay=63190568.0
//  Power=3030300.0

module popcount47_i2df(input [46:0] input_a, output [5:0] popcount47_i2df_out);
  wire popcount47_i2df_core_049;
  wire popcount47_i2df_core_050;
  wire popcount47_i2df_core_051;
  wire popcount47_i2df_core_052;
  wire popcount47_i2df_core_054;
  wire popcount47_i2df_core_056;
  wire popcount47_i2df_core_057_not;
  wire popcount47_i2df_core_062;
  wire popcount47_i2df_core_064;
  wire popcount47_i2df_core_065;
  wire popcount47_i2df_core_068;
  wire popcount47_i2df_core_069;
  wire popcount47_i2df_core_073;
  wire popcount47_i2df_core_079;
  wire popcount47_i2df_core_080_not;
  wire popcount47_i2df_core_081;
  wire popcount47_i2df_core_082;
  wire popcount47_i2df_core_083;
  wire popcount47_i2df_core_090;
  wire popcount47_i2df_core_091;
  wire popcount47_i2df_core_092;
  wire popcount47_i2df_core_094;
  wire popcount47_i2df_core_095;
  wire popcount47_i2df_core_096;
  wire popcount47_i2df_core_099;
  wire popcount47_i2df_core_100;
  wire popcount47_i2df_core_101;
  wire popcount47_i2df_core_104;
  wire popcount47_i2df_core_105;
  wire popcount47_i2df_core_107;
  wire popcount47_i2df_core_108;
  wire popcount47_i2df_core_109;
  wire popcount47_i2df_core_110;
  wire popcount47_i2df_core_111;
  wire popcount47_i2df_core_112;
  wire popcount47_i2df_core_113;
  wire popcount47_i2df_core_114;
  wire popcount47_i2df_core_115;
  wire popcount47_i2df_core_116;
  wire popcount47_i2df_core_117;
  wire popcount47_i2df_core_118;
  wire popcount47_i2df_core_119;
  wire popcount47_i2df_core_120;
  wire popcount47_i2df_core_121;
  wire popcount47_i2df_core_122;
  wire popcount47_i2df_core_123;
  wire popcount47_i2df_core_124;
  wire popcount47_i2df_core_125;
  wire popcount47_i2df_core_126;
  wire popcount47_i2df_core_127;
  wire popcount47_i2df_core_128;
  wire popcount47_i2df_core_129;
  wire popcount47_i2df_core_130;
  wire popcount47_i2df_core_131;
  wire popcount47_i2df_core_132;
  wire popcount47_i2df_core_133;
  wire popcount47_i2df_core_134;
  wire popcount47_i2df_core_137;
  wire popcount47_i2df_core_138;
  wire popcount47_i2df_core_139;
  wire popcount47_i2df_core_140;
  wire popcount47_i2df_core_142;
  wire popcount47_i2df_core_143;
  wire popcount47_i2df_core_144;
  wire popcount47_i2df_core_145;
  wire popcount47_i2df_core_146;
  wire popcount47_i2df_core_148;
  wire popcount47_i2df_core_149;
  wire popcount47_i2df_core_152;
  wire popcount47_i2df_core_153;
  wire popcount47_i2df_core_155;
  wire popcount47_i2df_core_156;
  wire popcount47_i2df_core_157;
  wire popcount47_i2df_core_158;
  wire popcount47_i2df_core_159;
  wire popcount47_i2df_core_160;
  wire popcount47_i2df_core_161;
  wire popcount47_i2df_core_162;
  wire popcount47_i2df_core_163;
  wire popcount47_i2df_core_164;
  wire popcount47_i2df_core_165;
  wire popcount47_i2df_core_166;
  wire popcount47_i2df_core_167;
  wire popcount47_i2df_core_168;
  wire popcount47_i2df_core_170;
  wire popcount47_i2df_core_171;
  wire popcount47_i2df_core_173;
  wire popcount47_i2df_core_175;
  wire popcount47_i2df_core_176;
  wire popcount47_i2df_core_179;
  wire popcount47_i2df_core_180;
  wire popcount47_i2df_core_181;
  wire popcount47_i2df_core_184_not;
  wire popcount47_i2df_core_187;
  wire popcount47_i2df_core_188;
  wire popcount47_i2df_core_189;
  wire popcount47_i2df_core_190;
  wire popcount47_i2df_core_191;
  wire popcount47_i2df_core_192;
  wire popcount47_i2df_core_193;
  wire popcount47_i2df_core_194;
  wire popcount47_i2df_core_195;
  wire popcount47_i2df_core_196;
  wire popcount47_i2df_core_197;
  wire popcount47_i2df_core_198;
  wire popcount47_i2df_core_199;
  wire popcount47_i2df_core_200;
  wire popcount47_i2df_core_201;
  wire popcount47_i2df_core_202;
  wire popcount47_i2df_core_203;
  wire popcount47_i2df_core_204;
  wire popcount47_i2df_core_205;
  wire popcount47_i2df_core_206;
  wire popcount47_i2df_core_207;
  wire popcount47_i2df_core_208;
  wire popcount47_i2df_core_209;
  wire popcount47_i2df_core_210;
  wire popcount47_i2df_core_211;
  wire popcount47_i2df_core_212;
  wire popcount47_i2df_core_213;
  wire popcount47_i2df_core_214;
  wire popcount47_i2df_core_215;
  wire popcount47_i2df_core_216;
  wire popcount47_i2df_core_217;
  wire popcount47_i2df_core_218;
  wire popcount47_i2df_core_219;
  wire popcount47_i2df_core_220;
  wire popcount47_i2df_core_221;
  wire popcount47_i2df_core_222;
  wire popcount47_i2df_core_223;
  wire popcount47_i2df_core_224;
  wire popcount47_i2df_core_225;
  wire popcount47_i2df_core_226;
  wire popcount47_i2df_core_227;
  wire popcount47_i2df_core_228;
  wire popcount47_i2df_core_229;
  wire popcount47_i2df_core_230;
  wire popcount47_i2df_core_231;
  wire popcount47_i2df_core_232;
  wire popcount47_i2df_core_235;
  wire popcount47_i2df_core_237;
  wire popcount47_i2df_core_238;
  wire popcount47_i2df_core_239;
  wire popcount47_i2df_core_240;
  wire popcount47_i2df_core_242;
  wire popcount47_i2df_core_244_not;
  wire popcount47_i2df_core_246;
  wire popcount47_i2df_core_249;
  wire popcount47_i2df_core_250;
  wire popcount47_i2df_core_251;
  wire popcount47_i2df_core_252;
  wire popcount47_i2df_core_253;
  wire popcount47_i2df_core_256;
  wire popcount47_i2df_core_257;
  wire popcount47_i2df_core_259;
  wire popcount47_i2df_core_260;
  wire popcount47_i2df_core_262;
  wire popcount47_i2df_core_263;
  wire popcount47_i2df_core_264;
  wire popcount47_i2df_core_265;
  wire popcount47_i2df_core_266;
  wire popcount47_i2df_core_267;
  wire popcount47_i2df_core_268;
  wire popcount47_i2df_core_270;
  wire popcount47_i2df_core_278_not;
  wire popcount47_i2df_core_279;
  wire popcount47_i2df_core_283;
  wire popcount47_i2df_core_284;
  wire popcount47_i2df_core_285;
  wire popcount47_i2df_core_286;
  wire popcount47_i2df_core_287;
  wire popcount47_i2df_core_290;
  wire popcount47_i2df_core_291;
  wire popcount47_i2df_core_292;
  wire popcount47_i2df_core_293;
  wire popcount47_i2df_core_294;
  wire popcount47_i2df_core_296;
  wire popcount47_i2df_core_298;
  wire popcount47_i2df_core_299;
  wire popcount47_i2df_core_302_not;
  wire popcount47_i2df_core_304_not;
  wire popcount47_i2df_core_306;
  wire popcount47_i2df_core_309;
  wire popcount47_i2df_core_310;
  wire popcount47_i2df_core_316;
  wire popcount47_i2df_core_317;
  wire popcount47_i2df_core_321;
  wire popcount47_i2df_core_322;
  wire popcount47_i2df_core_324;
  wire popcount47_i2df_core_326;
  wire popcount47_i2df_core_327;
  wire popcount47_i2df_core_331;
  wire popcount47_i2df_core_332;
  wire popcount47_i2df_core_333;
  wire popcount47_i2df_core_334;
  wire popcount47_i2df_core_336;
  wire popcount47_i2df_core_337;
  wire popcount47_i2df_core_344;
  wire popcount47_i2df_core_346;
  wire popcount47_i2df_core_347;
  wire popcount47_i2df_core_348;
  wire popcount47_i2df_core_349;
  wire popcount47_i2df_core_350;
  wire popcount47_i2df_core_351;
  wire popcount47_i2df_core_352;
  wire popcount47_i2df_core_353;
  wire popcount47_i2df_core_354;
  wire popcount47_i2df_core_355;
  wire popcount47_i2df_core_356;
  wire popcount47_i2df_core_357;
  wire popcount47_i2df_core_358;
  wire popcount47_i2df_core_359;
  wire popcount47_i2df_core_360;
  wire popcount47_i2df_core_361;
  wire popcount47_i2df_core_362;
  wire popcount47_i2df_core_365;
  wire popcount47_i2df_core_366;
  wire popcount47_i2df_core_368;
  wire popcount47_i2df_core_369;
  wire popcount47_i2df_core_370;
  wire popcount47_i2df_core_371;
  wire popcount47_i2df_core_372;

  assign popcount47_i2df_core_049 = input_a[0] ^ input_a[1];
  assign popcount47_i2df_core_050 = input_a[0] & input_a[1];
  assign popcount47_i2df_core_051 = input_a[3] ^ input_a[4];
  assign popcount47_i2df_core_052 = input_a[3] & input_a[4];
  assign popcount47_i2df_core_054 = input_a[2] & input_a[14];
  assign popcount47_i2df_core_056 = popcount47_i2df_core_052 & popcount47_i2df_core_054;
  assign popcount47_i2df_core_057_not = ~input_a[29];
  assign popcount47_i2df_core_062 = input_a[22] & input_a[42];
  assign popcount47_i2df_core_064 = popcount47_i2df_core_056 ^ popcount47_i2df_core_062;
  assign popcount47_i2df_core_065 = popcount47_i2df_core_056 & popcount47_i2df_core_062;
  assign popcount47_i2df_core_068 = input_a[5] ^ input_a[6];
  assign popcount47_i2df_core_069 = input_a[5] & input_a[6];
  assign popcount47_i2df_core_073 = input_a[9] & input_a[31];
  assign popcount47_i2df_core_079 = popcount47_i2df_core_068 & input_a[8];
  assign popcount47_i2df_core_080_not = ~popcount47_i2df_core_073;
  assign popcount47_i2df_core_081 = input_a[29] & popcount47_i2df_core_073;
  assign popcount47_i2df_core_082 = popcount47_i2df_core_080_not ^ input_a[26];
  assign popcount47_i2df_core_083 = popcount47_i2df_core_080_not & popcount47_i2df_core_079;
  assign popcount47_i2df_core_090 = ~(popcount47_i2df_core_057_not | input_a[1]);
  assign popcount47_i2df_core_091 = popcount47_i2df_core_057_not & input_a[5];
  assign popcount47_i2df_core_092 = input_a[26] ^ popcount47_i2df_core_082;
  assign popcount47_i2df_core_094 = input_a[9] ^ popcount47_i2df_core_091;
  assign popcount47_i2df_core_095 = popcount47_i2df_core_092 & popcount47_i2df_core_091;
  assign popcount47_i2df_core_096 = input_a[42] | popcount47_i2df_core_095;
  assign popcount47_i2df_core_099 = popcount47_i2df_core_064 ^ popcount47_i2df_core_096;
  assign popcount47_i2df_core_100 = popcount47_i2df_core_064 & popcount47_i2df_core_096;
  assign popcount47_i2df_core_101 = input_a[44] | popcount47_i2df_core_100;
  assign popcount47_i2df_core_104 = popcount47_i2df_core_065 ^ popcount47_i2df_core_101;
  assign popcount47_i2df_core_105 = popcount47_i2df_core_065 & popcount47_i2df_core_101;
  assign popcount47_i2df_core_107 = input_a[21] ^ input_a[13];
  assign popcount47_i2df_core_108 = input_a[12] & input_a[13];
  assign popcount47_i2df_core_109 = input_a[11] ^ popcount47_i2df_core_107;
  assign popcount47_i2df_core_110 = input_a[11] & popcount47_i2df_core_107;
  assign popcount47_i2df_core_111 = popcount47_i2df_core_108 ^ popcount47_i2df_core_110;
  assign popcount47_i2df_core_112 = popcount47_i2df_core_108 & popcount47_i2df_core_110;
  assign popcount47_i2df_core_113 = input_a[15] ^ input_a[16];
  assign popcount47_i2df_core_114 = input_a[33] & input_a[16];
  assign popcount47_i2df_core_115 = input_a[14] ^ popcount47_i2df_core_113;
  assign popcount47_i2df_core_116 = input_a[14] & popcount47_i2df_core_113;
  assign popcount47_i2df_core_117 = popcount47_i2df_core_114 ^ popcount47_i2df_core_116;
  assign popcount47_i2df_core_118 = popcount47_i2df_core_114 & popcount47_i2df_core_116;
  assign popcount47_i2df_core_119 = popcount47_i2df_core_109 & popcount47_i2df_core_115;
  assign popcount47_i2df_core_120 = popcount47_i2df_core_109 & popcount47_i2df_core_115;
  assign popcount47_i2df_core_121 = input_a[7] ^ popcount47_i2df_core_117;
  assign popcount47_i2df_core_122 = popcount47_i2df_core_111 & popcount47_i2df_core_117;
  assign popcount47_i2df_core_123 = popcount47_i2df_core_121 ^ popcount47_i2df_core_120;
  assign popcount47_i2df_core_124 = popcount47_i2df_core_121 & popcount47_i2df_core_120;
  assign popcount47_i2df_core_125 = popcount47_i2df_core_122 | popcount47_i2df_core_124;
  assign popcount47_i2df_core_126 = input_a[36] ^ popcount47_i2df_core_118;
  assign popcount47_i2df_core_127 = popcount47_i2df_core_112 & input_a[36];
  assign popcount47_i2df_core_128 = popcount47_i2df_core_126 & popcount47_i2df_core_125;
  assign popcount47_i2df_core_129 = popcount47_i2df_core_126 & popcount47_i2df_core_125;
  assign popcount47_i2df_core_130 = popcount47_i2df_core_127 | popcount47_i2df_core_129;
  assign popcount47_i2df_core_131 = input_a[18] ^ input_a[38];
  assign popcount47_i2df_core_132 = input_a[18] & input_a[19];
  assign popcount47_i2df_core_133 = input_a[17] ^ popcount47_i2df_core_131;
  assign popcount47_i2df_core_134 = input_a[17] & popcount47_i2df_core_131;
  assign popcount47_i2df_core_137 = input_a[21] ^ input_a[22];
  assign popcount47_i2df_core_138 = input_a[21] & input_a[22];
  assign popcount47_i2df_core_139 = input_a[20] ^ popcount47_i2df_core_137;
  assign popcount47_i2df_core_140 = input_a[20] & popcount47_i2df_core_137;
  assign popcount47_i2df_core_142 = popcount47_i2df_core_138 & input_a[29];
  assign popcount47_i2df_core_143 = popcount47_i2df_core_133 ^ popcount47_i2df_core_139;
  assign popcount47_i2df_core_144 = ~(popcount47_i2df_core_133 & popcount47_i2df_core_139);
  assign popcount47_i2df_core_145 = popcount47_i2df_core_132 ^ popcount47_i2df_core_138;
  assign popcount47_i2df_core_146 = popcount47_i2df_core_132 & popcount47_i2df_core_138;
  assign popcount47_i2df_core_148 = input_a[31] & popcount47_i2df_core_144;
  assign popcount47_i2df_core_149 = popcount47_i2df_core_146 | popcount47_i2df_core_148;
  assign popcount47_i2df_core_152 = input_a[46] ^ popcount47_i2df_core_149;
  assign popcount47_i2df_core_153 = popcount47_i2df_core_142 & popcount47_i2df_core_149;
  assign popcount47_i2df_core_155 = popcount47_i2df_core_119 ^ popcount47_i2df_core_143;
  assign popcount47_i2df_core_156 = ~popcount47_i2df_core_119;
  assign popcount47_i2df_core_157 = input_a[30] ^ input_a[32];
  assign popcount47_i2df_core_158 = popcount47_i2df_core_123 & popcount47_i2df_core_145;
  assign popcount47_i2df_core_159 = popcount47_i2df_core_157 ^ input_a[35];
  assign popcount47_i2df_core_160 = popcount47_i2df_core_157 & popcount47_i2df_core_156;
  assign popcount47_i2df_core_161 = popcount47_i2df_core_158 | popcount47_i2df_core_160;
  assign popcount47_i2df_core_162 = popcount47_i2df_core_128 ^ popcount47_i2df_core_152;
  assign popcount47_i2df_core_163 = popcount47_i2df_core_128 & input_a[40];
  assign popcount47_i2df_core_164 = popcount47_i2df_core_162 ^ popcount47_i2df_core_161;
  assign popcount47_i2df_core_165 = popcount47_i2df_core_162 & popcount47_i2df_core_161;
  assign popcount47_i2df_core_166 = popcount47_i2df_core_163 | input_a[4];
  assign popcount47_i2df_core_167 = popcount47_i2df_core_130 ^ popcount47_i2df_core_153;
  assign popcount47_i2df_core_168 = popcount47_i2df_core_130 & popcount47_i2df_core_153;
  assign popcount47_i2df_core_170 = popcount47_i2df_core_167 & popcount47_i2df_core_166;
  assign popcount47_i2df_core_171 = popcount47_i2df_core_168 | popcount47_i2df_core_170;
  assign popcount47_i2df_core_173 = popcount47_i2df_core_090 & input_a[34];
  assign popcount47_i2df_core_175 = popcount47_i2df_core_094 & popcount47_i2df_core_159;
  assign popcount47_i2df_core_176 = input_a[3] ^ popcount47_i2df_core_173;
  assign popcount47_i2df_core_179 = popcount47_i2df_core_099 ^ input_a[21];
  assign popcount47_i2df_core_180 = popcount47_i2df_core_099 & input_a[38];
  assign popcount47_i2df_core_181 = input_a[12] ^ popcount47_i2df_core_175;
  assign popcount47_i2df_core_184_not = ~popcount47_i2df_core_104;
  assign popcount47_i2df_core_187 = popcount47_i2df_core_184_not & input_a[1];
  assign popcount47_i2df_core_188 = popcount47_i2df_core_104 & popcount47_i2df_core_187;
  assign popcount47_i2df_core_189 = popcount47_i2df_core_105 ^ popcount47_i2df_core_171;
  assign popcount47_i2df_core_190 = popcount47_i2df_core_105 & popcount47_i2df_core_171;
  assign popcount47_i2df_core_191 = popcount47_i2df_core_189 ^ popcount47_i2df_core_188;
  assign popcount47_i2df_core_192 = popcount47_i2df_core_189 & popcount47_i2df_core_188;
  assign popcount47_i2df_core_193 = popcount47_i2df_core_190 | popcount47_i2df_core_192;
  assign popcount47_i2df_core_194 = input_a[24] ^ input_a[25];
  assign popcount47_i2df_core_195 = input_a[24] & input_a[43];
  assign popcount47_i2df_core_196 = input_a[23] ^ popcount47_i2df_core_194;
  assign popcount47_i2df_core_197 = input_a[23] & popcount47_i2df_core_194;
  assign popcount47_i2df_core_198 = ~(popcount47_i2df_core_195 | popcount47_i2df_core_197);
  assign popcount47_i2df_core_199 = popcount47_i2df_core_195 & popcount47_i2df_core_197;
  assign popcount47_i2df_core_200 = input_a[26] | input_a[28];
  assign popcount47_i2df_core_201 = input_a[27] & input_a[28];
  assign popcount47_i2df_core_202 = input_a[26] ^ popcount47_i2df_core_200;
  assign popcount47_i2df_core_203 = input_a[26] & popcount47_i2df_core_200;
  assign popcount47_i2df_core_204 = popcount47_i2df_core_201 ^ popcount47_i2df_core_203;
  assign popcount47_i2df_core_205 = popcount47_i2df_core_201 & popcount47_i2df_core_203;
  assign popcount47_i2df_core_206 = input_a[16] ^ popcount47_i2df_core_202;
  assign popcount47_i2df_core_207 = popcount47_i2df_core_196 & popcount47_i2df_core_202;
  assign popcount47_i2df_core_208 = popcount47_i2df_core_198 ^ popcount47_i2df_core_204;
  assign popcount47_i2df_core_209 = popcount47_i2df_core_198 & popcount47_i2df_core_204;
  assign popcount47_i2df_core_210 = popcount47_i2df_core_208 ^ popcount47_i2df_core_207;
  assign popcount47_i2df_core_211 = popcount47_i2df_core_208 & popcount47_i2df_core_207;
  assign popcount47_i2df_core_212 = popcount47_i2df_core_209 | popcount47_i2df_core_211;
  assign popcount47_i2df_core_213 = popcount47_i2df_core_199 & popcount47_i2df_core_205;
  assign popcount47_i2df_core_214 = popcount47_i2df_core_199 & popcount47_i2df_core_205;
  assign popcount47_i2df_core_215 = popcount47_i2df_core_213 ^ popcount47_i2df_core_212;
  assign popcount47_i2df_core_216 = popcount47_i2df_core_213 & popcount47_i2df_core_212;
  assign popcount47_i2df_core_217 = popcount47_i2df_core_214 | popcount47_i2df_core_216;
  assign popcount47_i2df_core_218 = ~input_a[30];
  assign popcount47_i2df_core_219 = input_a[30] & input_a[31];
  assign popcount47_i2df_core_220 = input_a[29] ^ popcount47_i2df_core_218;
  assign popcount47_i2df_core_221 = input_a[29] & popcount47_i2df_core_218;
  assign popcount47_i2df_core_222 = popcount47_i2df_core_219 ^ popcount47_i2df_core_221;
  assign popcount47_i2df_core_223 = popcount47_i2df_core_219 & popcount47_i2df_core_221;
  assign popcount47_i2df_core_224 = ~(input_a[33] | input_a[34]);
  assign popcount47_i2df_core_225 = input_a[33] & input_a[34];
  assign popcount47_i2df_core_226 = input_a[24] ^ popcount47_i2df_core_224;
  assign popcount47_i2df_core_227 = input_a[32] & popcount47_i2df_core_224;
  assign popcount47_i2df_core_228 = popcount47_i2df_core_225 ^ popcount47_i2df_core_227;
  assign popcount47_i2df_core_229 = popcount47_i2df_core_225 & popcount47_i2df_core_227;
  assign popcount47_i2df_core_230 = popcount47_i2df_core_220 & input_a[11];
  assign popcount47_i2df_core_231 = popcount47_i2df_core_220 & popcount47_i2df_core_226;
  assign popcount47_i2df_core_232 = popcount47_i2df_core_222 ^ popcount47_i2df_core_228;
  assign popcount47_i2df_core_235 = popcount47_i2df_core_232 & popcount47_i2df_core_231;
  assign popcount47_i2df_core_237 = popcount47_i2df_core_223 ^ input_a[25];
  assign popcount47_i2df_core_238 = popcount47_i2df_core_223 & popcount47_i2df_core_229;
  assign popcount47_i2df_core_239 = popcount47_i2df_core_237 ^ popcount47_i2df_core_235;
  assign popcount47_i2df_core_240 = popcount47_i2df_core_237 & popcount47_i2df_core_235;
  assign popcount47_i2df_core_242 = popcount47_i2df_core_206 ^ popcount47_i2df_core_230;
  assign popcount47_i2df_core_244_not = ~popcount47_i2df_core_210;
  assign popcount47_i2df_core_246 = ~(popcount47_i2df_core_244_not & input_a[42]);
  assign popcount47_i2df_core_249 = ~popcount47_i2df_core_215;
  assign popcount47_i2df_core_250 = popcount47_i2df_core_215 & popcount47_i2df_core_239;
  assign popcount47_i2df_core_251 = popcount47_i2df_core_249 ^ popcount47_i2df_core_210;
  assign popcount47_i2df_core_252 = ~(popcount47_i2df_core_249 & popcount47_i2df_core_210);
  assign popcount47_i2df_core_253 = ~(popcount47_i2df_core_250 | popcount47_i2df_core_252);
  assign popcount47_i2df_core_256 = popcount47_i2df_core_217 ^ popcount47_i2df_core_253;
  assign popcount47_i2df_core_257 = popcount47_i2df_core_217 & input_a[11];
  assign popcount47_i2df_core_259 = input_a[36] ^ input_a[37];
  assign popcount47_i2df_core_260 = input_a[36] & input_a[37];
  assign popcount47_i2df_core_262 = input_a[35] & popcount47_i2df_core_259;
  assign popcount47_i2df_core_263 = popcount47_i2df_core_260 ^ popcount47_i2df_core_262;
  assign popcount47_i2df_core_264 = popcount47_i2df_core_260 & popcount47_i2df_core_262;
  assign popcount47_i2df_core_265 = input_a[39] ^ input_a[40];
  assign popcount47_i2df_core_266 = input_a[39] & input_a[40];
  assign popcount47_i2df_core_267 = input_a[38] ^ popcount47_i2df_core_265;
  assign popcount47_i2df_core_268 = input_a[38] & popcount47_i2df_core_265;
  assign popcount47_i2df_core_270 = popcount47_i2df_core_266 & popcount47_i2df_core_268;
  assign popcount47_i2df_core_278_not = ~input_a[5];
  assign popcount47_i2df_core_279 = popcount47_i2df_core_264 & popcount47_i2df_core_270;
  assign popcount47_i2df_core_283 = input_a[42] ^ input_a[43];
  assign popcount47_i2df_core_284 = input_a[42] & input_a[43];
  assign popcount47_i2df_core_285 = input_a[41] ^ popcount47_i2df_core_283;
  assign popcount47_i2df_core_286 = input_a[41] & popcount47_i2df_core_283;
  assign popcount47_i2df_core_287 = popcount47_i2df_core_284 ^ input_a[18];
  assign popcount47_i2df_core_290 = ~(input_a[45] & input_a[46]);
  assign popcount47_i2df_core_291 = input_a[44] ^ input_a[45];
  assign popcount47_i2df_core_292 = input_a[44] & input_a[45];
  assign popcount47_i2df_core_293 = popcount47_i2df_core_290 ^ popcount47_i2df_core_292;
  assign popcount47_i2df_core_294 = popcount47_i2df_core_290 & popcount47_i2df_core_292;
  assign popcount47_i2df_core_296 = popcount47_i2df_core_285 & popcount47_i2df_core_291;
  assign popcount47_i2df_core_298 = popcount47_i2df_core_287 & popcount47_i2df_core_293;
  assign popcount47_i2df_core_299 = input_a[35] ^ popcount47_i2df_core_296;
  assign popcount47_i2df_core_302_not = ~popcount47_i2df_core_294;
  assign popcount47_i2df_core_304_not = ~popcount47_i2df_core_302_not;
  assign popcount47_i2df_core_306 = popcount47_i2df_core_294 | popcount47_i2df_core_302_not;
  assign popcount47_i2df_core_309 = input_a[15] & input_a[32];
  assign popcount47_i2df_core_310 = popcount47_i2df_core_263 & popcount47_i2df_core_299;
  assign popcount47_i2df_core_316 = popcount47_i2df_core_304_not ^ input_a[21];
  assign popcount47_i2df_core_317 = popcount47_i2df_core_304_not & input_a[21];
  assign popcount47_i2df_core_321 = popcount47_i2df_core_306 ^ input_a[19];
  assign popcount47_i2df_core_322 = popcount47_i2df_core_306 & popcount47_i2df_core_317;
  assign popcount47_i2df_core_324 = popcount47_i2df_core_242 ^ input_a[33];
  assign popcount47_i2df_core_326 = popcount47_i2df_core_246 ^ popcount47_i2df_core_309;
  assign popcount47_i2df_core_327 = popcount47_i2df_core_246 & popcount47_i2df_core_309;
  assign popcount47_i2df_core_331 = popcount47_i2df_core_251 ^ popcount47_i2df_core_316;
  assign popcount47_i2df_core_332 = ~popcount47_i2df_core_251;
  assign popcount47_i2df_core_333 = input_a[3] ^ popcount47_i2df_core_327;
  assign popcount47_i2df_core_334 = popcount47_i2df_core_331 & popcount47_i2df_core_327;
  assign popcount47_i2df_core_336 = popcount47_i2df_core_256 ^ popcount47_i2df_core_321;
  assign popcount47_i2df_core_337 = popcount47_i2df_core_256 & popcount47_i2df_core_321;
  assign popcount47_i2df_core_344 = popcount47_i2df_core_257 & input_a[25];
  assign popcount47_i2df_core_346 = popcount47_i2df_core_090 ^ popcount47_i2df_core_324;
  assign popcount47_i2df_core_347 = popcount47_i2df_core_090 & popcount47_i2df_core_324;
  assign popcount47_i2df_core_348 = popcount47_i2df_core_176 ^ popcount47_i2df_core_326;
  assign popcount47_i2df_core_349 = popcount47_i2df_core_176 & popcount47_i2df_core_326;
  assign popcount47_i2df_core_350 = popcount47_i2df_core_348 ^ popcount47_i2df_core_347;
  assign popcount47_i2df_core_351 = popcount47_i2df_core_348 & popcount47_i2df_core_347;
  assign popcount47_i2df_core_352 = input_a[32] | popcount47_i2df_core_351;
  assign popcount47_i2df_core_353 = popcount47_i2df_core_181 ^ popcount47_i2df_core_333;
  assign popcount47_i2df_core_354 = popcount47_i2df_core_181 & popcount47_i2df_core_333;
  assign popcount47_i2df_core_355 = popcount47_i2df_core_353 ^ popcount47_i2df_core_352;
  assign popcount47_i2df_core_356 = popcount47_i2df_core_353 & popcount47_i2df_core_352;
  assign popcount47_i2df_core_357 = popcount47_i2df_core_354 | popcount47_i2df_core_356;
  assign popcount47_i2df_core_358 = input_a[10] ^ popcount47_i2df_core_336;
  assign popcount47_i2df_core_359 = input_a[10] & popcount47_i2df_core_336;
  assign popcount47_i2df_core_360 = popcount47_i2df_core_358 ^ popcount47_i2df_core_357;
  assign popcount47_i2df_core_361 = popcount47_i2df_core_358 & popcount47_i2df_core_357;
  assign popcount47_i2df_core_362 = popcount47_i2df_core_359 | popcount47_i2df_core_361;
  assign popcount47_i2df_core_365 = popcount47_i2df_core_191 ^ popcount47_i2df_core_362;
  assign popcount47_i2df_core_366 = popcount47_i2df_core_191 & popcount47_i2df_core_362;
  assign popcount47_i2df_core_368 = popcount47_i2df_core_193 ^ popcount47_i2df_core_344;
  assign popcount47_i2df_core_369 = popcount47_i2df_core_193 & popcount47_i2df_core_344;
  assign popcount47_i2df_core_370 = popcount47_i2df_core_368 ^ popcount47_i2df_core_366;
  assign popcount47_i2df_core_371 = popcount47_i2df_core_368 & popcount47_i2df_core_366;
  assign popcount47_i2df_core_372 = popcount47_i2df_core_369 | popcount47_i2df_core_371;

  assign popcount47_i2df_out[0] = popcount47_i2df_core_346;
  assign popcount47_i2df_out[1] = 1'b1;
  assign popcount47_i2df_out[2] = popcount47_i2df_core_355;
  assign popcount47_i2df_out[3] = popcount47_i2df_core_360;
  assign popcount47_i2df_out[4] = popcount47_i2df_core_365;
  assign popcount47_i2df_out[5] = popcount47_i2df_core_370;
endmodule