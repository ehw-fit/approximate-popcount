// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.65305
// WCE=19.0
// EP=0.881976%
// Printed PDK parameters:
//  Area=4830570.0
//  Delay=15688585.0
//  Power=251410.0

module popcount38_h9vn(input [37:0] input_a, output [5:0] popcount38_h9vn_out);
  wire popcount38_h9vn_core_040;
  wire popcount38_h9vn_core_042;
  wire popcount38_h9vn_core_043;
  wire popcount38_h9vn_core_044;
  wire popcount38_h9vn_core_046;
  wire popcount38_h9vn_core_050;
  wire popcount38_h9vn_core_054;
  wire popcount38_h9vn_core_055;
  wire popcount38_h9vn_core_057;
  wire popcount38_h9vn_core_058;
  wire popcount38_h9vn_core_059;
  wire popcount38_h9vn_core_062;
  wire popcount38_h9vn_core_064;
  wire popcount38_h9vn_core_065;
  wire popcount38_h9vn_core_066;
  wire popcount38_h9vn_core_068;
  wire popcount38_h9vn_core_069;
  wire popcount38_h9vn_core_070;
  wire popcount38_h9vn_core_071;
  wire popcount38_h9vn_core_072;
  wire popcount38_h9vn_core_073;
  wire popcount38_h9vn_core_074;
  wire popcount38_h9vn_core_075;
  wire popcount38_h9vn_core_077;
  wire popcount38_h9vn_core_078;
  wire popcount38_h9vn_core_079;
  wire popcount38_h9vn_core_080;
  wire popcount38_h9vn_core_083;
  wire popcount38_h9vn_core_084;
  wire popcount38_h9vn_core_085;
  wire popcount38_h9vn_core_086;
  wire popcount38_h9vn_core_087;
  wire popcount38_h9vn_core_088;
  wire popcount38_h9vn_core_089;
  wire popcount38_h9vn_core_091;
  wire popcount38_h9vn_core_093;
  wire popcount38_h9vn_core_097;
  wire popcount38_h9vn_core_099;
  wire popcount38_h9vn_core_100;
  wire popcount38_h9vn_core_101;
  wire popcount38_h9vn_core_103;
  wire popcount38_h9vn_core_104;
  wire popcount38_h9vn_core_105;
  wire popcount38_h9vn_core_106;
  wire popcount38_h9vn_core_107;
  wire popcount38_h9vn_core_108;
  wire popcount38_h9vn_core_110;
  wire popcount38_h9vn_core_111;
  wire popcount38_h9vn_core_112;
  wire popcount38_h9vn_core_113;
  wire popcount38_h9vn_core_114;
  wire popcount38_h9vn_core_115;
  wire popcount38_h9vn_core_120;
  wire popcount38_h9vn_core_121;
  wire popcount38_h9vn_core_122;
  wire popcount38_h9vn_core_124;
  wire popcount38_h9vn_core_125;
  wire popcount38_h9vn_core_126;
  wire popcount38_h9vn_core_127;
  wire popcount38_h9vn_core_128;
  wire popcount38_h9vn_core_130;
  wire popcount38_h9vn_core_132;
  wire popcount38_h9vn_core_133;
  wire popcount38_h9vn_core_134;
  wire popcount38_h9vn_core_135;
  wire popcount38_h9vn_core_136;
  wire popcount38_h9vn_core_137;
  wire popcount38_h9vn_core_138;
  wire popcount38_h9vn_core_139;
  wire popcount38_h9vn_core_140;
  wire popcount38_h9vn_core_141;
  wire popcount38_h9vn_core_143;
  wire popcount38_h9vn_core_144;
  wire popcount38_h9vn_core_146;
  wire popcount38_h9vn_core_150;
  wire popcount38_h9vn_core_154;
  wire popcount38_h9vn_core_155;
  wire popcount38_h9vn_core_156;
  wire popcount38_h9vn_core_157;
  wire popcount38_h9vn_core_158;
  wire popcount38_h9vn_core_159;
  wire popcount38_h9vn_core_162;
  wire popcount38_h9vn_core_165;
  wire popcount38_h9vn_core_166;
  wire popcount38_h9vn_core_167;
  wire popcount38_h9vn_core_169;
  wire popcount38_h9vn_core_170;
  wire popcount38_h9vn_core_172;
  wire popcount38_h9vn_core_174;
  wire popcount38_h9vn_core_178;
  wire popcount38_h9vn_core_180;
  wire popcount38_h9vn_core_181;
  wire popcount38_h9vn_core_183;
  wire popcount38_h9vn_core_184;
  wire popcount38_h9vn_core_187;
  wire popcount38_h9vn_core_188;
  wire popcount38_h9vn_core_190;
  wire popcount38_h9vn_core_191;
  wire popcount38_h9vn_core_194;
  wire popcount38_h9vn_core_195;
  wire popcount38_h9vn_core_196;
  wire popcount38_h9vn_core_197;
  wire popcount38_h9vn_core_198;
  wire popcount38_h9vn_core_200;
  wire popcount38_h9vn_core_201;
  wire popcount38_h9vn_core_202;
  wire popcount38_h9vn_core_203;
  wire popcount38_h9vn_core_205;
  wire popcount38_h9vn_core_206;
  wire popcount38_h9vn_core_207;
  wire popcount38_h9vn_core_208;
  wire popcount38_h9vn_core_209;
  wire popcount38_h9vn_core_211;
  wire popcount38_h9vn_core_212;
  wire popcount38_h9vn_core_218;
  wire popcount38_h9vn_core_219;
  wire popcount38_h9vn_core_220;
  wire popcount38_h9vn_core_221;
  wire popcount38_h9vn_core_224;
  wire popcount38_h9vn_core_225;
  wire popcount38_h9vn_core_226;
  wire popcount38_h9vn_core_227;
  wire popcount38_h9vn_core_228;
  wire popcount38_h9vn_core_229;
  wire popcount38_h9vn_core_231;
  wire popcount38_h9vn_core_232;
  wire popcount38_h9vn_core_233;
  wire popcount38_h9vn_core_235;
  wire popcount38_h9vn_core_237;
  wire popcount38_h9vn_core_238;
  wire popcount38_h9vn_core_240;
  wire popcount38_h9vn_core_241;
  wire popcount38_h9vn_core_242;
  wire popcount38_h9vn_core_243;
  wire popcount38_h9vn_core_244;
  wire popcount38_h9vn_core_245;
  wire popcount38_h9vn_core_248;
  wire popcount38_h9vn_core_249;
  wire popcount38_h9vn_core_251;
  wire popcount38_h9vn_core_252;
  wire popcount38_h9vn_core_254;
  wire popcount38_h9vn_core_255;
  wire popcount38_h9vn_core_256;
  wire popcount38_h9vn_core_257;
  wire popcount38_h9vn_core_258;
  wire popcount38_h9vn_core_259;
  wire popcount38_h9vn_core_260_not;
  wire popcount38_h9vn_core_261;
  wire popcount38_h9vn_core_262;
  wire popcount38_h9vn_core_263;
  wire popcount38_h9vn_core_265;
  wire popcount38_h9vn_core_266;
  wire popcount38_h9vn_core_270;
  wire popcount38_h9vn_core_273;
  wire popcount38_h9vn_core_274;
  wire popcount38_h9vn_core_275;
  wire popcount38_h9vn_core_279;
  wire popcount38_h9vn_core_280;
  wire popcount38_h9vn_core_282_not;
  wire popcount38_h9vn_core_284;
  wire popcount38_h9vn_core_289;
  wire popcount38_h9vn_core_290;
  wire popcount38_h9vn_core_292;
  wire popcount38_h9vn_core_293_not;
  wire popcount38_h9vn_core_295;
  wire popcount38_h9vn_core_296;

  assign popcount38_h9vn_core_040 = ~(input_a[32] | input_a[25]);
  assign popcount38_h9vn_core_042 = input_a[37] ^ input_a[33];
  assign popcount38_h9vn_core_043 = input_a[0] ^ input_a[11];
  assign popcount38_h9vn_core_044 = ~(input_a[20] ^ input_a[9]);
  assign popcount38_h9vn_core_046 = input_a[4] ^ input_a[9];
  assign popcount38_h9vn_core_050 = input_a[15] ^ input_a[28];
  assign popcount38_h9vn_core_054 = input_a[2] | input_a[6];
  assign popcount38_h9vn_core_055 = ~input_a[31];
  assign popcount38_h9vn_core_057 = input_a[9] ^ input_a[17];
  assign popcount38_h9vn_core_058 = ~(input_a[5] | input_a[23]);
  assign popcount38_h9vn_core_059 = ~(input_a[28] ^ input_a[9]);
  assign popcount38_h9vn_core_062 = ~(input_a[27] | input_a[10]);
  assign popcount38_h9vn_core_064 = ~(input_a[37] & input_a[29]);
  assign popcount38_h9vn_core_065 = input_a[27] ^ input_a[13];
  assign popcount38_h9vn_core_066 = ~(input_a[10] ^ input_a[9]);
  assign popcount38_h9vn_core_068 = ~(input_a[13] ^ input_a[21]);
  assign popcount38_h9vn_core_069 = input_a[32] & input_a[3];
  assign popcount38_h9vn_core_070 = ~(input_a[3] | input_a[11]);
  assign popcount38_h9vn_core_071 = ~(input_a[17] & input_a[21]);
  assign popcount38_h9vn_core_072 = input_a[29] & input_a[25];
  assign popcount38_h9vn_core_073 = input_a[31] ^ input_a[16];
  assign popcount38_h9vn_core_074 = ~input_a[7];
  assign popcount38_h9vn_core_075 = ~(input_a[4] & input_a[27]);
  assign popcount38_h9vn_core_077 = ~(input_a[32] ^ input_a[9]);
  assign popcount38_h9vn_core_078 = ~(input_a[33] | input_a[37]);
  assign popcount38_h9vn_core_079 = input_a[4] ^ input_a[9];
  assign popcount38_h9vn_core_080 = ~(input_a[12] | input_a[2]);
  assign popcount38_h9vn_core_083 = input_a[3] ^ input_a[36];
  assign popcount38_h9vn_core_084 = ~input_a[6];
  assign popcount38_h9vn_core_085 = input_a[33] | input_a[12];
  assign popcount38_h9vn_core_086 = input_a[18] | input_a[19];
  assign popcount38_h9vn_core_087 = ~(input_a[33] | input_a[31]);
  assign popcount38_h9vn_core_088 = ~(input_a[13] & input_a[16]);
  assign popcount38_h9vn_core_089 = ~(input_a[28] | input_a[29]);
  assign popcount38_h9vn_core_091 = input_a[14] ^ input_a[24];
  assign popcount38_h9vn_core_093 = ~(input_a[35] | input_a[7]);
  assign popcount38_h9vn_core_097 = input_a[16] ^ input_a[21];
  assign popcount38_h9vn_core_099 = ~input_a[10];
  assign popcount38_h9vn_core_100 = ~(input_a[6] & input_a[21]);
  assign popcount38_h9vn_core_101 = input_a[30] & input_a[5];
  assign popcount38_h9vn_core_103 = ~(input_a[28] ^ input_a[17]);
  assign popcount38_h9vn_core_104 = input_a[21] & input_a[24];
  assign popcount38_h9vn_core_105 = input_a[12] ^ input_a[29];
  assign popcount38_h9vn_core_106 = input_a[31] | input_a[4];
  assign popcount38_h9vn_core_107 = input_a[16] | input_a[18];
  assign popcount38_h9vn_core_108 = input_a[27] & input_a[33];
  assign popcount38_h9vn_core_110 = input_a[17] | input_a[11];
  assign popcount38_h9vn_core_111 = input_a[7] ^ input_a[37];
  assign popcount38_h9vn_core_112 = input_a[18] ^ input_a[30];
  assign popcount38_h9vn_core_113 = ~(input_a[23] & input_a[22]);
  assign popcount38_h9vn_core_114 = ~input_a[26];
  assign popcount38_h9vn_core_115 = input_a[11] ^ input_a[10];
  assign popcount38_h9vn_core_120 = ~(input_a[32] | input_a[7]);
  assign popcount38_h9vn_core_121 = input_a[20] | input_a[3];
  assign popcount38_h9vn_core_122 = ~(input_a[35] & input_a[24]);
  assign popcount38_h9vn_core_124 = input_a[14] | input_a[11];
  assign popcount38_h9vn_core_125 = ~(input_a[33] & input_a[15]);
  assign popcount38_h9vn_core_126 = ~(input_a[5] & input_a[13]);
  assign popcount38_h9vn_core_127 = ~(input_a[7] | input_a[31]);
  assign popcount38_h9vn_core_128 = input_a[14] ^ input_a[29];
  assign popcount38_h9vn_core_130 = ~(input_a[16] | input_a[1]);
  assign popcount38_h9vn_core_132 = ~(input_a[37] & input_a[9]);
  assign popcount38_h9vn_core_133 = ~(input_a[25] | input_a[15]);
  assign popcount38_h9vn_core_134 = input_a[18] & input_a[35];
  assign popcount38_h9vn_core_135 = ~input_a[31];
  assign popcount38_h9vn_core_136 = input_a[24] | input_a[17];
  assign popcount38_h9vn_core_137 = ~(input_a[34] | input_a[33]);
  assign popcount38_h9vn_core_138 = input_a[27] | input_a[3];
  assign popcount38_h9vn_core_139 = input_a[5] | input_a[5];
  assign popcount38_h9vn_core_140 = ~input_a[26];
  assign popcount38_h9vn_core_141 = ~(input_a[14] | input_a[23]);
  assign popcount38_h9vn_core_143 = ~(input_a[33] ^ input_a[13]);
  assign popcount38_h9vn_core_144 = input_a[24] | input_a[31];
  assign popcount38_h9vn_core_146 = input_a[20] & input_a[34];
  assign popcount38_h9vn_core_150 = input_a[19] & input_a[18];
  assign popcount38_h9vn_core_154 = ~input_a[12];
  assign popcount38_h9vn_core_155 = ~(input_a[31] ^ input_a[5]);
  assign popcount38_h9vn_core_156 = ~(input_a[4] & input_a[6]);
  assign popcount38_h9vn_core_157 = input_a[13] ^ input_a[21];
  assign popcount38_h9vn_core_158 = ~input_a[23];
  assign popcount38_h9vn_core_159 = ~(input_a[28] & input_a[1]);
  assign popcount38_h9vn_core_162 = input_a[16] ^ input_a[35];
  assign popcount38_h9vn_core_165 = ~(input_a[29] & input_a[9]);
  assign popcount38_h9vn_core_166 = ~(input_a[27] ^ input_a[10]);
  assign popcount38_h9vn_core_167 = ~input_a[31];
  assign popcount38_h9vn_core_169 = input_a[2] | input_a[28];
  assign popcount38_h9vn_core_170 = ~(input_a[15] & input_a[21]);
  assign popcount38_h9vn_core_172 = ~(input_a[13] | input_a[3]);
  assign popcount38_h9vn_core_174 = input_a[27] & input_a[20];
  assign popcount38_h9vn_core_178 = input_a[36] & input_a[25];
  assign popcount38_h9vn_core_180 = ~input_a[20];
  assign popcount38_h9vn_core_181 = ~(input_a[7] ^ input_a[30]);
  assign popcount38_h9vn_core_183 = ~(input_a[21] ^ input_a[8]);
  assign popcount38_h9vn_core_184 = ~(input_a[12] ^ input_a[1]);
  assign popcount38_h9vn_core_187 = ~input_a[12];
  assign popcount38_h9vn_core_188 = input_a[8] | input_a[22];
  assign popcount38_h9vn_core_190 = ~input_a[20];
  assign popcount38_h9vn_core_191 = ~(input_a[7] & input_a[25]);
  assign popcount38_h9vn_core_194 = ~input_a[36];
  assign popcount38_h9vn_core_195 = ~input_a[7];
  assign popcount38_h9vn_core_196 = input_a[26] ^ input_a[9];
  assign popcount38_h9vn_core_197 = input_a[9] & input_a[27];
  assign popcount38_h9vn_core_198 = input_a[27] | input_a[11];
  assign popcount38_h9vn_core_200 = input_a[25] ^ input_a[27];
  assign popcount38_h9vn_core_201 = input_a[28] ^ input_a[21];
  assign popcount38_h9vn_core_202 = input_a[8] ^ input_a[30];
  assign popcount38_h9vn_core_203 = ~(input_a[22] | input_a[37]);
  assign popcount38_h9vn_core_205 = input_a[1] ^ input_a[27];
  assign popcount38_h9vn_core_206 = input_a[10] | input_a[13];
  assign popcount38_h9vn_core_207 = ~(input_a[37] & input_a[36]);
  assign popcount38_h9vn_core_208 = input_a[23] ^ input_a[14];
  assign popcount38_h9vn_core_209 = ~(input_a[23] ^ input_a[22]);
  assign popcount38_h9vn_core_211 = input_a[9] | input_a[37];
  assign popcount38_h9vn_core_212 = ~(input_a[16] | input_a[7]);
  assign popcount38_h9vn_core_218 = input_a[30] ^ input_a[10];
  assign popcount38_h9vn_core_219 = input_a[17] ^ input_a[12];
  assign popcount38_h9vn_core_220 = ~(input_a[4] ^ input_a[16]);
  assign popcount38_h9vn_core_221 = input_a[27] ^ input_a[29];
  assign popcount38_h9vn_core_224 = ~input_a[19];
  assign popcount38_h9vn_core_225 = input_a[24] & input_a[23];
  assign popcount38_h9vn_core_226 = ~(input_a[16] ^ input_a[25]);
  assign popcount38_h9vn_core_227 = ~(input_a[19] ^ input_a[22]);
  assign popcount38_h9vn_core_228 = input_a[7] | input_a[23];
  assign popcount38_h9vn_core_229 = input_a[28] & input_a[21];
  assign popcount38_h9vn_core_231 = input_a[17] ^ input_a[35];
  assign popcount38_h9vn_core_232 = ~(input_a[6] | input_a[13]);
  assign popcount38_h9vn_core_233 = input_a[8] ^ input_a[27];
  assign popcount38_h9vn_core_235 = input_a[16] & input_a[37];
  assign popcount38_h9vn_core_237 = input_a[14] | input_a[30];
  assign popcount38_h9vn_core_238 = input_a[0] | input_a[5];
  assign popcount38_h9vn_core_240 = input_a[25] & input_a[7];
  assign popcount38_h9vn_core_241 = ~input_a[25];
  assign popcount38_h9vn_core_242 = input_a[15] | input_a[11];
  assign popcount38_h9vn_core_243 = input_a[26] ^ input_a[30];
  assign popcount38_h9vn_core_244 = input_a[25] & input_a[4];
  assign popcount38_h9vn_core_245 = input_a[10] & input_a[21];
  assign popcount38_h9vn_core_248 = input_a[29] ^ input_a[10];
  assign popcount38_h9vn_core_249 = input_a[20] & input_a[23];
  assign popcount38_h9vn_core_251 = ~(input_a[11] | input_a[28]);
  assign popcount38_h9vn_core_252 = ~input_a[37];
  assign popcount38_h9vn_core_254 = input_a[36] | input_a[9];
  assign popcount38_h9vn_core_255 = ~(input_a[21] & popcount38_h9vn_core_240);
  assign popcount38_h9vn_core_256 = input_a[21] & popcount38_h9vn_core_240;
  assign popcount38_h9vn_core_257 = popcount38_h9vn_core_255 ^ popcount38_h9vn_core_254;
  assign popcount38_h9vn_core_258 = ~(input_a[2] ^ input_a[8]);
  assign popcount38_h9vn_core_259 = popcount38_h9vn_core_256 | input_a[9];
  assign popcount38_h9vn_core_260_not = ~input_a[37];
  assign popcount38_h9vn_core_261 = input_a[27] & input_a[34];
  assign popcount38_h9vn_core_262 = input_a[36] | popcount38_h9vn_core_259;
  assign popcount38_h9vn_core_263 = input_a[31] & input_a[34];
  assign popcount38_h9vn_core_265 = ~(input_a[29] ^ input_a[2]);
  assign popcount38_h9vn_core_266 = input_a[21] ^ input_a[20];
  assign popcount38_h9vn_core_270 = input_a[12] & input_a[5];
  assign popcount38_h9vn_core_273 = ~(input_a[5] ^ input_a[29]);
  assign popcount38_h9vn_core_274 = input_a[34] | input_a[2];
  assign popcount38_h9vn_core_275 = input_a[33] ^ input_a[9];
  assign popcount38_h9vn_core_279 = ~(popcount38_h9vn_core_257 & input_a[0]);
  assign popcount38_h9vn_core_280 = popcount38_h9vn_core_257 & input_a[0];
  assign popcount38_h9vn_core_282_not = ~popcount38_h9vn_core_262;
  assign popcount38_h9vn_core_284 = popcount38_h9vn_core_282_not ^ popcount38_h9vn_core_280;
  assign popcount38_h9vn_core_289 = input_a[0] | popcount38_h9vn_core_262;
  assign popcount38_h9vn_core_290 = ~(input_a[2] & input_a[33]);
  assign popcount38_h9vn_core_292 = input_a[25] ^ input_a[0];
  assign popcount38_h9vn_core_293_not = ~input_a[6];
  assign popcount38_h9vn_core_295 = ~input_a[14];
  assign popcount38_h9vn_core_296 = input_a[0] ^ input_a[29];

  assign popcount38_h9vn_out[0] = input_a[37];
  assign popcount38_h9vn_out[1] = popcount38_h9vn_core_282_not;
  assign popcount38_h9vn_out[2] = popcount38_h9vn_core_279;
  assign popcount38_h9vn_out[3] = popcount38_h9vn_core_284;
  assign popcount38_h9vn_out[4] = popcount38_h9vn_core_289;
  assign popcount38_h9vn_out[5] = 1'b0;
endmodule