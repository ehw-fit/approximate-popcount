// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.88739
// WCE=20.0
// EP=0.93127%
// Printed PDK parameters:
//  Area=19068938.0
//  Delay=40225548.0
//  Power=783400.0

module popcount39_je9w(input [38:0] input_a, output [5:0] popcount39_je9w_out);
  wire popcount39_je9w_core_041;
  wire popcount39_je9w_core_042;
  wire popcount39_je9w_core_043;
  wire popcount39_je9w_core_044;
  wire popcount39_je9w_core_045;
  wire popcount39_je9w_core_049;
  wire popcount39_je9w_core_050;
  wire popcount39_je9w_core_051;
  wire popcount39_je9w_core_052;
  wire popcount39_je9w_core_053;
  wire popcount39_je9w_core_054;
  wire popcount39_je9w_core_055;
  wire popcount39_je9w_core_056;
  wire popcount39_je9w_core_057;
  wire popcount39_je9w_core_058;
  wire popcount39_je9w_core_059;
  wire popcount39_je9w_core_060;
  wire popcount39_je9w_core_061;
  wire popcount39_je9w_core_063;
  wire popcount39_je9w_core_064;
  wire popcount39_je9w_core_065;
  wire popcount39_je9w_core_067;
  wire popcount39_je9w_core_068;
  wire popcount39_je9w_core_069;
  wire popcount39_je9w_core_070;
  wire popcount39_je9w_core_071;
  wire popcount39_je9w_core_072;
  wire popcount39_je9w_core_075;
  wire popcount39_je9w_core_076;
  wire popcount39_je9w_core_077;
  wire popcount39_je9w_core_078;
  wire popcount39_je9w_core_079;
  wire popcount39_je9w_core_081;
  wire popcount39_je9w_core_082;
  wire popcount39_je9w_core_083;
  wire popcount39_je9w_core_084;
  wire popcount39_je9w_core_087;
  wire popcount39_je9w_core_088;
  wire popcount39_je9w_core_089;
  wire popcount39_je9w_core_091;
  wire popcount39_je9w_core_093;
  wire popcount39_je9w_core_094;
  wire popcount39_je9w_core_095;
  wire popcount39_je9w_core_096;
  wire popcount39_je9w_core_097;
  wire popcount39_je9w_core_100;
  wire popcount39_je9w_core_101;
  wire popcount39_je9w_core_103;
  wire popcount39_je9w_core_108;
  wire popcount39_je9w_core_109;
  wire popcount39_je9w_core_110;
  wire popcount39_je9w_core_111;
  wire popcount39_je9w_core_113;
  wire popcount39_je9w_core_116_not;
  wire popcount39_je9w_core_117;
  wire popcount39_je9w_core_118;
  wire popcount39_je9w_core_119;
  wire popcount39_je9w_core_121;
  wire popcount39_je9w_core_122;
  wire popcount39_je9w_core_123;
  wire popcount39_je9w_core_124;
  wire popcount39_je9w_core_125;
  wire popcount39_je9w_core_126;
  wire popcount39_je9w_core_127;
  wire popcount39_je9w_core_128;
  wire popcount39_je9w_core_130;
  wire popcount39_je9w_core_133;
  wire popcount39_je9w_core_134;
  wire popcount39_je9w_core_136;
  wire popcount39_je9w_core_137;
  wire popcount39_je9w_core_138;
  wire popcount39_je9w_core_141;
  wire popcount39_je9w_core_142;
  wire popcount39_je9w_core_144;
  wire popcount39_je9w_core_146;
  wire popcount39_je9w_core_147;
  wire popcount39_je9w_core_148;
  wire popcount39_je9w_core_149;
  wire popcount39_je9w_core_150;
  wire popcount39_je9w_core_152;
  wire popcount39_je9w_core_154;
  wire popcount39_je9w_core_155;
  wire popcount39_je9w_core_157;
  wire popcount39_je9w_core_158;
  wire popcount39_je9w_core_159;
  wire popcount39_je9w_core_160;
  wire popcount39_je9w_core_161;
  wire popcount39_je9w_core_162;
  wire popcount39_je9w_core_163;
  wire popcount39_je9w_core_164;
  wire popcount39_je9w_core_167;
  wire popcount39_je9w_core_168;
  wire popcount39_je9w_core_169;
  wire popcount39_je9w_core_170;
  wire popcount39_je9w_core_171_not;
  wire popcount39_je9w_core_172;
  wire popcount39_je9w_core_174;
  wire popcount39_je9w_core_175;
  wire popcount39_je9w_core_178;
  wire popcount39_je9w_core_181;
  wire popcount39_je9w_core_182;
  wire popcount39_je9w_core_183;
  wire popcount39_je9w_core_185;
  wire popcount39_je9w_core_186;
  wire popcount39_je9w_core_187;
  wire popcount39_je9w_core_188;
  wire popcount39_je9w_core_193;
  wire popcount39_je9w_core_194;
  wire popcount39_je9w_core_196;
  wire popcount39_je9w_core_197;
  wire popcount39_je9w_core_202;
  wire popcount39_je9w_core_203;
  wire popcount39_je9w_core_204;
  wire popcount39_je9w_core_205;
  wire popcount39_je9w_core_206;
  wire popcount39_je9w_core_207;
  wire popcount39_je9w_core_208;
  wire popcount39_je9w_core_209;
  wire popcount39_je9w_core_212;
  wire popcount39_je9w_core_213;
  wire popcount39_je9w_core_216;
  wire popcount39_je9w_core_217;
  wire popcount39_je9w_core_219;
  wire popcount39_je9w_core_220;
  wire popcount39_je9w_core_222;
  wire popcount39_je9w_core_223;
  wire popcount39_je9w_core_226;
  wire popcount39_je9w_core_228;
  wire popcount39_je9w_core_229;
  wire popcount39_je9w_core_231;
  wire popcount39_je9w_core_232;
  wire popcount39_je9w_core_233;
  wire popcount39_je9w_core_236;
  wire popcount39_je9w_core_237;
  wire popcount39_je9w_core_240;
  wire popcount39_je9w_core_243;
  wire popcount39_je9w_core_244;
  wire popcount39_je9w_core_245;
  wire popcount39_je9w_core_246;
  wire popcount39_je9w_core_247_not;
  wire popcount39_je9w_core_248;
  wire popcount39_je9w_core_249;
  wire popcount39_je9w_core_250;
  wire popcount39_je9w_core_252;
  wire popcount39_je9w_core_253;
  wire popcount39_je9w_core_254;
  wire popcount39_je9w_core_255;
  wire popcount39_je9w_core_257;
  wire popcount39_je9w_core_259;
  wire popcount39_je9w_core_260_not;
  wire popcount39_je9w_core_262;
  wire popcount39_je9w_core_263;
  wire popcount39_je9w_core_264;
  wire popcount39_je9w_core_265;
  wire popcount39_je9w_core_266;
  wire popcount39_je9w_core_267;
  wire popcount39_je9w_core_270;
  wire popcount39_je9w_core_271;
  wire popcount39_je9w_core_272;
  wire popcount39_je9w_core_274;
  wire popcount39_je9w_core_275;
  wire popcount39_je9w_core_277;
  wire popcount39_je9w_core_278;
  wire popcount39_je9w_core_281;
  wire popcount39_je9w_core_282;
  wire popcount39_je9w_core_283;
  wire popcount39_je9w_core_284;
  wire popcount39_je9w_core_285;
  wire popcount39_je9w_core_286;
  wire popcount39_je9w_core_287;
  wire popcount39_je9w_core_289;
  wire popcount39_je9w_core_290;
  wire popcount39_je9w_core_291;
  wire popcount39_je9w_core_294;
  wire popcount39_je9w_core_295;
  wire popcount39_je9w_core_298;
  wire popcount39_je9w_core_299;
  wire popcount39_je9w_core_300_not;
  wire popcount39_je9w_core_301;
  wire popcount39_je9w_core_303;
  wire popcount39_je9w_core_304;
  wire popcount39_je9w_core_305;

  assign popcount39_je9w_core_041 = ~(input_a[7] & input_a[8]);
  assign popcount39_je9w_core_042 = input_a[12] & input_a[22];
  assign popcount39_je9w_core_043 = ~(input_a[24] & input_a[4]);
  assign popcount39_je9w_core_044 = input_a[19] & input_a[10];
  assign popcount39_je9w_core_045 = input_a[9] & input_a[29];
  assign popcount39_je9w_core_049 = ~(input_a[33] | input_a[25]);
  assign popcount39_je9w_core_050 = ~(input_a[12] ^ input_a[3]);
  assign popcount39_je9w_core_051 = input_a[18] & input_a[19];
  assign popcount39_je9w_core_052 = input_a[22] ^ input_a[26];
  assign popcount39_je9w_core_053 = input_a[34] | input_a[27];
  assign popcount39_je9w_core_054 = input_a[7] | input_a[2];
  assign popcount39_je9w_core_055 = input_a[13] | input_a[29];
  assign popcount39_je9w_core_056 = ~(input_a[9] & input_a[5]);
  assign popcount39_je9w_core_057 = ~(input_a[12] | input_a[9]);
  assign popcount39_je9w_core_058 = input_a[2] & input_a[0];
  assign popcount39_je9w_core_059 = ~input_a[6];
  assign popcount39_je9w_core_060 = ~input_a[31];
  assign popcount39_je9w_core_061 = ~input_a[11];
  assign popcount39_je9w_core_063 = ~(input_a[26] ^ input_a[3]);
  assign popcount39_je9w_core_064 = ~(input_a[12] | input_a[6]);
  assign popcount39_je9w_core_065 = ~(input_a[22] & input_a[38]);
  assign popcount39_je9w_core_067 = input_a[27] ^ input_a[29];
  assign popcount39_je9w_core_068 = ~(input_a[28] ^ input_a[28]);
  assign popcount39_je9w_core_069 = input_a[17] | input_a[16];
  assign popcount39_je9w_core_070 = ~input_a[2];
  assign popcount39_je9w_core_071 = ~(input_a[17] ^ input_a[30]);
  assign popcount39_je9w_core_072 = ~(input_a[19] & input_a[20]);
  assign popcount39_je9w_core_075 = input_a[30] & input_a[14];
  assign popcount39_je9w_core_076 = input_a[28] & input_a[6];
  assign popcount39_je9w_core_077 = input_a[0] | input_a[35];
  assign popcount39_je9w_core_078 = input_a[18] | input_a[23];
  assign popcount39_je9w_core_079 = input_a[5] ^ input_a[31];
  assign popcount39_je9w_core_081 = input_a[28] | input_a[17];
  assign popcount39_je9w_core_082 = input_a[20] ^ input_a[15];
  assign popcount39_je9w_core_083 = input_a[9] ^ input_a[10];
  assign popcount39_je9w_core_084 = input_a[9] & input_a[10];
  assign popcount39_je9w_core_087 = input_a[33] ^ input_a[30];
  assign popcount39_je9w_core_088 = ~(input_a[12] & input_a[35]);
  assign popcount39_je9w_core_089 = input_a[21] | input_a[14];
  assign popcount39_je9w_core_091 = ~(input_a[16] & input_a[0]);
  assign popcount39_je9w_core_093 = popcount39_je9w_core_084 ^ popcount39_je9w_core_089;
  assign popcount39_je9w_core_094 = input_a[9] & popcount39_je9w_core_089;
  assign popcount39_je9w_core_095 = popcount39_je9w_core_093 ^ popcount39_je9w_core_083;
  assign popcount39_je9w_core_096 = popcount39_je9w_core_093 & popcount39_je9w_core_083;
  assign popcount39_je9w_core_097 = popcount39_je9w_core_094 | popcount39_je9w_core_096;
  assign popcount39_je9w_core_100 = input_a[0] ^ input_a[36];
  assign popcount39_je9w_core_101 = input_a[29] & input_a[31];
  assign popcount39_je9w_core_103 = input_a[6] & input_a[25];
  assign popcount39_je9w_core_108 = input_a[3] | input_a[10];
  assign popcount39_je9w_core_109 = input_a[30] & input_a[8];
  assign popcount39_je9w_core_110 = popcount39_je9w_core_101 ^ popcount39_je9w_core_103;
  assign popcount39_je9w_core_111 = popcount39_je9w_core_101 & popcount39_je9w_core_103;
  assign popcount39_je9w_core_113 = ~(input_a[18] | input_a[30]);
  assign popcount39_je9w_core_116_not = ~input_a[28];
  assign popcount39_je9w_core_117 = input_a[18] & input_a[13];
  assign popcount39_je9w_core_118 = input_a[16] | input_a[36];
  assign popcount39_je9w_core_119 = popcount39_je9w_core_095 | popcount39_je9w_core_110;
  assign popcount39_je9w_core_121 = input_a[11] | input_a[11];
  assign popcount39_je9w_core_122 = popcount39_je9w_core_119 & input_a[1];
  assign popcount39_je9w_core_123 = popcount39_je9w_core_095 | popcount39_je9w_core_122;
  assign popcount39_je9w_core_124 = popcount39_je9w_core_097 ^ popcount39_je9w_core_111;
  assign popcount39_je9w_core_125 = popcount39_je9w_core_097 & popcount39_je9w_core_111;
  assign popcount39_je9w_core_126 = popcount39_je9w_core_124 ^ popcount39_je9w_core_123;
  assign popcount39_je9w_core_127 = popcount39_je9w_core_124 & popcount39_je9w_core_123;
  assign popcount39_je9w_core_128 = popcount39_je9w_core_125 | popcount39_je9w_core_127;
  assign popcount39_je9w_core_130 = input_a[36] ^ input_a[33];
  assign popcount39_je9w_core_133 = ~(input_a[32] & input_a[12]);
  assign popcount39_je9w_core_134 = ~(input_a[4] & input_a[8]);
  assign popcount39_je9w_core_136 = input_a[0] ^ input_a[15];
  assign popcount39_je9w_core_137 = input_a[31] | input_a[16];
  assign popcount39_je9w_core_138 = input_a[23] ^ input_a[31];
  assign popcount39_je9w_core_141 = popcount39_je9w_core_078 ^ popcount39_je9w_core_126;
  assign popcount39_je9w_core_142 = popcount39_je9w_core_078 & popcount39_je9w_core_126;
  assign popcount39_je9w_core_144 = ~(input_a[3] | input_a[15]);
  assign popcount39_je9w_core_146 = popcount39_je9w_core_081 ^ popcount39_je9w_core_128;
  assign popcount39_je9w_core_147 = popcount39_je9w_core_081 & popcount39_je9w_core_128;
  assign popcount39_je9w_core_148 = popcount39_je9w_core_146 ^ popcount39_je9w_core_142;
  assign popcount39_je9w_core_149 = popcount39_je9w_core_146 & popcount39_je9w_core_142;
  assign popcount39_je9w_core_150 = popcount39_je9w_core_147 | popcount39_je9w_core_149;
  assign popcount39_je9w_core_152 = ~(input_a[27] | input_a[20]);
  assign popcount39_je9w_core_154 = ~input_a[6];
  assign popcount39_je9w_core_155 = input_a[32] & input_a[28];
  assign popcount39_je9w_core_157 = input_a[13] | input_a[1];
  assign popcount39_je9w_core_158 = input_a[34] | input_a[23];
  assign popcount39_je9w_core_159 = ~(input_a[17] ^ input_a[20]);
  assign popcount39_je9w_core_160 = ~input_a[11];
  assign popcount39_je9w_core_161 = ~input_a[10];
  assign popcount39_je9w_core_162 = ~(input_a[6] ^ input_a[18]);
  assign popcount39_je9w_core_163 = input_a[32] ^ input_a[20];
  assign popcount39_je9w_core_164 = input_a[4] ^ input_a[18];
  assign popcount39_je9w_core_167 = input_a[38] & input_a[35];
  assign popcount39_je9w_core_168 = ~(input_a[32] & input_a[13]);
  assign popcount39_je9w_core_169 = ~(input_a[13] ^ input_a[16]);
  assign popcount39_je9w_core_170 = ~(input_a[32] ^ input_a[14]);
  assign popcount39_je9w_core_171_not = ~input_a[14];
  assign popcount39_je9w_core_172 = input_a[5] | input_a[1];
  assign popcount39_je9w_core_174 = input_a[3] & input_a[36];
  assign popcount39_je9w_core_175 = input_a[15] | input_a[17];
  assign popcount39_je9w_core_178 = input_a[19] | input_a[37];
  assign popcount39_je9w_core_181 = ~input_a[36];
  assign popcount39_je9w_core_182 = ~(input_a[2] | input_a[25]);
  assign popcount39_je9w_core_183 = input_a[6] ^ input_a[36];
  assign popcount39_je9w_core_185 = ~(input_a[25] & input_a[6]);
  assign popcount39_je9w_core_186 = ~(input_a[0] & input_a[35]);
  assign popcount39_je9w_core_187 = ~(input_a[14] | input_a[20]);
  assign popcount39_je9w_core_188 = input_a[5] ^ input_a[36];
  assign popcount39_je9w_core_193 = ~(input_a[9] | input_a[25]);
  assign popcount39_je9w_core_194 = input_a[12] & input_a[13];
  assign popcount39_je9w_core_196 = input_a[10] | input_a[34];
  assign popcount39_je9w_core_197 = input_a[38] | input_a[36];
  assign popcount39_je9w_core_202 = input_a[6] | input_a[27];
  assign popcount39_je9w_core_203 = input_a[23] | input_a[1];
  assign popcount39_je9w_core_204 = ~(input_a[11] | input_a[36]);
  assign popcount39_je9w_core_205 = input_a[16] | input_a[8];
  assign popcount39_je9w_core_206 = input_a[22] ^ input_a[35];
  assign popcount39_je9w_core_207 = input_a[15] | input_a[12];
  assign popcount39_je9w_core_208 = ~(input_a[14] | input_a[13]);
  assign popcount39_je9w_core_209 = ~(input_a[10] | input_a[0]);
  assign popcount39_je9w_core_212 = ~(input_a[5] & input_a[3]);
  assign popcount39_je9w_core_213 = ~input_a[24];
  assign popcount39_je9w_core_216 = input_a[36] ^ input_a[3];
  assign popcount39_je9w_core_217 = input_a[16] ^ input_a[26];
  assign popcount39_je9w_core_219 = input_a[25] | input_a[3];
  assign popcount39_je9w_core_220 = input_a[14] | input_a[33];
  assign popcount39_je9w_core_222 = ~(input_a[4] & input_a[8]);
  assign popcount39_je9w_core_223 = ~(input_a[22] & input_a[21]);
  assign popcount39_je9w_core_226 = input_a[0] | input_a[16];
  assign popcount39_je9w_core_228 = ~(input_a[34] & input_a[31]);
  assign popcount39_je9w_core_229 = ~(input_a[11] ^ input_a[18]);
  assign popcount39_je9w_core_231 = input_a[36] ^ input_a[29];
  assign popcount39_je9w_core_232 = ~(input_a[25] | input_a[3]);
  assign popcount39_je9w_core_233 = ~input_a[17];
  assign popcount39_je9w_core_236 = input_a[24] & input_a[14];
  assign popcount39_je9w_core_237 = input_a[38] & input_a[0];
  assign popcount39_je9w_core_240 = ~(input_a[20] | input_a[7]);
  assign popcount39_je9w_core_243 = ~(input_a[7] | input_a[20]);
  assign popcount39_je9w_core_244 = ~(input_a[1] & input_a[34]);
  assign popcount39_je9w_core_245 = input_a[28] ^ input_a[0];
  assign popcount39_je9w_core_246 = ~input_a[20];
  assign popcount39_je9w_core_247_not = ~input_a[8];
  assign popcount39_je9w_core_248 = ~(input_a[36] | input_a[27]);
  assign popcount39_je9w_core_249 = ~input_a[31];
  assign popcount39_je9w_core_250 = ~(input_a[37] ^ input_a[30]);
  assign popcount39_je9w_core_252 = input_a[8] | input_a[31];
  assign popcount39_je9w_core_253 = ~(input_a[19] | input_a[17]);
  assign popcount39_je9w_core_254 = ~(input_a[31] | input_a[18]);
  assign popcount39_je9w_core_255 = ~(input_a[17] ^ input_a[2]);
  assign popcount39_je9w_core_257 = input_a[32] & input_a[24];
  assign popcount39_je9w_core_259 = ~(input_a[21] ^ input_a[7]);
  assign popcount39_je9w_core_260_not = ~input_a[1];
  assign popcount39_je9w_core_262 = input_a[28] & input_a[31];
  assign popcount39_je9w_core_263 = ~(input_a[5] | input_a[10]);
  assign popcount39_je9w_core_264 = ~(input_a[17] ^ input_a[21]);
  assign popcount39_je9w_core_265 = ~(input_a[13] | input_a[32]);
  assign popcount39_je9w_core_266 = ~input_a[29];
  assign popcount39_je9w_core_267 = ~input_a[20];
  assign popcount39_je9w_core_270 = ~input_a[15];
  assign popcount39_je9w_core_271 = ~input_a[38];
  assign popcount39_je9w_core_272 = input_a[26] ^ input_a[13];
  assign popcount39_je9w_core_274 = input_a[32] | input_a[28];
  assign popcount39_je9w_core_275 = input_a[0] & input_a[24];
  assign popcount39_je9w_core_277 = ~(input_a[38] ^ input_a[24]);
  assign popcount39_je9w_core_278 = input_a[1] | input_a[31];
  assign popcount39_je9w_core_281 = input_a[34] & input_a[5];
  assign popcount39_je9w_core_282 = ~input_a[38];
  assign popcount39_je9w_core_283 = input_a[37] | input_a[32];
  assign popcount39_je9w_core_284 = popcount39_je9w_core_282 ^ popcount39_je9w_core_281;
  assign popcount39_je9w_core_285 = input_a[34] & input_a[5];
  assign popcount39_je9w_core_286 = input_a[38] | popcount39_je9w_core_285;
  assign popcount39_je9w_core_287 = ~popcount39_je9w_core_141;
  assign popcount39_je9w_core_289 = popcount39_je9w_core_287 ^ popcount39_je9w_core_286;
  assign popcount39_je9w_core_290 = popcount39_je9w_core_287 & popcount39_je9w_core_286;
  assign popcount39_je9w_core_291 = popcount39_je9w_core_141 | popcount39_je9w_core_290;
  assign popcount39_je9w_core_294 = popcount39_je9w_core_148 ^ popcount39_je9w_core_291;
  assign popcount39_je9w_core_295 = popcount39_je9w_core_148 & popcount39_je9w_core_291;
  assign popcount39_je9w_core_298 = input_a[34] ^ input_a[34];
  assign popcount39_je9w_core_299 = popcount39_je9w_core_150 | popcount39_je9w_core_295;
  assign popcount39_je9w_core_300_not = ~input_a[34];
  assign popcount39_je9w_core_301 = ~(input_a[3] ^ input_a[26]);
  assign popcount39_je9w_core_303 = input_a[13] ^ input_a[36];
  assign popcount39_je9w_core_304 = input_a[25] & input_a[24];
  assign popcount39_je9w_core_305 = input_a[1] ^ input_a[10];

  assign popcount39_je9w_out[0] = input_a[20];
  assign popcount39_je9w_out[1] = popcount39_je9w_core_284;
  assign popcount39_je9w_out[2] = popcount39_je9w_core_289;
  assign popcount39_je9w_out[3] = popcount39_je9w_core_294;
  assign popcount39_je9w_out[4] = popcount39_je9w_core_299;
  assign popcount39_je9w_out[5] = 1'b0;
endmodule