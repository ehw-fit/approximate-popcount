// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=11.0013
// WCE=27.0
// EP=0.998417%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_ajog(input [23:0] input_a, output [4:0] popcount24_ajog_out);
  wire popcount24_ajog_core_026;
  wire popcount24_ajog_core_027;
  wire popcount24_ajog_core_028;
  wire popcount24_ajog_core_029;
  wire popcount24_ajog_core_030;
  wire popcount24_ajog_core_031;
  wire popcount24_ajog_core_032;
  wire popcount24_ajog_core_035;
  wire popcount24_ajog_core_036;
  wire popcount24_ajog_core_038;
  wire popcount24_ajog_core_039;
  wire popcount24_ajog_core_040;
  wire popcount24_ajog_core_041;
  wire popcount24_ajog_core_042;
  wire popcount24_ajog_core_043;
  wire popcount24_ajog_core_046;
  wire popcount24_ajog_core_048;
  wire popcount24_ajog_core_049;
  wire popcount24_ajog_core_051;
  wire popcount24_ajog_core_052;
  wire popcount24_ajog_core_053;
  wire popcount24_ajog_core_054;
  wire popcount24_ajog_core_056;
  wire popcount24_ajog_core_058;
  wire popcount24_ajog_core_060;
  wire popcount24_ajog_core_061;
  wire popcount24_ajog_core_062;
  wire popcount24_ajog_core_063;
  wire popcount24_ajog_core_066;
  wire popcount24_ajog_core_067;
  wire popcount24_ajog_core_069_not;
  wire popcount24_ajog_core_071;
  wire popcount24_ajog_core_072;
  wire popcount24_ajog_core_073_not;
  wire popcount24_ajog_core_075;
  wire popcount24_ajog_core_076;
  wire popcount24_ajog_core_077;
  wire popcount24_ajog_core_080;
  wire popcount24_ajog_core_081;
  wire popcount24_ajog_core_083_not;
  wire popcount24_ajog_core_087;
  wire popcount24_ajog_core_091;
  wire popcount24_ajog_core_094;
  wire popcount24_ajog_core_096;
  wire popcount24_ajog_core_097;
  wire popcount24_ajog_core_099;
  wire popcount24_ajog_core_100_not;
  wire popcount24_ajog_core_101;
  wire popcount24_ajog_core_102;
  wire popcount24_ajog_core_103;
  wire popcount24_ajog_core_104_not;
  wire popcount24_ajog_core_105;
  wire popcount24_ajog_core_107_not;
  wire popcount24_ajog_core_110;
  wire popcount24_ajog_core_111;
  wire popcount24_ajog_core_113;
  wire popcount24_ajog_core_114;
  wire popcount24_ajog_core_115;
  wire popcount24_ajog_core_116;
  wire popcount24_ajog_core_117;
  wire popcount24_ajog_core_118;
  wire popcount24_ajog_core_120;
  wire popcount24_ajog_core_122;
  wire popcount24_ajog_core_123;
  wire popcount24_ajog_core_124;
  wire popcount24_ajog_core_125;
  wire popcount24_ajog_core_126;
  wire popcount24_ajog_core_128;
  wire popcount24_ajog_core_130;
  wire popcount24_ajog_core_134;
  wire popcount24_ajog_core_135;
  wire popcount24_ajog_core_136;
  wire popcount24_ajog_core_138;
  wire popcount24_ajog_core_139;
  wire popcount24_ajog_core_142;
  wire popcount24_ajog_core_143;
  wire popcount24_ajog_core_145;
  wire popcount24_ajog_core_146;
  wire popcount24_ajog_core_147;
  wire popcount24_ajog_core_149;
  wire popcount24_ajog_core_150;
  wire popcount24_ajog_core_151;
  wire popcount24_ajog_core_152;
  wire popcount24_ajog_core_154;
  wire popcount24_ajog_core_156;
  wire popcount24_ajog_core_158;
  wire popcount24_ajog_core_162;
  wire popcount24_ajog_core_164;
  wire popcount24_ajog_core_166;
  wire popcount24_ajog_core_167;
  wire popcount24_ajog_core_171;
  wire popcount24_ajog_core_172;
  wire popcount24_ajog_core_173;
  wire popcount24_ajog_core_175;
  wire popcount24_ajog_core_176_not;
  wire popcount24_ajog_core_177;

  assign popcount24_ajog_core_026 = ~(input_a[18] & input_a[3]);
  assign popcount24_ajog_core_027 = input_a[17] ^ input_a[4];
  assign popcount24_ajog_core_028 = input_a[4] & input_a[10];
  assign popcount24_ajog_core_029 = ~(input_a[6] ^ input_a[0]);
  assign popcount24_ajog_core_030 = input_a[3] & input_a[4];
  assign popcount24_ajog_core_031 = input_a[19] ^ input_a[17];
  assign popcount24_ajog_core_032 = input_a[16] ^ input_a[14];
  assign popcount24_ajog_core_035 = ~input_a[2];
  assign popcount24_ajog_core_036 = input_a[13] ^ input_a[2];
  assign popcount24_ajog_core_038 = ~(input_a[2] ^ input_a[4]);
  assign popcount24_ajog_core_039 = ~(input_a[7] & input_a[21]);
  assign popcount24_ajog_core_040 = ~input_a[20];
  assign popcount24_ajog_core_041 = ~(input_a[3] & input_a[18]);
  assign popcount24_ajog_core_042 = input_a[2] | input_a[20];
  assign popcount24_ajog_core_043 = ~input_a[0];
  assign popcount24_ajog_core_046 = ~(input_a[15] ^ input_a[5]);
  assign popcount24_ajog_core_048 = input_a[9] | input_a[4];
  assign popcount24_ajog_core_049 = input_a[7] ^ input_a[9];
  assign popcount24_ajog_core_051 = ~(input_a[21] & input_a[3]);
  assign popcount24_ajog_core_052 = input_a[22] ^ input_a[23];
  assign popcount24_ajog_core_053 = input_a[19] ^ input_a[13];
  assign popcount24_ajog_core_054 = input_a[4] ^ input_a[22];
  assign popcount24_ajog_core_056 = input_a[8] ^ input_a[11];
  assign popcount24_ajog_core_058 = input_a[14] ^ input_a[16];
  assign popcount24_ajog_core_060 = input_a[20] & input_a[22];
  assign popcount24_ajog_core_061 = ~(input_a[22] | input_a[15]);
  assign popcount24_ajog_core_062 = input_a[1] | input_a[2];
  assign popcount24_ajog_core_063 = ~(input_a[10] & input_a[14]);
  assign popcount24_ajog_core_066 = ~(input_a[14] ^ input_a[2]);
  assign popcount24_ajog_core_067 = input_a[11] & input_a[6];
  assign popcount24_ajog_core_069_not = ~input_a[10];
  assign popcount24_ajog_core_071 = input_a[10] & input_a[11];
  assign popcount24_ajog_core_072 = input_a[3] ^ input_a[1];
  assign popcount24_ajog_core_073_not = ~input_a[22];
  assign popcount24_ajog_core_075 = input_a[4] & input_a[1];
  assign popcount24_ajog_core_076 = ~(input_a[17] ^ input_a[15]);
  assign popcount24_ajog_core_077 = ~(input_a[6] | input_a[7]);
  assign popcount24_ajog_core_080 = ~input_a[10];
  assign popcount24_ajog_core_081 = ~(input_a[12] & input_a[1]);
  assign popcount24_ajog_core_083_not = ~input_a[20];
  assign popcount24_ajog_core_087 = ~(input_a[23] ^ input_a[10]);
  assign popcount24_ajog_core_091 = ~(input_a[18] | input_a[7]);
  assign popcount24_ajog_core_094 = ~(input_a[19] ^ input_a[17]);
  assign popcount24_ajog_core_096 = input_a[5] | input_a[21];
  assign popcount24_ajog_core_097 = ~input_a[1];
  assign popcount24_ajog_core_099 = input_a[20] | input_a[12];
  assign popcount24_ajog_core_100_not = ~input_a[10];
  assign popcount24_ajog_core_101 = ~(input_a[11] & input_a[7]);
  assign popcount24_ajog_core_102 = ~(input_a[5] | input_a[7]);
  assign popcount24_ajog_core_103 = ~(input_a[4] ^ input_a[2]);
  assign popcount24_ajog_core_104_not = ~input_a[21];
  assign popcount24_ajog_core_105 = ~(input_a[3] ^ input_a[9]);
  assign popcount24_ajog_core_107_not = ~input_a[9];
  assign popcount24_ajog_core_110 = input_a[12] & input_a[14];
  assign popcount24_ajog_core_111 = ~input_a[19];
  assign popcount24_ajog_core_113 = ~(input_a[10] ^ input_a[13]);
  assign popcount24_ajog_core_114 = ~input_a[9];
  assign popcount24_ajog_core_115 = ~(input_a[22] ^ input_a[14]);
  assign popcount24_ajog_core_116 = ~input_a[0];
  assign popcount24_ajog_core_117 = ~input_a[1];
  assign popcount24_ajog_core_118 = input_a[19] | input_a[17];
  assign popcount24_ajog_core_120 = input_a[18] ^ input_a[4];
  assign popcount24_ajog_core_122 = input_a[20] & input_a[19];
  assign popcount24_ajog_core_123 = input_a[8] | input_a[3];
  assign popcount24_ajog_core_124 = ~input_a[4];
  assign popcount24_ajog_core_125 = ~(input_a[18] ^ input_a[2]);
  assign popcount24_ajog_core_126 = input_a[16] & input_a[12];
  assign popcount24_ajog_core_128 = input_a[14] & input_a[5];
  assign popcount24_ajog_core_130 = input_a[11] & input_a[5];
  assign popcount24_ajog_core_134 = input_a[20] ^ input_a[5];
  assign popcount24_ajog_core_135 = ~(input_a[19] | input_a[6]);
  assign popcount24_ajog_core_136 = input_a[7] ^ input_a[5];
  assign popcount24_ajog_core_138 = ~input_a[22];
  assign popcount24_ajog_core_139 = ~(input_a[4] | input_a[9]);
  assign popcount24_ajog_core_142 = input_a[22] & input_a[21];
  assign popcount24_ajog_core_143 = ~(input_a[3] ^ input_a[20]);
  assign popcount24_ajog_core_145 = ~(input_a[2] ^ input_a[6]);
  assign popcount24_ajog_core_146 = ~(input_a[19] ^ input_a[14]);
  assign popcount24_ajog_core_147 = input_a[11] | input_a[13];
  assign popcount24_ajog_core_149 = input_a[14] & input_a[6];
  assign popcount24_ajog_core_150 = ~(input_a[23] | input_a[3]);
  assign popcount24_ajog_core_151 = ~(input_a[6] ^ input_a[9]);
  assign popcount24_ajog_core_152 = input_a[7] ^ input_a[22];
  assign popcount24_ajog_core_154 = ~(input_a[2] ^ input_a[9]);
  assign popcount24_ajog_core_156 = input_a[21] ^ input_a[13];
  assign popcount24_ajog_core_158 = ~(input_a[5] & input_a[8]);
  assign popcount24_ajog_core_162 = input_a[3] | input_a[22];
  assign popcount24_ajog_core_164 = ~input_a[8];
  assign popcount24_ajog_core_166 = input_a[8] ^ input_a[14];
  assign popcount24_ajog_core_167 = ~(input_a[3] & input_a[0]);
  assign popcount24_ajog_core_171 = ~input_a[16];
  assign popcount24_ajog_core_172 = input_a[16] | input_a[21];
  assign popcount24_ajog_core_173 = ~input_a[4];
  assign popcount24_ajog_core_175 = ~input_a[4];
  assign popcount24_ajog_core_176_not = ~input_a[7];
  assign popcount24_ajog_core_177 = input_a[6] ^ input_a[10];

  assign popcount24_ajog_out[0] = 1'b0;
  assign popcount24_ajog_out[1] = input_a[19];
  assign popcount24_ajog_out[2] = input_a[15];
  assign popcount24_ajog_out[3] = input_a[23];
  assign popcount24_ajog_out[4] = 1'b1;
endmodule