// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.89636
// WCE=20.0
// EP=0.930242%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_b0rq(input [31:0] input_a, output [5:0] popcount32_b0rq_out);
  wire popcount32_b0rq_core_035;
  wire popcount32_b0rq_core_041_not;
  wire popcount32_b0rq_core_045;
  wire popcount32_b0rq_core_046;
  wire popcount32_b0rq_core_047;
  wire popcount32_b0rq_core_048_not;
  wire popcount32_b0rq_core_049;
  wire popcount32_b0rq_core_051;
  wire popcount32_b0rq_core_053;
  wire popcount32_b0rq_core_054;
  wire popcount32_b0rq_core_056;
  wire popcount32_b0rq_core_059;
  wire popcount32_b0rq_core_063;
  wire popcount32_b0rq_core_066;
  wire popcount32_b0rq_core_068;
  wire popcount32_b0rq_core_070;
  wire popcount32_b0rq_core_071;
  wire popcount32_b0rq_core_072;
  wire popcount32_b0rq_core_073;
  wire popcount32_b0rq_core_075;
  wire popcount32_b0rq_core_076;
  wire popcount32_b0rq_core_077;
  wire popcount32_b0rq_core_078;
  wire popcount32_b0rq_core_079;
  wire popcount32_b0rq_core_082;
  wire popcount32_b0rq_core_083;
  wire popcount32_b0rq_core_084;
  wire popcount32_b0rq_core_085;
  wire popcount32_b0rq_core_086;
  wire popcount32_b0rq_core_087;
  wire popcount32_b0rq_core_091;
  wire popcount32_b0rq_core_092;
  wire popcount32_b0rq_core_093;
  wire popcount32_b0rq_core_096;
  wire popcount32_b0rq_core_097_not;
  wire popcount32_b0rq_core_098;
  wire popcount32_b0rq_core_100;
  wire popcount32_b0rq_core_102;
  wire popcount32_b0rq_core_105;
  wire popcount32_b0rq_core_106;
  wire popcount32_b0rq_core_107;
  wire popcount32_b0rq_core_110;
  wire popcount32_b0rq_core_111;
  wire popcount32_b0rq_core_112;
  wire popcount32_b0rq_core_113;
  wire popcount32_b0rq_core_114;
  wire popcount32_b0rq_core_115;
  wire popcount32_b0rq_core_116_not;
  wire popcount32_b0rq_core_118;
  wire popcount32_b0rq_core_119;
  wire popcount32_b0rq_core_122;
  wire popcount32_b0rq_core_123;
  wire popcount32_b0rq_core_124;
  wire popcount32_b0rq_core_125;
  wire popcount32_b0rq_core_127;
  wire popcount32_b0rq_core_130;
  wire popcount32_b0rq_core_131_not;
  wire popcount32_b0rq_core_132;
  wire popcount32_b0rq_core_133;
  wire popcount32_b0rq_core_136;
  wire popcount32_b0rq_core_137;
  wire popcount32_b0rq_core_139;
  wire popcount32_b0rq_core_140_not;
  wire popcount32_b0rq_core_142;
  wire popcount32_b0rq_core_143;
  wire popcount32_b0rq_core_144;
  wire popcount32_b0rq_core_145;
  wire popcount32_b0rq_core_147;
  wire popcount32_b0rq_core_148;
  wire popcount32_b0rq_core_150;
  wire popcount32_b0rq_core_153;
  wire popcount32_b0rq_core_154;
  wire popcount32_b0rq_core_155;
  wire popcount32_b0rq_core_157_not;
  wire popcount32_b0rq_core_159;
  wire popcount32_b0rq_core_160;
  wire popcount32_b0rq_core_164;
  wire popcount32_b0rq_core_165;
  wire popcount32_b0rq_core_166;
  wire popcount32_b0rq_core_167;
  wire popcount32_b0rq_core_168;
  wire popcount32_b0rq_core_171;
  wire popcount32_b0rq_core_172;
  wire popcount32_b0rq_core_173;
  wire popcount32_b0rq_core_176;
  wire popcount32_b0rq_core_178;
  wire popcount32_b0rq_core_179;
  wire popcount32_b0rq_core_181;
  wire popcount32_b0rq_core_182;
  wire popcount32_b0rq_core_183;
  wire popcount32_b0rq_core_184;
  wire popcount32_b0rq_core_185;
  wire popcount32_b0rq_core_186;
  wire popcount32_b0rq_core_187_not;
  wire popcount32_b0rq_core_188;
  wire popcount32_b0rq_core_189;
  wire popcount32_b0rq_core_190;
  wire popcount32_b0rq_core_195;
  wire popcount32_b0rq_core_197;
  wire popcount32_b0rq_core_199;
  wire popcount32_b0rq_core_200;
  wire popcount32_b0rq_core_201;
  wire popcount32_b0rq_core_203;
  wire popcount32_b0rq_core_207;
  wire popcount32_b0rq_core_208;
  wire popcount32_b0rq_core_209;
  wire popcount32_b0rq_core_212;
  wire popcount32_b0rq_core_213;
  wire popcount32_b0rq_core_214;
  wire popcount32_b0rq_core_216;
  wire popcount32_b0rq_core_217;
  wire popcount32_b0rq_core_219;
  wire popcount32_b0rq_core_221;
  wire popcount32_b0rq_core_222;
  wire popcount32_b0rq_core_223;
  wire popcount32_b0rq_core_224_not;
  wire popcount32_b0rq_core_225;

  assign popcount32_b0rq_core_035 = input_a[16] ^ input_a[28];
  assign popcount32_b0rq_core_041_not = ~input_a[27];
  assign popcount32_b0rq_core_045 = ~(input_a[25] | input_a[30]);
  assign popcount32_b0rq_core_046 = input_a[25] & input_a[12];
  assign popcount32_b0rq_core_047 = ~(input_a[22] & input_a[25]);
  assign popcount32_b0rq_core_048_not = ~input_a[20];
  assign popcount32_b0rq_core_049 = input_a[28] & input_a[15];
  assign popcount32_b0rq_core_051 = input_a[2] & input_a[18];
  assign popcount32_b0rq_core_053 = ~input_a[18];
  assign popcount32_b0rq_core_054 = input_a[14] ^ input_a[1];
  assign popcount32_b0rq_core_056 = ~(input_a[31] | input_a[26]);
  assign popcount32_b0rq_core_059 = ~(input_a[28] ^ input_a[14]);
  assign popcount32_b0rq_core_063 = ~(input_a[22] | input_a[30]);
  assign popcount32_b0rq_core_066 = ~input_a[30];
  assign popcount32_b0rq_core_068 = ~(input_a[4] | input_a[20]);
  assign popcount32_b0rq_core_070 = input_a[3] & input_a[18];
  assign popcount32_b0rq_core_071 = ~(input_a[19] ^ input_a[19]);
  assign popcount32_b0rq_core_072 = ~(input_a[4] & input_a[8]);
  assign popcount32_b0rq_core_073 = input_a[14] | input_a[2];
  assign popcount32_b0rq_core_075 = ~(input_a[17] ^ input_a[16]);
  assign popcount32_b0rq_core_076 = input_a[12] & input_a[18];
  assign popcount32_b0rq_core_077 = ~(input_a[26] & input_a[5]);
  assign popcount32_b0rq_core_078 = input_a[13] ^ input_a[7];
  assign popcount32_b0rq_core_079 = ~(input_a[3] | input_a[16]);
  assign popcount32_b0rq_core_082 = input_a[4] & input_a[15];
  assign popcount32_b0rq_core_083 = input_a[10] | input_a[7];
  assign popcount32_b0rq_core_084 = input_a[7] & input_a[19];
  assign popcount32_b0rq_core_085 = ~(input_a[14] ^ input_a[24]);
  assign popcount32_b0rq_core_086 = ~(input_a[4] | input_a[20]);
  assign popcount32_b0rq_core_087 = ~(input_a[14] | input_a[18]);
  assign popcount32_b0rq_core_091 = input_a[28] & input_a[14];
  assign popcount32_b0rq_core_092 = input_a[19] & input_a[13];
  assign popcount32_b0rq_core_093 = ~(input_a[16] ^ input_a[30]);
  assign popcount32_b0rq_core_096 = ~(input_a[30] | input_a[26]);
  assign popcount32_b0rq_core_097_not = ~input_a[20];
  assign popcount32_b0rq_core_098 = input_a[10] | input_a[18];
  assign popcount32_b0rq_core_100 = ~(input_a[18] ^ input_a[26]);
  assign popcount32_b0rq_core_102 = ~(input_a[25] ^ input_a[2]);
  assign popcount32_b0rq_core_105 = input_a[11] ^ input_a[2];
  assign popcount32_b0rq_core_106 = input_a[12] & input_a[16];
  assign popcount32_b0rq_core_107 = ~input_a[7];
  assign popcount32_b0rq_core_110 = input_a[4] ^ input_a[16];
  assign popcount32_b0rq_core_111 = ~(input_a[8] & input_a[30]);
  assign popcount32_b0rq_core_112 = ~(input_a[12] & input_a[27]);
  assign popcount32_b0rq_core_113 = ~(input_a[20] & input_a[20]);
  assign popcount32_b0rq_core_114 = ~(input_a[5] ^ input_a[22]);
  assign popcount32_b0rq_core_115 = ~(input_a[1] ^ input_a[1]);
  assign popcount32_b0rq_core_116_not = ~input_a[25];
  assign popcount32_b0rq_core_118 = ~(input_a[25] ^ input_a[14]);
  assign popcount32_b0rq_core_119 = input_a[25] | input_a[30];
  assign popcount32_b0rq_core_122 = ~(input_a[22] | input_a[12]);
  assign popcount32_b0rq_core_123 = input_a[0] & input_a[0];
  assign popcount32_b0rq_core_124 = ~input_a[16];
  assign popcount32_b0rq_core_125 = ~(input_a[28] | input_a[29]);
  assign popcount32_b0rq_core_127 = ~(input_a[17] | input_a[17]);
  assign popcount32_b0rq_core_130 = input_a[14] | input_a[14];
  assign popcount32_b0rq_core_131_not = ~input_a[29];
  assign popcount32_b0rq_core_132 = ~input_a[19];
  assign popcount32_b0rq_core_133 = input_a[20] | input_a[7];
  assign popcount32_b0rq_core_136 = ~(input_a[6] ^ input_a[9]);
  assign popcount32_b0rq_core_137 = input_a[26] | input_a[25];
  assign popcount32_b0rq_core_139 = ~input_a[12];
  assign popcount32_b0rq_core_140_not = ~input_a[0];
  assign popcount32_b0rq_core_142 = input_a[26] & input_a[13];
  assign popcount32_b0rq_core_143 = ~input_a[17];
  assign popcount32_b0rq_core_144 = input_a[15] & input_a[2];
  assign popcount32_b0rq_core_145 = ~(input_a[8] & input_a[19]);
  assign popcount32_b0rq_core_147 = ~(input_a[29] | input_a[0]);
  assign popcount32_b0rq_core_148 = input_a[6] & input_a[7];
  assign popcount32_b0rq_core_150 = ~input_a[29];
  assign popcount32_b0rq_core_153 = ~(input_a[1] ^ input_a[14]);
  assign popcount32_b0rq_core_154 = input_a[11] | input_a[24];
  assign popcount32_b0rq_core_155 = ~(input_a[13] & input_a[11]);
  assign popcount32_b0rq_core_157_not = ~input_a[13];
  assign popcount32_b0rq_core_159 = input_a[1] & input_a[5];
  assign popcount32_b0rq_core_160 = ~(input_a[16] | input_a[15]);
  assign popcount32_b0rq_core_164 = ~input_a[10];
  assign popcount32_b0rq_core_165 = input_a[31] & input_a[13];
  assign popcount32_b0rq_core_166 = ~(input_a[13] & input_a[9]);
  assign popcount32_b0rq_core_167 = input_a[12] | input_a[2];
  assign popcount32_b0rq_core_168 = ~input_a[8];
  assign popcount32_b0rq_core_171 = input_a[26] ^ input_a[2];
  assign popcount32_b0rq_core_172 = ~(input_a[21] & input_a[17]);
  assign popcount32_b0rq_core_173 = ~(input_a[2] | input_a[19]);
  assign popcount32_b0rq_core_176 = ~input_a[1];
  assign popcount32_b0rq_core_178 = ~input_a[21];
  assign popcount32_b0rq_core_179 = ~(input_a[14] ^ input_a[22]);
  assign popcount32_b0rq_core_181 = input_a[16] | input_a[30];
  assign popcount32_b0rq_core_182 = ~(input_a[20] | input_a[24]);
  assign popcount32_b0rq_core_183 = ~(input_a[6] ^ input_a[27]);
  assign popcount32_b0rq_core_184 = ~(input_a[0] & input_a[4]);
  assign popcount32_b0rq_core_185 = input_a[10] ^ input_a[27];
  assign popcount32_b0rq_core_186 = input_a[26] & input_a[10];
  assign popcount32_b0rq_core_187_not = ~input_a[16];
  assign popcount32_b0rq_core_188 = input_a[30] ^ input_a[3];
  assign popcount32_b0rq_core_189 = ~(input_a[11] ^ input_a[10]);
  assign popcount32_b0rq_core_190 = ~(input_a[14] | input_a[7]);
  assign popcount32_b0rq_core_195 = ~(input_a[9] ^ input_a[22]);
  assign popcount32_b0rq_core_197 = ~(input_a[22] ^ input_a[27]);
  assign popcount32_b0rq_core_199 = input_a[26] & input_a[13];
  assign popcount32_b0rq_core_200 = input_a[13] ^ input_a[2];
  assign popcount32_b0rq_core_201 = input_a[10] | input_a[4];
  assign popcount32_b0rq_core_203 = ~(input_a[23] & input_a[12]);
  assign popcount32_b0rq_core_207 = ~(input_a[9] | input_a[6]);
  assign popcount32_b0rq_core_208 = input_a[0] & input_a[12];
  assign popcount32_b0rq_core_209 = ~(input_a[21] ^ input_a[7]);
  assign popcount32_b0rq_core_212 = ~input_a[12];
  assign popcount32_b0rq_core_213 = ~(input_a[3] & input_a[26]);
  assign popcount32_b0rq_core_214 = ~(input_a[0] & input_a[18]);
  assign popcount32_b0rq_core_216 = ~(input_a[28] | input_a[6]);
  assign popcount32_b0rq_core_217 = input_a[14] ^ input_a[7];
  assign popcount32_b0rq_core_219 = input_a[1] | input_a[11];
  assign popcount32_b0rq_core_221 = input_a[14] ^ input_a[30];
  assign popcount32_b0rq_core_222 = input_a[21] | input_a[15];
  assign popcount32_b0rq_core_223 = ~(input_a[28] & input_a[1]);
  assign popcount32_b0rq_core_224_not = ~input_a[10];
  assign popcount32_b0rq_core_225 = ~(input_a[17] ^ input_a[11]);

  assign popcount32_b0rq_out[0] = input_a[2];
  assign popcount32_b0rq_out[1] = input_a[19];
  assign popcount32_b0rq_out[2] = input_a[1];
  assign popcount32_b0rq_out[3] = 1'b0;
  assign popcount32_b0rq_out[4] = 1'b1;
  assign popcount32_b0rq_out[5] = 1'b0;
endmodule