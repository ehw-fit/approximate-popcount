// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.31143
// WCE=16.0
// EP=0.864565%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_xsys(input [30:0] input_a, output [4:0] popcount31_xsys_out);
  wire popcount31_xsys_core_036;
  wire popcount31_xsys_core_038_not;
  wire popcount31_xsys_core_039;
  wire popcount31_xsys_core_040;
  wire popcount31_xsys_core_041;
  wire popcount31_xsys_core_042;
  wire popcount31_xsys_core_043;
  wire popcount31_xsys_core_044;
  wire popcount31_xsys_core_045;
  wire popcount31_xsys_core_047;
  wire popcount31_xsys_core_048;
  wire popcount31_xsys_core_049;
  wire popcount31_xsys_core_050;
  wire popcount31_xsys_core_051;
  wire popcount31_xsys_core_052;
  wire popcount31_xsys_core_053;
  wire popcount31_xsys_core_057;
  wire popcount31_xsys_core_058;
  wire popcount31_xsys_core_060;
  wire popcount31_xsys_core_062;
  wire popcount31_xsys_core_063;
  wire popcount31_xsys_core_064;
  wire popcount31_xsys_core_065;
  wire popcount31_xsys_core_066;
  wire popcount31_xsys_core_067;
  wire popcount31_xsys_core_068;
  wire popcount31_xsys_core_072;
  wire popcount31_xsys_core_073;
  wire popcount31_xsys_core_075;
  wire popcount31_xsys_core_076;
  wire popcount31_xsys_core_078;
  wire popcount31_xsys_core_079;
  wire popcount31_xsys_core_080;
  wire popcount31_xsys_core_081_not;
  wire popcount31_xsys_core_082;
  wire popcount31_xsys_core_085;
  wire popcount31_xsys_core_088;
  wire popcount31_xsys_core_091;
  wire popcount31_xsys_core_092;
  wire popcount31_xsys_core_095;
  wire popcount31_xsys_core_097;
  wire popcount31_xsys_core_098;
  wire popcount31_xsys_core_099;
  wire popcount31_xsys_core_101;
  wire popcount31_xsys_core_102;
  wire popcount31_xsys_core_103;
  wire popcount31_xsys_core_104;
  wire popcount31_xsys_core_105;
  wire popcount31_xsys_core_106;
  wire popcount31_xsys_core_107;
  wire popcount31_xsys_core_108;
  wire popcount31_xsys_core_109;
  wire popcount31_xsys_core_111;
  wire popcount31_xsys_core_113;
  wire popcount31_xsys_core_114;
  wire popcount31_xsys_core_117;
  wire popcount31_xsys_core_119;
  wire popcount31_xsys_core_120;
  wire popcount31_xsys_core_121;
  wire popcount31_xsys_core_124;
  wire popcount31_xsys_core_127;
  wire popcount31_xsys_core_129;
  wire popcount31_xsys_core_133;
  wire popcount31_xsys_core_135;
  wire popcount31_xsys_core_136;
  wire popcount31_xsys_core_138;
  wire popcount31_xsys_core_140;
  wire popcount31_xsys_core_142;
  wire popcount31_xsys_core_143;
  wire popcount31_xsys_core_144;
  wire popcount31_xsys_core_145;
  wire popcount31_xsys_core_148;
  wire popcount31_xsys_core_150;
  wire popcount31_xsys_core_151_not;
  wire popcount31_xsys_core_152;
  wire popcount31_xsys_core_153;
  wire popcount31_xsys_core_154;
  wire popcount31_xsys_core_155;
  wire popcount31_xsys_core_156;
  wire popcount31_xsys_core_158;
  wire popcount31_xsys_core_159;
  wire popcount31_xsys_core_160;
  wire popcount31_xsys_core_161;
  wire popcount31_xsys_core_162;
  wire popcount31_xsys_core_163;
  wire popcount31_xsys_core_166;
  wire popcount31_xsys_core_167;
  wire popcount31_xsys_core_168;
  wire popcount31_xsys_core_169;
  wire popcount31_xsys_core_171;
  wire popcount31_xsys_core_172;
  wire popcount31_xsys_core_173;
  wire popcount31_xsys_core_176;
  wire popcount31_xsys_core_179;
  wire popcount31_xsys_core_180;
  wire popcount31_xsys_core_182;
  wire popcount31_xsys_core_183;
  wire popcount31_xsys_core_184;
  wire popcount31_xsys_core_185;
  wire popcount31_xsys_core_186;
  wire popcount31_xsys_core_187;
  wire popcount31_xsys_core_188;
  wire popcount31_xsys_core_190;
  wire popcount31_xsys_core_192;
  wire popcount31_xsys_core_193;
  wire popcount31_xsys_core_194;
  wire popcount31_xsys_core_195;
  wire popcount31_xsys_core_196;
  wire popcount31_xsys_core_197;
  wire popcount31_xsys_core_198;
  wire popcount31_xsys_core_199;
  wire popcount31_xsys_core_200;
  wire popcount31_xsys_core_201;
  wire popcount31_xsys_core_202;
  wire popcount31_xsys_core_206;
  wire popcount31_xsys_core_208;
  wire popcount31_xsys_core_211;
  wire popcount31_xsys_core_212;
  wire popcount31_xsys_core_213;
  wire popcount31_xsys_core_214_not;
  wire popcount31_xsys_core_215;
  wire popcount31_xsys_core_216;
  wire popcount31_xsys_core_218;

  assign popcount31_xsys_core_036 = input_a[26] & input_a[14];
  assign popcount31_xsys_core_038_not = ~input_a[28];
  assign popcount31_xsys_core_039 = ~(input_a[15] & input_a[23]);
  assign popcount31_xsys_core_040 = input_a[19] & input_a[5];
  assign popcount31_xsys_core_041 = ~(input_a[12] & input_a[10]);
  assign popcount31_xsys_core_042 = ~input_a[2];
  assign popcount31_xsys_core_043 = ~(input_a[20] ^ input_a[15]);
  assign popcount31_xsys_core_044 = ~input_a[12];
  assign popcount31_xsys_core_045 = ~(input_a[3] & input_a[22]);
  assign popcount31_xsys_core_047 = ~(input_a[15] & input_a[23]);
  assign popcount31_xsys_core_048 = ~input_a[16];
  assign popcount31_xsys_core_049 = ~(input_a[29] | input_a[25]);
  assign popcount31_xsys_core_050 = ~(input_a[6] ^ input_a[29]);
  assign popcount31_xsys_core_051 = ~(input_a[28] & input_a[26]);
  assign popcount31_xsys_core_052 = ~(input_a[2] & input_a[1]);
  assign popcount31_xsys_core_053 = input_a[2] | input_a[5];
  assign popcount31_xsys_core_057 = input_a[1] & input_a[21];
  assign popcount31_xsys_core_058 = ~(input_a[23] & input_a[2]);
  assign popcount31_xsys_core_060 = input_a[3] | input_a[7];
  assign popcount31_xsys_core_062 = input_a[25] ^ input_a[29];
  assign popcount31_xsys_core_063 = input_a[17] & input_a[2];
  assign popcount31_xsys_core_064 = input_a[27] & input_a[7];
  assign popcount31_xsys_core_065 = input_a[21] & input_a[4];
  assign popcount31_xsys_core_066 = input_a[16] & input_a[29];
  assign popcount31_xsys_core_067 = ~input_a[28];
  assign popcount31_xsys_core_068 = ~(input_a[9] | input_a[22]);
  assign popcount31_xsys_core_072 = ~(input_a[2] ^ input_a[3]);
  assign popcount31_xsys_core_073 = ~(input_a[20] ^ input_a[26]);
  assign popcount31_xsys_core_075 = ~input_a[8];
  assign popcount31_xsys_core_076 = ~(input_a[16] & input_a[27]);
  assign popcount31_xsys_core_078 = ~(input_a[9] & input_a[0]);
  assign popcount31_xsys_core_079 = ~(input_a[4] ^ input_a[4]);
  assign popcount31_xsys_core_080 = ~input_a[14];
  assign popcount31_xsys_core_081_not = ~input_a[6];
  assign popcount31_xsys_core_082 = ~(input_a[23] & input_a[15]);
  assign popcount31_xsys_core_085 = ~input_a[6];
  assign popcount31_xsys_core_088 = ~(input_a[13] & input_a[2]);
  assign popcount31_xsys_core_091 = ~(input_a[24] & input_a[13]);
  assign popcount31_xsys_core_092 = input_a[25] ^ input_a[28];
  assign popcount31_xsys_core_095 = input_a[6] & input_a[11];
  assign popcount31_xsys_core_097 = ~(input_a[28] ^ input_a[9]);
  assign popcount31_xsys_core_098 = input_a[3] | input_a[1];
  assign popcount31_xsys_core_099 = ~(input_a[27] & input_a[28]);
  assign popcount31_xsys_core_101 = input_a[29] | input_a[15];
  assign popcount31_xsys_core_102 = input_a[26] ^ input_a[22];
  assign popcount31_xsys_core_103 = input_a[10] ^ input_a[18];
  assign popcount31_xsys_core_104 = ~(input_a[19] ^ input_a[0]);
  assign popcount31_xsys_core_105 = ~(input_a[11] | input_a[20]);
  assign popcount31_xsys_core_106 = input_a[14] ^ input_a[30];
  assign popcount31_xsys_core_107 = ~input_a[19];
  assign popcount31_xsys_core_108 = input_a[1] | input_a[2];
  assign popcount31_xsys_core_109 = input_a[5] & input_a[16];
  assign popcount31_xsys_core_111 = ~input_a[9];
  assign popcount31_xsys_core_113 = ~(input_a[10] | input_a[17]);
  assign popcount31_xsys_core_114 = input_a[22] ^ input_a[24];
  assign popcount31_xsys_core_117 = input_a[8] & input_a[28];
  assign popcount31_xsys_core_119 = ~(input_a[6] & input_a[22]);
  assign popcount31_xsys_core_120 = input_a[2] & input_a[23];
  assign popcount31_xsys_core_121 = input_a[19] & input_a[25];
  assign popcount31_xsys_core_124 = ~(input_a[7] ^ input_a[27]);
  assign popcount31_xsys_core_127 = input_a[4] & input_a[4];
  assign popcount31_xsys_core_129 = input_a[16] | input_a[17];
  assign popcount31_xsys_core_133 = input_a[11] | input_a[17];
  assign popcount31_xsys_core_135 = input_a[11] | input_a[5];
  assign popcount31_xsys_core_136 = input_a[7] ^ input_a[13];
  assign popcount31_xsys_core_138 = ~input_a[12];
  assign popcount31_xsys_core_140 = ~(input_a[29] & input_a[1]);
  assign popcount31_xsys_core_142 = input_a[27] ^ input_a[28];
  assign popcount31_xsys_core_143 = ~(input_a[1] | input_a[28]);
  assign popcount31_xsys_core_144 = ~input_a[12];
  assign popcount31_xsys_core_145 = input_a[27] & input_a[13];
  assign popcount31_xsys_core_148 = input_a[11] | input_a[15];
  assign popcount31_xsys_core_150 = ~input_a[26];
  assign popcount31_xsys_core_151_not = ~input_a[14];
  assign popcount31_xsys_core_152 = ~(input_a[29] & input_a[22]);
  assign popcount31_xsys_core_153 = ~(input_a[5] | input_a[16]);
  assign popcount31_xsys_core_154 = ~(input_a[23] ^ input_a[5]);
  assign popcount31_xsys_core_155 = ~input_a[11];
  assign popcount31_xsys_core_156 = ~(input_a[17] ^ input_a[8]);
  assign popcount31_xsys_core_158 = ~(input_a[19] ^ input_a[14]);
  assign popcount31_xsys_core_159 = ~(input_a[21] | input_a[6]);
  assign popcount31_xsys_core_160 = input_a[26] ^ input_a[23];
  assign popcount31_xsys_core_161 = ~(input_a[21] | input_a[25]);
  assign popcount31_xsys_core_162 = ~(input_a[6] & input_a[5]);
  assign popcount31_xsys_core_163 = input_a[24] & input_a[24];
  assign popcount31_xsys_core_166 = input_a[17] ^ input_a[2];
  assign popcount31_xsys_core_167 = ~(input_a[23] & input_a[21]);
  assign popcount31_xsys_core_168 = ~(input_a[7] & input_a[11]);
  assign popcount31_xsys_core_169 = ~(input_a[29] & input_a[21]);
  assign popcount31_xsys_core_171 = ~(input_a[25] | input_a[23]);
  assign popcount31_xsys_core_172 = ~(input_a[30] ^ input_a[10]);
  assign popcount31_xsys_core_173 = ~input_a[23];
  assign popcount31_xsys_core_176 = input_a[23] | input_a[25];
  assign popcount31_xsys_core_179 = input_a[27] & input_a[3];
  assign popcount31_xsys_core_180 = ~input_a[19];
  assign popcount31_xsys_core_182 = input_a[3] ^ input_a[21];
  assign popcount31_xsys_core_183 = input_a[15] & input_a[16];
  assign popcount31_xsys_core_184 = ~(input_a[10] | input_a[5]);
  assign popcount31_xsys_core_185 = input_a[11] ^ input_a[2];
  assign popcount31_xsys_core_186 = input_a[22] & input_a[1];
  assign popcount31_xsys_core_187 = ~(input_a[1] & input_a[10]);
  assign popcount31_xsys_core_188 = input_a[29] | input_a[12];
  assign popcount31_xsys_core_190 = input_a[21] ^ input_a[21];
  assign popcount31_xsys_core_192 = ~(input_a[1] & input_a[14]);
  assign popcount31_xsys_core_193 = ~(input_a[0] & input_a[8]);
  assign popcount31_xsys_core_194 = ~(input_a[21] ^ input_a[6]);
  assign popcount31_xsys_core_195 = input_a[3] ^ input_a[7];
  assign popcount31_xsys_core_196 = ~(input_a[30] & input_a[12]);
  assign popcount31_xsys_core_197 = ~input_a[20];
  assign popcount31_xsys_core_198 = ~input_a[28];
  assign popcount31_xsys_core_199 = ~(input_a[30] ^ input_a[22]);
  assign popcount31_xsys_core_200 = ~(input_a[29] | input_a[2]);
  assign popcount31_xsys_core_201 = input_a[1] & input_a[18];
  assign popcount31_xsys_core_202 = ~(input_a[4] | input_a[30]);
  assign popcount31_xsys_core_206 = input_a[21] & input_a[24];
  assign popcount31_xsys_core_208 = ~(input_a[21] | input_a[19]);
  assign popcount31_xsys_core_211 = input_a[17] ^ input_a[9];
  assign popcount31_xsys_core_212 = ~(input_a[15] & input_a[7]);
  assign popcount31_xsys_core_213 = ~(input_a[15] | input_a[4]);
  assign popcount31_xsys_core_214_not = ~input_a[10];
  assign popcount31_xsys_core_215 = input_a[14] ^ input_a[6];
  assign popcount31_xsys_core_216 = ~(input_a[6] & input_a[15]);
  assign popcount31_xsys_core_218 = ~(input_a[0] | input_a[15]);

  assign popcount31_xsys_out[0] = input_a[11];
  assign popcount31_xsys_out[1] = 1'b0;
  assign popcount31_xsys_out[2] = 1'b0;
  assign popcount31_xsys_out[3] = 1'b0;
  assign popcount31_xsys_out[4] = 1'b1;
endmodule