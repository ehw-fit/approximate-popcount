// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.58084
// WCE=18.0
// EP=0.879259%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_ysq8(input [32:0] input_a, output [5:0] popcount33_ysq8_out);
  wire popcount33_ysq8_core_035;
  wire popcount33_ysq8_core_036;
  wire popcount33_ysq8_core_040;
  wire popcount33_ysq8_core_041;
  wire popcount33_ysq8_core_044;
  wire popcount33_ysq8_core_046;
  wire popcount33_ysq8_core_047;
  wire popcount33_ysq8_core_048;
  wire popcount33_ysq8_core_051;
  wire popcount33_ysq8_core_052;
  wire popcount33_ysq8_core_055;
  wire popcount33_ysq8_core_056;
  wire popcount33_ysq8_core_057;
  wire popcount33_ysq8_core_058;
  wire popcount33_ysq8_core_059;
  wire popcount33_ysq8_core_061;
  wire popcount33_ysq8_core_064;
  wire popcount33_ysq8_core_065;
  wire popcount33_ysq8_core_066;
  wire popcount33_ysq8_core_068;
  wire popcount33_ysq8_core_069;
  wire popcount33_ysq8_core_070;
  wire popcount33_ysq8_core_076;
  wire popcount33_ysq8_core_079;
  wire popcount33_ysq8_core_080;
  wire popcount33_ysq8_core_081;
  wire popcount33_ysq8_core_083;
  wire popcount33_ysq8_core_084;
  wire popcount33_ysq8_core_087;
  wire popcount33_ysq8_core_088;
  wire popcount33_ysq8_core_089;
  wire popcount33_ysq8_core_090;
  wire popcount33_ysq8_core_091;
  wire popcount33_ysq8_core_092;
  wire popcount33_ysq8_core_094;
  wire popcount33_ysq8_core_096;
  wire popcount33_ysq8_core_097;
  wire popcount33_ysq8_core_098;
  wire popcount33_ysq8_core_099;
  wire popcount33_ysq8_core_102;
  wire popcount33_ysq8_core_103;
  wire popcount33_ysq8_core_105;
  wire popcount33_ysq8_core_108;
  wire popcount33_ysq8_core_109;
  wire popcount33_ysq8_core_111_not;
  wire popcount33_ysq8_core_112;
  wire popcount33_ysq8_core_113;
  wire popcount33_ysq8_core_115;
  wire popcount33_ysq8_core_117;
  wire popcount33_ysq8_core_118;
  wire popcount33_ysq8_core_119;
  wire popcount33_ysq8_core_121;
  wire popcount33_ysq8_core_123;
  wire popcount33_ysq8_core_125;
  wire popcount33_ysq8_core_126;
  wire popcount33_ysq8_core_128;
  wire popcount33_ysq8_core_130;
  wire popcount33_ysq8_core_132;
  wire popcount33_ysq8_core_133;
  wire popcount33_ysq8_core_134_not;
  wire popcount33_ysq8_core_142;
  wire popcount33_ysq8_core_143_not;
  wire popcount33_ysq8_core_144;
  wire popcount33_ysq8_core_145;
  wire popcount33_ysq8_core_146;
  wire popcount33_ysq8_core_147;
  wire popcount33_ysq8_core_148;
  wire popcount33_ysq8_core_152;
  wire popcount33_ysq8_core_155;
  wire popcount33_ysq8_core_156;
  wire popcount33_ysq8_core_157;
  wire popcount33_ysq8_core_158;
  wire popcount33_ysq8_core_159;
  wire popcount33_ysq8_core_160;
  wire popcount33_ysq8_core_162;
  wire popcount33_ysq8_core_163;
  wire popcount33_ysq8_core_164;
  wire popcount33_ysq8_core_165;
  wire popcount33_ysq8_core_166;
  wire popcount33_ysq8_core_167;
  wire popcount33_ysq8_core_168;
  wire popcount33_ysq8_core_169;
  wire popcount33_ysq8_core_172;
  wire popcount33_ysq8_core_173;
  wire popcount33_ysq8_core_175;
  wire popcount33_ysq8_core_176;
  wire popcount33_ysq8_core_177;
  wire popcount33_ysq8_core_179;
  wire popcount33_ysq8_core_180;
  wire popcount33_ysq8_core_182;
  wire popcount33_ysq8_core_183;
  wire popcount33_ysq8_core_185;
  wire popcount33_ysq8_core_186;
  wire popcount33_ysq8_core_187;
  wire popcount33_ysq8_core_188;
  wire popcount33_ysq8_core_190;
  wire popcount33_ysq8_core_192;
  wire popcount33_ysq8_core_194;
  wire popcount33_ysq8_core_195;
  wire popcount33_ysq8_core_196;
  wire popcount33_ysq8_core_197;
  wire popcount33_ysq8_core_198;
  wire popcount33_ysq8_core_200;
  wire popcount33_ysq8_core_202;
  wire popcount33_ysq8_core_203;
  wire popcount33_ysq8_core_204;
  wire popcount33_ysq8_core_206;
  wire popcount33_ysq8_core_212;
  wire popcount33_ysq8_core_216;
  wire popcount33_ysq8_core_217;
  wire popcount33_ysq8_core_218;
  wire popcount33_ysq8_core_219;
  wire popcount33_ysq8_core_220;
  wire popcount33_ysq8_core_221;
  wire popcount33_ysq8_core_222;
  wire popcount33_ysq8_core_224;
  wire popcount33_ysq8_core_228;
  wire popcount33_ysq8_core_230;
  wire popcount33_ysq8_core_231;
  wire popcount33_ysq8_core_232;
  wire popcount33_ysq8_core_234;
  wire popcount33_ysq8_core_235;
  wire popcount33_ysq8_core_237;
  wire popcount33_ysq8_core_238;

  assign popcount33_ysq8_core_035 = ~input_a[15];
  assign popcount33_ysq8_core_036 = input_a[24] ^ input_a[12];
  assign popcount33_ysq8_core_040 = input_a[23] | input_a[9];
  assign popcount33_ysq8_core_041 = ~(input_a[14] | input_a[10]);
  assign popcount33_ysq8_core_044 = ~(input_a[7] & input_a[32]);
  assign popcount33_ysq8_core_046 = ~(input_a[14] | input_a[16]);
  assign popcount33_ysq8_core_047 = input_a[1] | input_a[13];
  assign popcount33_ysq8_core_048 = ~input_a[5];
  assign popcount33_ysq8_core_051 = ~(input_a[17] | input_a[8]);
  assign popcount33_ysq8_core_052 = ~(input_a[1] & input_a[22]);
  assign popcount33_ysq8_core_055 = ~(input_a[2] | input_a[22]);
  assign popcount33_ysq8_core_056 = ~(input_a[13] & input_a[18]);
  assign popcount33_ysq8_core_057 = ~(input_a[27] & input_a[26]);
  assign popcount33_ysq8_core_058 = ~(input_a[17] ^ input_a[6]);
  assign popcount33_ysq8_core_059 = ~input_a[17];
  assign popcount33_ysq8_core_061 = input_a[8] ^ input_a[9];
  assign popcount33_ysq8_core_064 = ~input_a[28];
  assign popcount33_ysq8_core_065 = ~input_a[3];
  assign popcount33_ysq8_core_066 = input_a[3] & input_a[21];
  assign popcount33_ysq8_core_068 = ~(input_a[2] | input_a[8]);
  assign popcount33_ysq8_core_069 = ~(input_a[26] & input_a[17]);
  assign popcount33_ysq8_core_070 = ~(input_a[4] & input_a[25]);
  assign popcount33_ysq8_core_076 = input_a[20] & input_a[11];
  assign popcount33_ysq8_core_079 = ~input_a[24];
  assign popcount33_ysq8_core_080 = input_a[27] | input_a[32];
  assign popcount33_ysq8_core_081 = ~(input_a[31] ^ input_a[19]);
  assign popcount33_ysq8_core_083 = ~(input_a[18] ^ input_a[31]);
  assign popcount33_ysq8_core_084 = input_a[23] | input_a[27];
  assign popcount33_ysq8_core_087 = input_a[12] & input_a[24];
  assign popcount33_ysq8_core_088 = input_a[30] | input_a[29];
  assign popcount33_ysq8_core_089 = input_a[21] | input_a[4];
  assign popcount33_ysq8_core_090 = ~(input_a[3] | input_a[7]);
  assign popcount33_ysq8_core_091 = ~(input_a[6] | input_a[25]);
  assign popcount33_ysq8_core_092 = input_a[2] | input_a[2];
  assign popcount33_ysq8_core_094 = ~(input_a[18] ^ input_a[21]);
  assign popcount33_ysq8_core_096 = input_a[4] | input_a[32];
  assign popcount33_ysq8_core_097 = ~input_a[30];
  assign popcount33_ysq8_core_098 = ~(input_a[0] | input_a[7]);
  assign popcount33_ysq8_core_099 = input_a[15] | input_a[2];
  assign popcount33_ysq8_core_102 = input_a[9] ^ input_a[4];
  assign popcount33_ysq8_core_103 = ~input_a[30];
  assign popcount33_ysq8_core_105 = input_a[8] & input_a[4];
  assign popcount33_ysq8_core_108 = input_a[19] | input_a[30];
  assign popcount33_ysq8_core_109 = ~(input_a[27] ^ input_a[31]);
  assign popcount33_ysq8_core_111_not = ~input_a[16];
  assign popcount33_ysq8_core_112 = input_a[6] ^ input_a[26];
  assign popcount33_ysq8_core_113 = input_a[5] & input_a[7];
  assign popcount33_ysq8_core_115 = ~input_a[8];
  assign popcount33_ysq8_core_117 = ~(input_a[27] & input_a[19]);
  assign popcount33_ysq8_core_118 = input_a[7] & input_a[16];
  assign popcount33_ysq8_core_119 = ~(input_a[25] ^ input_a[2]);
  assign popcount33_ysq8_core_121 = input_a[23] & input_a[31];
  assign popcount33_ysq8_core_123 = ~(input_a[4] & input_a[11]);
  assign popcount33_ysq8_core_125 = ~input_a[27];
  assign popcount33_ysq8_core_126 = input_a[17] | input_a[12];
  assign popcount33_ysq8_core_128 = ~(input_a[9] & input_a[7]);
  assign popcount33_ysq8_core_130 = input_a[3] & input_a[8];
  assign popcount33_ysq8_core_132 = ~input_a[28];
  assign popcount33_ysq8_core_133 = input_a[30] ^ input_a[17];
  assign popcount33_ysq8_core_134_not = ~input_a[22];
  assign popcount33_ysq8_core_142 = ~(input_a[22] & input_a[31]);
  assign popcount33_ysq8_core_143_not = ~input_a[1];
  assign popcount33_ysq8_core_144 = ~input_a[14];
  assign popcount33_ysq8_core_145 = input_a[30] ^ input_a[3];
  assign popcount33_ysq8_core_146 = input_a[20] ^ input_a[15];
  assign popcount33_ysq8_core_147 = input_a[4] ^ input_a[13];
  assign popcount33_ysq8_core_148 = input_a[9] ^ input_a[1];
  assign popcount33_ysq8_core_152 = input_a[17] | input_a[1];
  assign popcount33_ysq8_core_155 = input_a[11] & input_a[8];
  assign popcount33_ysq8_core_156 = ~(input_a[29] & input_a[10]);
  assign popcount33_ysq8_core_157 = ~(input_a[14] ^ input_a[26]);
  assign popcount33_ysq8_core_158 = ~(input_a[3] ^ input_a[8]);
  assign popcount33_ysq8_core_159 = input_a[15] | input_a[28];
  assign popcount33_ysq8_core_160 = ~(input_a[11] ^ input_a[27]);
  assign popcount33_ysq8_core_162 = ~(input_a[21] | input_a[20]);
  assign popcount33_ysq8_core_163 = ~(input_a[29] & input_a[16]);
  assign popcount33_ysq8_core_164 = ~input_a[0];
  assign popcount33_ysq8_core_165 = input_a[6] & input_a[31];
  assign popcount33_ysq8_core_166 = input_a[26] & input_a[22];
  assign popcount33_ysq8_core_167 = input_a[20] | input_a[3];
  assign popcount33_ysq8_core_168 = ~(input_a[11] | input_a[13]);
  assign popcount33_ysq8_core_169 = input_a[25] ^ input_a[28];
  assign popcount33_ysq8_core_172 = input_a[2] & input_a[8];
  assign popcount33_ysq8_core_173 = ~(input_a[1] & input_a[8]);
  assign popcount33_ysq8_core_175 = ~(input_a[17] ^ input_a[30]);
  assign popcount33_ysq8_core_176 = ~input_a[0];
  assign popcount33_ysq8_core_177 = ~input_a[31];
  assign popcount33_ysq8_core_179 = ~input_a[9];
  assign popcount33_ysq8_core_180 = input_a[31] & input_a[31];
  assign popcount33_ysq8_core_182 = input_a[32] | input_a[0];
  assign popcount33_ysq8_core_183 = input_a[9] & input_a[17];
  assign popcount33_ysq8_core_185 = input_a[6] | input_a[15];
  assign popcount33_ysq8_core_186 = ~(input_a[16] & input_a[2]);
  assign popcount33_ysq8_core_187 = ~(input_a[30] | input_a[29]);
  assign popcount33_ysq8_core_188 = input_a[11] | input_a[21];
  assign popcount33_ysq8_core_190 = input_a[23] | input_a[17];
  assign popcount33_ysq8_core_192 = ~(input_a[12] ^ input_a[1]);
  assign popcount33_ysq8_core_194 = input_a[21] & input_a[17];
  assign popcount33_ysq8_core_195 = ~(input_a[25] ^ input_a[15]);
  assign popcount33_ysq8_core_196 = ~(input_a[24] & input_a[25]);
  assign popcount33_ysq8_core_197 = input_a[31] | input_a[3];
  assign popcount33_ysq8_core_198 = input_a[20] & input_a[8];
  assign popcount33_ysq8_core_200 = ~(input_a[19] & input_a[10]);
  assign popcount33_ysq8_core_202 = ~input_a[6];
  assign popcount33_ysq8_core_203 = ~(input_a[14] ^ input_a[1]);
  assign popcount33_ysq8_core_204 = ~(input_a[26] | input_a[25]);
  assign popcount33_ysq8_core_206 = ~(input_a[25] & input_a[2]);
  assign popcount33_ysq8_core_212 = ~input_a[16];
  assign popcount33_ysq8_core_216 = ~(input_a[24] & input_a[13]);
  assign popcount33_ysq8_core_217 = ~input_a[31];
  assign popcount33_ysq8_core_218 = ~(input_a[27] & input_a[24]);
  assign popcount33_ysq8_core_219 = ~(input_a[26] ^ input_a[25]);
  assign popcount33_ysq8_core_220 = ~(input_a[6] | input_a[4]);
  assign popcount33_ysq8_core_221 = ~input_a[27];
  assign popcount33_ysq8_core_222 = input_a[12] | input_a[15];
  assign popcount33_ysq8_core_224 = input_a[21] & input_a[5];
  assign popcount33_ysq8_core_228 = ~(input_a[23] | input_a[7]);
  assign popcount33_ysq8_core_230 = input_a[30] ^ input_a[27];
  assign popcount33_ysq8_core_231 = input_a[19] ^ input_a[16];
  assign popcount33_ysq8_core_232 = ~(input_a[4] | input_a[6]);
  assign popcount33_ysq8_core_234 = input_a[20] ^ input_a[7];
  assign popcount33_ysq8_core_235 = input_a[5] & input_a[7];
  assign popcount33_ysq8_core_237 = input_a[29] & input_a[24];
  assign popcount33_ysq8_core_238 = input_a[13] | input_a[15];

  assign popcount33_ysq8_out[0] = 1'b0;
  assign popcount33_ysq8_out[1] = 1'b1;
  assign popcount33_ysq8_out[2] = 1'b0;
  assign popcount33_ysq8_out[3] = 1'b0;
  assign popcount33_ysq8_out[4] = 1'b1;
  assign popcount33_ysq8_out[5] = 1'b0;
endmodule