// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=16.5806
// WCE=50.0
// EP=0.972395%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_im4v(input [34:0] input_a, output [5:0] popcount35_im4v_out);
  wire popcount35_im4v_core_037;
  wire popcount35_im4v_core_039;
  wire popcount35_im4v_core_041;
  wire popcount35_im4v_core_043;
  wire popcount35_im4v_core_045;
  wire popcount35_im4v_core_048;
  wire popcount35_im4v_core_049;
  wire popcount35_im4v_core_050;
  wire popcount35_im4v_core_051;
  wire popcount35_im4v_core_052;
  wire popcount35_im4v_core_054;
  wire popcount35_im4v_core_057;
  wire popcount35_im4v_core_059;
  wire popcount35_im4v_core_060;
  wire popcount35_im4v_core_062;
  wire popcount35_im4v_core_066;
  wire popcount35_im4v_core_068;
  wire popcount35_im4v_core_071;
  wire popcount35_im4v_core_072;
  wire popcount35_im4v_core_073;
  wire popcount35_im4v_core_075;
  wire popcount35_im4v_core_076;
  wire popcount35_im4v_core_077;
  wire popcount35_im4v_core_078;
  wire popcount35_im4v_core_079;
  wire popcount35_im4v_core_081;
  wire popcount35_im4v_core_082;
  wire popcount35_im4v_core_083_not;
  wire popcount35_im4v_core_086;
  wire popcount35_im4v_core_087;
  wire popcount35_im4v_core_088;
  wire popcount35_im4v_core_091;
  wire popcount35_im4v_core_092;
  wire popcount35_im4v_core_093;
  wire popcount35_im4v_core_095;
  wire popcount35_im4v_core_096;
  wire popcount35_im4v_core_098;
  wire popcount35_im4v_core_100;
  wire popcount35_im4v_core_102;
  wire popcount35_im4v_core_103;
  wire popcount35_im4v_core_104;
  wire popcount35_im4v_core_107;
  wire popcount35_im4v_core_108;
  wire popcount35_im4v_core_109;
  wire popcount35_im4v_core_111;
  wire popcount35_im4v_core_112;
  wire popcount35_im4v_core_113;
  wire popcount35_im4v_core_114;
  wire popcount35_im4v_core_115;
  wire popcount35_im4v_core_116;
  wire popcount35_im4v_core_118;
  wire popcount35_im4v_core_121;
  wire popcount35_im4v_core_123;
  wire popcount35_im4v_core_125;
  wire popcount35_im4v_core_127;
  wire popcount35_im4v_core_129;
  wire popcount35_im4v_core_130;
  wire popcount35_im4v_core_131;
  wire popcount35_im4v_core_132;
  wire popcount35_im4v_core_133;
  wire popcount35_im4v_core_134;
  wire popcount35_im4v_core_135;
  wire popcount35_im4v_core_136;
  wire popcount35_im4v_core_137;
  wire popcount35_im4v_core_138;
  wire popcount35_im4v_core_139;
  wire popcount35_im4v_core_140;
  wire popcount35_im4v_core_141;
  wire popcount35_im4v_core_142;
  wire popcount35_im4v_core_143;
  wire popcount35_im4v_core_145;
  wire popcount35_im4v_core_146;
  wire popcount35_im4v_core_148;
  wire popcount35_im4v_core_150;
  wire popcount35_im4v_core_151;
  wire popcount35_im4v_core_154;
  wire popcount35_im4v_core_155;
  wire popcount35_im4v_core_158;
  wire popcount35_im4v_core_159;
  wire popcount35_im4v_core_160;
  wire popcount35_im4v_core_162;
  wire popcount35_im4v_core_163;
  wire popcount35_im4v_core_164;
  wire popcount35_im4v_core_165;
  wire popcount35_im4v_core_166;
  wire popcount35_im4v_core_167;
  wire popcount35_im4v_core_168;
  wire popcount35_im4v_core_170;
  wire popcount35_im4v_core_171;
  wire popcount35_im4v_core_174;
  wire popcount35_im4v_core_176;
  wire popcount35_im4v_core_177;
  wire popcount35_im4v_core_180;
  wire popcount35_im4v_core_181;
  wire popcount35_im4v_core_182;
  wire popcount35_im4v_core_183;
  wire popcount35_im4v_core_184;
  wire popcount35_im4v_core_186;
  wire popcount35_im4v_core_187;
  wire popcount35_im4v_core_188;
  wire popcount35_im4v_core_189;
  wire popcount35_im4v_core_190;
  wire popcount35_im4v_core_192;
  wire popcount35_im4v_core_193;
  wire popcount35_im4v_core_194;
  wire popcount35_im4v_core_195;
  wire popcount35_im4v_core_197;
  wire popcount35_im4v_core_198;
  wire popcount35_im4v_core_199;
  wire popcount35_im4v_core_201;
  wire popcount35_im4v_core_204;
  wire popcount35_im4v_core_206;
  wire popcount35_im4v_core_211;
  wire popcount35_im4v_core_212_not;
  wire popcount35_im4v_core_213;
  wire popcount35_im4v_core_214;
  wire popcount35_im4v_core_215;
  wire popcount35_im4v_core_216;
  wire popcount35_im4v_core_219;
  wire popcount35_im4v_core_222;
  wire popcount35_im4v_core_223;
  wire popcount35_im4v_core_224;
  wire popcount35_im4v_core_225_not;
  wire popcount35_im4v_core_226;
  wire popcount35_im4v_core_227;
  wire popcount35_im4v_core_228;
  wire popcount35_im4v_core_230;
  wire popcount35_im4v_core_231;
  wire popcount35_im4v_core_232;
  wire popcount35_im4v_core_233;
  wire popcount35_im4v_core_234;
  wire popcount35_im4v_core_237;
  wire popcount35_im4v_core_238;
  wire popcount35_im4v_core_239;
  wire popcount35_im4v_core_243;
  wire popcount35_im4v_core_245_not;
  wire popcount35_im4v_core_246;
  wire popcount35_im4v_core_247;
  wire popcount35_im4v_core_248;
  wire popcount35_im4v_core_249;
  wire popcount35_im4v_core_251;
  wire popcount35_im4v_core_252;
  wire popcount35_im4v_core_260;
  wire popcount35_im4v_core_261;
  wire popcount35_im4v_core_262;
  wire popcount35_im4v_core_263;
  wire popcount35_im4v_core_264;

  assign popcount35_im4v_core_037 = input_a[2] | input_a[30];
  assign popcount35_im4v_core_039 = input_a[20] & input_a[12];
  assign popcount35_im4v_core_041 = input_a[14] & input_a[16];
  assign popcount35_im4v_core_043 = ~(input_a[2] | input_a[9]);
  assign popcount35_im4v_core_045 = ~(input_a[32] ^ input_a[5]);
  assign popcount35_im4v_core_048 = input_a[18] & input_a[0];
  assign popcount35_im4v_core_049 = ~input_a[22];
  assign popcount35_im4v_core_050 = ~(input_a[12] | input_a[14]);
  assign popcount35_im4v_core_051 = ~(input_a[23] & input_a[6]);
  assign popcount35_im4v_core_052 = ~(input_a[17] & input_a[30]);
  assign popcount35_im4v_core_054 = ~(input_a[2] & input_a[12]);
  assign popcount35_im4v_core_057 = input_a[31] | input_a[6];
  assign popcount35_im4v_core_059 = input_a[0] ^ input_a[23];
  assign popcount35_im4v_core_060 = input_a[32] & input_a[1];
  assign popcount35_im4v_core_062 = input_a[18] & input_a[18];
  assign popcount35_im4v_core_066 = input_a[30] | input_a[34];
  assign popcount35_im4v_core_068 = ~(input_a[0] & input_a[34]);
  assign popcount35_im4v_core_071 = ~input_a[17];
  assign popcount35_im4v_core_072 = ~(input_a[13] & input_a[9]);
  assign popcount35_im4v_core_073 = ~(input_a[4] ^ input_a[1]);
  assign popcount35_im4v_core_075 = ~(input_a[31] ^ input_a[0]);
  assign popcount35_im4v_core_076 = ~(input_a[3] & input_a[0]);
  assign popcount35_im4v_core_077 = input_a[5] | input_a[10];
  assign popcount35_im4v_core_078 = input_a[1] & input_a[6];
  assign popcount35_im4v_core_079 = input_a[21] ^ input_a[13];
  assign popcount35_im4v_core_081 = ~(input_a[22] ^ input_a[18]);
  assign popcount35_im4v_core_082 = input_a[14] ^ input_a[21];
  assign popcount35_im4v_core_083_not = ~input_a[25];
  assign popcount35_im4v_core_086 = ~(input_a[26] | input_a[4]);
  assign popcount35_im4v_core_087 = ~(input_a[15] | input_a[8]);
  assign popcount35_im4v_core_088 = input_a[30] ^ input_a[28];
  assign popcount35_im4v_core_091 = input_a[28] | input_a[29];
  assign popcount35_im4v_core_092 = ~(input_a[5] | input_a[15]);
  assign popcount35_im4v_core_093 = ~(input_a[10] & input_a[30]);
  assign popcount35_im4v_core_095 = ~(input_a[15] | input_a[18]);
  assign popcount35_im4v_core_096 = ~input_a[0];
  assign popcount35_im4v_core_098 = input_a[13] | input_a[32];
  assign popcount35_im4v_core_100 = input_a[17] ^ input_a[12];
  assign popcount35_im4v_core_102 = input_a[11] ^ input_a[1];
  assign popcount35_im4v_core_103 = input_a[32] | input_a[2];
  assign popcount35_im4v_core_104 = ~(input_a[7] ^ input_a[11]);
  assign popcount35_im4v_core_107 = input_a[18] | input_a[21];
  assign popcount35_im4v_core_108 = ~(input_a[9] | input_a[31]);
  assign popcount35_im4v_core_109 = ~(input_a[5] ^ input_a[19]);
  assign popcount35_im4v_core_111 = ~input_a[10];
  assign popcount35_im4v_core_112 = ~input_a[15];
  assign popcount35_im4v_core_113 = ~(input_a[27] & input_a[17]);
  assign popcount35_im4v_core_114 = ~(input_a[25] ^ input_a[31]);
  assign popcount35_im4v_core_115 = ~input_a[26];
  assign popcount35_im4v_core_116 = input_a[33] & input_a[21];
  assign popcount35_im4v_core_118 = ~(input_a[18] ^ input_a[33]);
  assign popcount35_im4v_core_121 = input_a[21] | input_a[1];
  assign popcount35_im4v_core_123 = ~(input_a[2] | input_a[26]);
  assign popcount35_im4v_core_125 = ~input_a[7];
  assign popcount35_im4v_core_127 = ~(input_a[12] & input_a[33]);
  assign popcount35_im4v_core_129 = input_a[8] | input_a[4];
  assign popcount35_im4v_core_130 = ~(input_a[16] | input_a[11]);
  assign popcount35_im4v_core_131 = input_a[0] & input_a[26];
  assign popcount35_im4v_core_132 = input_a[10] ^ input_a[1];
  assign popcount35_im4v_core_133 = input_a[17] & input_a[11];
  assign popcount35_im4v_core_134 = input_a[12] ^ input_a[12];
  assign popcount35_im4v_core_135 = input_a[31] | input_a[33];
  assign popcount35_im4v_core_136 = ~(input_a[32] ^ input_a[27]);
  assign popcount35_im4v_core_137 = input_a[24] ^ input_a[10];
  assign popcount35_im4v_core_138 = ~(input_a[19] ^ input_a[33]);
  assign popcount35_im4v_core_139 = ~(input_a[23] ^ input_a[26]);
  assign popcount35_im4v_core_140 = input_a[21] ^ input_a[26];
  assign popcount35_im4v_core_141 = ~(input_a[7] | input_a[32]);
  assign popcount35_im4v_core_142 = input_a[34] | input_a[16];
  assign popcount35_im4v_core_143 = ~input_a[2];
  assign popcount35_im4v_core_145 = ~(input_a[22] ^ input_a[17]);
  assign popcount35_im4v_core_146 = ~(input_a[13] | input_a[7]);
  assign popcount35_im4v_core_148 = input_a[10] | input_a[19];
  assign popcount35_im4v_core_150 = ~(input_a[1] & input_a[32]);
  assign popcount35_im4v_core_151 = input_a[7] ^ input_a[30];
  assign popcount35_im4v_core_154 = input_a[0] & input_a[29];
  assign popcount35_im4v_core_155 = input_a[7] ^ input_a[24];
  assign popcount35_im4v_core_158 = input_a[16] ^ input_a[11];
  assign popcount35_im4v_core_159 = ~input_a[29];
  assign popcount35_im4v_core_160 = ~(input_a[28] | input_a[31]);
  assign popcount35_im4v_core_162 = ~(input_a[32] ^ input_a[8]);
  assign popcount35_im4v_core_163 = ~(input_a[3] ^ input_a[28]);
  assign popcount35_im4v_core_164 = ~input_a[19];
  assign popcount35_im4v_core_165 = ~input_a[31];
  assign popcount35_im4v_core_166 = ~(input_a[27] & input_a[1]);
  assign popcount35_im4v_core_167 = ~(input_a[3] & input_a[10]);
  assign popcount35_im4v_core_168 = input_a[31] & input_a[19];
  assign popcount35_im4v_core_170 = ~(input_a[16] ^ input_a[20]);
  assign popcount35_im4v_core_171 = ~(input_a[11] & input_a[13]);
  assign popcount35_im4v_core_174 = input_a[9] | input_a[0];
  assign popcount35_im4v_core_176 = ~(input_a[5] | input_a[5]);
  assign popcount35_im4v_core_177 = input_a[33] | input_a[10];
  assign popcount35_im4v_core_180 = ~(input_a[2] ^ input_a[5]);
  assign popcount35_im4v_core_181 = ~(input_a[22] & input_a[31]);
  assign popcount35_im4v_core_182 = ~input_a[24];
  assign popcount35_im4v_core_183 = ~(input_a[0] & input_a[13]);
  assign popcount35_im4v_core_184 = input_a[25] | input_a[1];
  assign popcount35_im4v_core_186 = ~(input_a[17] ^ input_a[26]);
  assign popcount35_im4v_core_187 = input_a[29] | input_a[27];
  assign popcount35_im4v_core_188 = ~(input_a[9] ^ input_a[29]);
  assign popcount35_im4v_core_189 = ~(input_a[30] & input_a[12]);
  assign popcount35_im4v_core_190 = ~(input_a[19] | input_a[1]);
  assign popcount35_im4v_core_192 = ~(input_a[16] | input_a[19]);
  assign popcount35_im4v_core_193 = ~input_a[3];
  assign popcount35_im4v_core_194 = input_a[32] ^ input_a[2];
  assign popcount35_im4v_core_195 = input_a[31] | input_a[33];
  assign popcount35_im4v_core_197 = ~input_a[18];
  assign popcount35_im4v_core_198 = ~(input_a[33] | input_a[22]);
  assign popcount35_im4v_core_199 = input_a[7] | input_a[11];
  assign popcount35_im4v_core_201 = input_a[27] ^ input_a[11];
  assign popcount35_im4v_core_204 = ~input_a[0];
  assign popcount35_im4v_core_206 = input_a[24] | input_a[22];
  assign popcount35_im4v_core_211 = ~input_a[12];
  assign popcount35_im4v_core_212_not = ~input_a[16];
  assign popcount35_im4v_core_213 = ~(input_a[1] ^ input_a[29]);
  assign popcount35_im4v_core_214 = input_a[18] & input_a[27];
  assign popcount35_im4v_core_215 = ~(input_a[3] & input_a[7]);
  assign popcount35_im4v_core_216 = input_a[11] ^ input_a[4];
  assign popcount35_im4v_core_219 = ~(input_a[0] ^ input_a[1]);
  assign popcount35_im4v_core_222 = input_a[25] ^ input_a[34];
  assign popcount35_im4v_core_223 = ~(input_a[17] | input_a[1]);
  assign popcount35_im4v_core_224 = ~input_a[8];
  assign popcount35_im4v_core_225_not = ~input_a[4];
  assign popcount35_im4v_core_226 = input_a[25] ^ input_a[16];
  assign popcount35_im4v_core_227 = input_a[18] | input_a[11];
  assign popcount35_im4v_core_228 = ~(input_a[30] ^ input_a[4]);
  assign popcount35_im4v_core_230 = ~(input_a[9] | input_a[12]);
  assign popcount35_im4v_core_231 = input_a[31] ^ input_a[8];
  assign popcount35_im4v_core_232 = ~(input_a[3] | input_a[21]);
  assign popcount35_im4v_core_233 = ~(input_a[11] | input_a[5]);
  assign popcount35_im4v_core_234 = ~input_a[2];
  assign popcount35_im4v_core_237 = input_a[27] ^ input_a[28];
  assign popcount35_im4v_core_238 = ~(input_a[2] & input_a[34]);
  assign popcount35_im4v_core_239 = input_a[32] & input_a[29];
  assign popcount35_im4v_core_243 = ~(input_a[23] ^ input_a[28]);
  assign popcount35_im4v_core_245_not = ~input_a[6];
  assign popcount35_im4v_core_246 = input_a[14] & input_a[30];
  assign popcount35_im4v_core_247 = input_a[0] ^ input_a[24];
  assign popcount35_im4v_core_248 = input_a[15] & input_a[18];
  assign popcount35_im4v_core_249 = input_a[18] & input_a[32];
  assign popcount35_im4v_core_251 = ~input_a[8];
  assign popcount35_im4v_core_252 = ~(input_a[7] & input_a[9]);
  assign popcount35_im4v_core_260 = input_a[0] & input_a[13];
  assign popcount35_im4v_core_261 = ~(input_a[29] & input_a[21]);
  assign popcount35_im4v_core_262 = input_a[5] | input_a[2];
  assign popcount35_im4v_core_263 = ~(input_a[8] ^ input_a[4]);
  assign popcount35_im4v_core_264 = ~(input_a[3] | input_a[9]);

  assign popcount35_im4v_out[0] = 1'b0;
  assign popcount35_im4v_out[1] = input_a[28];
  assign popcount35_im4v_out[2] = input_a[21];
  assign popcount35_im4v_out[3] = 1'b0;
  assign popcount35_im4v_out[4] = input_a[23];
  assign popcount35_im4v_out[5] = input_a[24];
endmodule