// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.53964
// WCE=28.0
// EP=0.986587%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_7upc(input [38:0] input_a, output [5:0] popcount39_7upc_out);
  wire popcount39_7upc_core_041;
  wire popcount39_7upc_core_044;
  wire popcount39_7upc_core_046;
  wire popcount39_7upc_core_047;
  wire popcount39_7upc_core_048;
  wire popcount39_7upc_core_049;
  wire popcount39_7upc_core_053;
  wire popcount39_7upc_core_054;
  wire popcount39_7upc_core_055;
  wire popcount39_7upc_core_056;
  wire popcount39_7upc_core_058;
  wire popcount39_7upc_core_059;
  wire popcount39_7upc_core_060;
  wire popcount39_7upc_core_061;
  wire popcount39_7upc_core_063;
  wire popcount39_7upc_core_064;
  wire popcount39_7upc_core_069;
  wire popcount39_7upc_core_071;
  wire popcount39_7upc_core_072;
  wire popcount39_7upc_core_073;
  wire popcount39_7upc_core_074;
  wire popcount39_7upc_core_075;
  wire popcount39_7upc_core_077;
  wire popcount39_7upc_core_079;
  wire popcount39_7upc_core_080;
  wire popcount39_7upc_core_081;
  wire popcount39_7upc_core_082;
  wire popcount39_7upc_core_083;
  wire popcount39_7upc_core_084;
  wire popcount39_7upc_core_085;
  wire popcount39_7upc_core_086;
  wire popcount39_7upc_core_089;
  wire popcount39_7upc_core_090;
  wire popcount39_7upc_core_091;
  wire popcount39_7upc_core_092;
  wire popcount39_7upc_core_095;
  wire popcount39_7upc_core_097;
  wire popcount39_7upc_core_098;
  wire popcount39_7upc_core_099;
  wire popcount39_7upc_core_100;
  wire popcount39_7upc_core_101;
  wire popcount39_7upc_core_105;
  wire popcount39_7upc_core_107;
  wire popcount39_7upc_core_109;
  wire popcount39_7upc_core_110;
  wire popcount39_7upc_core_111;
  wire popcount39_7upc_core_112;
  wire popcount39_7upc_core_114;
  wire popcount39_7upc_core_116;
  wire popcount39_7upc_core_117;
  wire popcount39_7upc_core_121;
  wire popcount39_7upc_core_122;
  wire popcount39_7upc_core_124;
  wire popcount39_7upc_core_125;
  wire popcount39_7upc_core_127;
  wire popcount39_7upc_core_130;
  wire popcount39_7upc_core_132;
  wire popcount39_7upc_core_133;
  wire popcount39_7upc_core_134;
  wire popcount39_7upc_core_136;
  wire popcount39_7upc_core_139;
  wire popcount39_7upc_core_140;
  wire popcount39_7upc_core_141;
  wire popcount39_7upc_core_142;
  wire popcount39_7upc_core_144;
  wire popcount39_7upc_core_145;
  wire popcount39_7upc_core_146;
  wire popcount39_7upc_core_147;
  wire popcount39_7upc_core_148;
  wire popcount39_7upc_core_149;
  wire popcount39_7upc_core_150;
  wire popcount39_7upc_core_151;
  wire popcount39_7upc_core_152;
  wire popcount39_7upc_core_158_not;
  wire popcount39_7upc_core_159;
  wire popcount39_7upc_core_160;
  wire popcount39_7upc_core_161;
  wire popcount39_7upc_core_162;
  wire popcount39_7upc_core_163;
  wire popcount39_7upc_core_164;
  wire popcount39_7upc_core_165;
  wire popcount39_7upc_core_166;
  wire popcount39_7upc_core_167;
  wire popcount39_7upc_core_171;
  wire popcount39_7upc_core_173_not;
  wire popcount39_7upc_core_174;
  wire popcount39_7upc_core_176;
  wire popcount39_7upc_core_180;
  wire popcount39_7upc_core_182;
  wire popcount39_7upc_core_183;
  wire popcount39_7upc_core_184;
  wire popcount39_7upc_core_185;
  wire popcount39_7upc_core_186;
  wire popcount39_7upc_core_187;
  wire popcount39_7upc_core_188;
  wire popcount39_7upc_core_189;
  wire popcount39_7upc_core_190;
  wire popcount39_7upc_core_192;
  wire popcount39_7upc_core_193;
  wire popcount39_7upc_core_194;
  wire popcount39_7upc_core_196;
  wire popcount39_7upc_core_197;
  wire popcount39_7upc_core_198;
  wire popcount39_7upc_core_199;
  wire popcount39_7upc_core_200;
  wire popcount39_7upc_core_202_not;
  wire popcount39_7upc_core_203;
  wire popcount39_7upc_core_205;
  wire popcount39_7upc_core_206;
  wire popcount39_7upc_core_207;
  wire popcount39_7upc_core_208;
  wire popcount39_7upc_core_209;
  wire popcount39_7upc_core_212;
  wire popcount39_7upc_core_213;
  wire popcount39_7upc_core_215;
  wire popcount39_7upc_core_217;
  wire popcount39_7upc_core_218;
  wire popcount39_7upc_core_219;
  wire popcount39_7upc_core_221;
  wire popcount39_7upc_core_223;
  wire popcount39_7upc_core_230_not;
  wire popcount39_7upc_core_232;
  wire popcount39_7upc_core_233;
  wire popcount39_7upc_core_235;
  wire popcount39_7upc_core_236;
  wire popcount39_7upc_core_241;
  wire popcount39_7upc_core_242;
  wire popcount39_7upc_core_243;
  wire popcount39_7upc_core_244;
  wire popcount39_7upc_core_246;
  wire popcount39_7upc_core_247;
  wire popcount39_7upc_core_248;
  wire popcount39_7upc_core_249;
  wire popcount39_7upc_core_250;
  wire popcount39_7upc_core_252;
  wire popcount39_7upc_core_253;
  wire popcount39_7upc_core_254;
  wire popcount39_7upc_core_255;
  wire popcount39_7upc_core_257;
  wire popcount39_7upc_core_258;
  wire popcount39_7upc_core_259;
  wire popcount39_7upc_core_262_not;
  wire popcount39_7upc_core_264;
  wire popcount39_7upc_core_265;
  wire popcount39_7upc_core_266;
  wire popcount39_7upc_core_268;
  wire popcount39_7upc_core_269;
  wire popcount39_7upc_core_273_not;
  wire popcount39_7upc_core_274;
  wire popcount39_7upc_core_276;
  wire popcount39_7upc_core_277;
  wire popcount39_7upc_core_278;
  wire popcount39_7upc_core_279;
  wire popcount39_7upc_core_280;
  wire popcount39_7upc_core_282;
  wire popcount39_7upc_core_284;
  wire popcount39_7upc_core_285;
  wire popcount39_7upc_core_290;
  wire popcount39_7upc_core_295;
  wire popcount39_7upc_core_296;
  wire popcount39_7upc_core_300;
  wire popcount39_7upc_core_302;
  wire popcount39_7upc_core_303;
  wire popcount39_7upc_core_304_not;
  wire popcount39_7upc_core_305;

  assign popcount39_7upc_core_041 = ~(input_a[28] ^ input_a[23]);
  assign popcount39_7upc_core_044 = input_a[2] ^ input_a[12];
  assign popcount39_7upc_core_046 = ~(input_a[34] | input_a[14]);
  assign popcount39_7upc_core_047 = input_a[23] ^ input_a[6];
  assign popcount39_7upc_core_048 = ~(input_a[29] ^ input_a[9]);
  assign popcount39_7upc_core_049 = input_a[34] ^ input_a[29];
  assign popcount39_7upc_core_053 = input_a[29] & input_a[36];
  assign popcount39_7upc_core_054 = input_a[9] | input_a[34];
  assign popcount39_7upc_core_055 = ~(input_a[14] | input_a[11]);
  assign popcount39_7upc_core_056 = ~(input_a[31] ^ input_a[24]);
  assign popcount39_7upc_core_058 = input_a[19] | input_a[27];
  assign popcount39_7upc_core_059 = input_a[11] | input_a[0];
  assign popcount39_7upc_core_060 = input_a[24] & input_a[21];
  assign popcount39_7upc_core_061 = input_a[12] & input_a[6];
  assign popcount39_7upc_core_063 = input_a[0] ^ input_a[12];
  assign popcount39_7upc_core_064 = ~(input_a[30] | input_a[31]);
  assign popcount39_7upc_core_069 = ~(input_a[20] | input_a[32]);
  assign popcount39_7upc_core_071 = input_a[17] ^ input_a[38];
  assign popcount39_7upc_core_072 = ~(input_a[20] & input_a[24]);
  assign popcount39_7upc_core_073 = ~(input_a[9] | input_a[25]);
  assign popcount39_7upc_core_074 = ~input_a[18];
  assign popcount39_7upc_core_075 = input_a[29] | input_a[23];
  assign popcount39_7upc_core_077 = ~input_a[38];
  assign popcount39_7upc_core_079 = ~(input_a[1] | input_a[2]);
  assign popcount39_7upc_core_080 = ~(input_a[9] | input_a[4]);
  assign popcount39_7upc_core_081 = input_a[14] | input_a[19];
  assign popcount39_7upc_core_082 = input_a[25] ^ input_a[35];
  assign popcount39_7upc_core_083 = input_a[15] | input_a[7];
  assign popcount39_7upc_core_084 = ~input_a[14];
  assign popcount39_7upc_core_085 = ~(input_a[27] ^ input_a[31]);
  assign popcount39_7upc_core_086 = input_a[15] ^ input_a[34];
  assign popcount39_7upc_core_089 = ~(input_a[38] | input_a[15]);
  assign popcount39_7upc_core_090 = ~input_a[5];
  assign popcount39_7upc_core_091 = ~(input_a[5] ^ input_a[38]);
  assign popcount39_7upc_core_092 = ~(input_a[27] ^ input_a[30]);
  assign popcount39_7upc_core_095 = input_a[26] ^ input_a[6];
  assign popcount39_7upc_core_097 = ~(input_a[1] & input_a[11]);
  assign popcount39_7upc_core_098 = input_a[13] | input_a[16];
  assign popcount39_7upc_core_099 = ~(input_a[32] & input_a[27]);
  assign popcount39_7upc_core_100 = ~input_a[37];
  assign popcount39_7upc_core_101 = input_a[12] ^ input_a[16];
  assign popcount39_7upc_core_105 = ~(input_a[0] | input_a[8]);
  assign popcount39_7upc_core_107 = ~(input_a[10] | input_a[34]);
  assign popcount39_7upc_core_109 = ~(input_a[33] | input_a[16]);
  assign popcount39_7upc_core_110 = ~(input_a[29] & input_a[30]);
  assign popcount39_7upc_core_111 = ~input_a[34];
  assign popcount39_7upc_core_112 = input_a[28] ^ input_a[27];
  assign popcount39_7upc_core_114 = input_a[19] ^ input_a[18];
  assign popcount39_7upc_core_116 = input_a[15] ^ input_a[17];
  assign popcount39_7upc_core_117 = ~(input_a[32] | input_a[31]);
  assign popcount39_7upc_core_121 = input_a[35] | input_a[18];
  assign popcount39_7upc_core_122 = input_a[10] & input_a[7];
  assign popcount39_7upc_core_124 = ~(input_a[7] ^ input_a[33]);
  assign popcount39_7upc_core_125 = ~(input_a[10] | input_a[6]);
  assign popcount39_7upc_core_127 = ~(input_a[23] ^ input_a[31]);
  assign popcount39_7upc_core_130 = ~input_a[4];
  assign popcount39_7upc_core_132 = ~input_a[21];
  assign popcount39_7upc_core_133 = ~input_a[29];
  assign popcount39_7upc_core_134 = input_a[36] & input_a[38];
  assign popcount39_7upc_core_136 = input_a[10] | input_a[5];
  assign popcount39_7upc_core_139 = ~(input_a[38] & input_a[37]);
  assign popcount39_7upc_core_140 = ~(input_a[6] | input_a[27]);
  assign popcount39_7upc_core_141 = ~(input_a[35] | input_a[5]);
  assign popcount39_7upc_core_142 = ~input_a[20];
  assign popcount39_7upc_core_144 = input_a[14] | input_a[4];
  assign popcount39_7upc_core_145 = input_a[37] & input_a[32];
  assign popcount39_7upc_core_146 = ~(input_a[36] | input_a[33]);
  assign popcount39_7upc_core_147 = ~(input_a[9] & input_a[29]);
  assign popcount39_7upc_core_148 = ~input_a[18];
  assign popcount39_7upc_core_149 = input_a[0] & input_a[16];
  assign popcount39_7upc_core_150 = input_a[34] | input_a[28];
  assign popcount39_7upc_core_151 = ~(input_a[7] & input_a[11]);
  assign popcount39_7upc_core_152 = ~(input_a[3] ^ input_a[36]);
  assign popcount39_7upc_core_158_not = ~input_a[21];
  assign popcount39_7upc_core_159 = ~input_a[7];
  assign popcount39_7upc_core_160 = ~(input_a[32] ^ input_a[3]);
  assign popcount39_7upc_core_161 = input_a[33] ^ input_a[15];
  assign popcount39_7upc_core_162 = input_a[27] & input_a[13];
  assign popcount39_7upc_core_163 = input_a[24] ^ input_a[30];
  assign popcount39_7upc_core_164 = input_a[25] | input_a[23];
  assign popcount39_7upc_core_165 = ~(input_a[17] | input_a[33]);
  assign popcount39_7upc_core_166 = ~input_a[0];
  assign popcount39_7upc_core_167 = ~(input_a[8] & input_a[19]);
  assign popcount39_7upc_core_171 = ~(input_a[25] ^ input_a[26]);
  assign popcount39_7upc_core_173_not = ~input_a[33];
  assign popcount39_7upc_core_174 = ~input_a[9];
  assign popcount39_7upc_core_176 = input_a[33] | input_a[19];
  assign popcount39_7upc_core_180 = ~(input_a[30] | input_a[35]);
  assign popcount39_7upc_core_182 = ~(input_a[15] | input_a[16]);
  assign popcount39_7upc_core_183 = ~(input_a[4] ^ input_a[36]);
  assign popcount39_7upc_core_184 = ~(input_a[3] ^ input_a[0]);
  assign popcount39_7upc_core_185 = ~(input_a[28] & input_a[9]);
  assign popcount39_7upc_core_186 = ~input_a[34];
  assign popcount39_7upc_core_187 = ~(input_a[19] ^ input_a[29]);
  assign popcount39_7upc_core_188 = input_a[33] ^ input_a[21];
  assign popcount39_7upc_core_189 = ~input_a[23];
  assign popcount39_7upc_core_190 = ~(input_a[25] & input_a[4]);
  assign popcount39_7upc_core_192 = input_a[38] ^ input_a[17];
  assign popcount39_7upc_core_193 = input_a[7] ^ input_a[33];
  assign popcount39_7upc_core_194 = ~(input_a[6] & input_a[22]);
  assign popcount39_7upc_core_196 = ~(input_a[17] ^ input_a[7]);
  assign popcount39_7upc_core_197 = ~input_a[4];
  assign popcount39_7upc_core_198 = ~(input_a[3] ^ input_a[17]);
  assign popcount39_7upc_core_199 = ~(input_a[25] | input_a[18]);
  assign popcount39_7upc_core_200 = input_a[36] & input_a[25];
  assign popcount39_7upc_core_202_not = ~input_a[33];
  assign popcount39_7upc_core_203 = input_a[35] & input_a[33];
  assign popcount39_7upc_core_205 = ~(input_a[9] & input_a[24]);
  assign popcount39_7upc_core_206 = ~(input_a[1] & input_a[25]);
  assign popcount39_7upc_core_207 = ~(input_a[12] ^ input_a[23]);
  assign popcount39_7upc_core_208 = input_a[17] | input_a[7];
  assign popcount39_7upc_core_209 = input_a[13] & input_a[18];
  assign popcount39_7upc_core_212 = input_a[34] ^ input_a[26];
  assign popcount39_7upc_core_213 = ~(input_a[3] | input_a[3]);
  assign popcount39_7upc_core_215 = ~input_a[17];
  assign popcount39_7upc_core_217 = input_a[26] | input_a[11];
  assign popcount39_7upc_core_218 = ~(input_a[28] & input_a[2]);
  assign popcount39_7upc_core_219 = ~(input_a[10] & input_a[38]);
  assign popcount39_7upc_core_221 = ~input_a[18];
  assign popcount39_7upc_core_223 = ~(input_a[8] ^ input_a[23]);
  assign popcount39_7upc_core_230_not = ~input_a[23];
  assign popcount39_7upc_core_232 = input_a[12] ^ input_a[6];
  assign popcount39_7upc_core_233 = input_a[20] ^ input_a[28];
  assign popcount39_7upc_core_235 = ~(input_a[0] & input_a[20]);
  assign popcount39_7upc_core_236 = ~input_a[20];
  assign popcount39_7upc_core_241 = input_a[35] | input_a[14];
  assign popcount39_7upc_core_242 = ~input_a[38];
  assign popcount39_7upc_core_243 = input_a[14] | input_a[13];
  assign popcount39_7upc_core_244 = input_a[21] ^ input_a[15];
  assign popcount39_7upc_core_246 = input_a[0] | input_a[36];
  assign popcount39_7upc_core_247 = input_a[4] & input_a[24];
  assign popcount39_7upc_core_248 = input_a[35] ^ input_a[18];
  assign popcount39_7upc_core_249 = ~(input_a[0] ^ input_a[19]);
  assign popcount39_7upc_core_250 = input_a[10] | input_a[1];
  assign popcount39_7upc_core_252 = input_a[5] & input_a[26];
  assign popcount39_7upc_core_253 = ~(input_a[9] ^ input_a[26]);
  assign popcount39_7upc_core_254 = input_a[18] ^ input_a[1];
  assign popcount39_7upc_core_255 = input_a[31] ^ input_a[18];
  assign popcount39_7upc_core_257 = ~(input_a[28] ^ input_a[23]);
  assign popcount39_7upc_core_258 = ~input_a[32];
  assign popcount39_7upc_core_259 = input_a[22] ^ input_a[7];
  assign popcount39_7upc_core_262_not = ~input_a[9];
  assign popcount39_7upc_core_264 = input_a[19] | input_a[5];
  assign popcount39_7upc_core_265 = ~(input_a[8] ^ input_a[28]);
  assign popcount39_7upc_core_266 = ~input_a[25];
  assign popcount39_7upc_core_268 = ~input_a[26];
  assign popcount39_7upc_core_269 = input_a[21] & input_a[3];
  assign popcount39_7upc_core_273_not = ~input_a[36];
  assign popcount39_7upc_core_274 = ~input_a[7];
  assign popcount39_7upc_core_276 = ~(input_a[30] | input_a[25]);
  assign popcount39_7upc_core_277 = ~(input_a[23] | input_a[36]);
  assign popcount39_7upc_core_278 = input_a[2] | input_a[20];
  assign popcount39_7upc_core_279 = input_a[17] | input_a[3];
  assign popcount39_7upc_core_280 = input_a[2] & input_a[12];
  assign popcount39_7upc_core_282 = ~input_a[21];
  assign popcount39_7upc_core_284 = ~input_a[5];
  assign popcount39_7upc_core_285 = ~(input_a[32] & input_a[14]);
  assign popcount39_7upc_core_290 = input_a[32] & input_a[18];
  assign popcount39_7upc_core_295 = ~(input_a[31] & input_a[25]);
  assign popcount39_7upc_core_296 = input_a[5] ^ input_a[36];
  assign popcount39_7upc_core_300 = input_a[37] | input_a[26];
  assign popcount39_7upc_core_302 = ~(input_a[24] & input_a[10]);
  assign popcount39_7upc_core_303 = ~(input_a[5] & input_a[10]);
  assign popcount39_7upc_core_304_not = ~input_a[13];
  assign popcount39_7upc_core_305 = ~(input_a[30] ^ input_a[3]);

  assign popcount39_7upc_out[0] = input_a[38];
  assign popcount39_7upc_out[1] = input_a[1];
  assign popcount39_7upc_out[2] = 1'b0;
  assign popcount39_7upc_out[3] = 1'b1;
  assign popcount39_7upc_out[4] = input_a[37];
  assign popcount39_7upc_out[5] = 1'b0;
endmodule