// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.84769
// WCE=16.0
// EP=0.92507%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_fggb(input [22:0] input_a, output [4:0] popcount23_fggb_out);
  wire popcount23_fggb_core_026;
  wire popcount23_fggb_core_027;
  wire popcount23_fggb_core_029;
  wire popcount23_fggb_core_031;
  wire popcount23_fggb_core_033;
  wire popcount23_fggb_core_034;
  wire popcount23_fggb_core_036;
  wire popcount23_fggb_core_037;
  wire popcount23_fggb_core_038;
  wire popcount23_fggb_core_040;
  wire popcount23_fggb_core_041;
  wire popcount23_fggb_core_043;
  wire popcount23_fggb_core_044;
  wire popcount23_fggb_core_045;
  wire popcount23_fggb_core_046;
  wire popcount23_fggb_core_048;
  wire popcount23_fggb_core_049;
  wire popcount23_fggb_core_050;
  wire popcount23_fggb_core_052;
  wire popcount23_fggb_core_053;
  wire popcount23_fggb_core_055;
  wire popcount23_fggb_core_059;
  wire popcount23_fggb_core_061;
  wire popcount23_fggb_core_063;
  wire popcount23_fggb_core_065;
  wire popcount23_fggb_core_067;
  wire popcount23_fggb_core_068;
  wire popcount23_fggb_core_069;
  wire popcount23_fggb_core_071;
  wire popcount23_fggb_core_078;
  wire popcount23_fggb_core_079;
  wire popcount23_fggb_core_080;
  wire popcount23_fggb_core_081;
  wire popcount23_fggb_core_082;
  wire popcount23_fggb_core_084;
  wire popcount23_fggb_core_085;
  wire popcount23_fggb_core_086;
  wire popcount23_fggb_core_087;
  wire popcount23_fggb_core_088;
  wire popcount23_fggb_core_089;
  wire popcount23_fggb_core_090;
  wire popcount23_fggb_core_093;
  wire popcount23_fggb_core_094;
  wire popcount23_fggb_core_095_not;
  wire popcount23_fggb_core_096;
  wire popcount23_fggb_core_097;
  wire popcount23_fggb_core_099;
  wire popcount23_fggb_core_100_not;
  wire popcount23_fggb_core_101;
  wire popcount23_fggb_core_103;
  wire popcount23_fggb_core_106;
  wire popcount23_fggb_core_107;
  wire popcount23_fggb_core_109;
  wire popcount23_fggb_core_110;
  wire popcount23_fggb_core_111;
  wire popcount23_fggb_core_112_not;
  wire popcount23_fggb_core_115;
  wire popcount23_fggb_core_116;
  wire popcount23_fggb_core_118;
  wire popcount23_fggb_core_119;
  wire popcount23_fggb_core_121;
  wire popcount23_fggb_core_122;
  wire popcount23_fggb_core_124;
  wire popcount23_fggb_core_126;
  wire popcount23_fggb_core_127;
  wire popcount23_fggb_core_128;
  wire popcount23_fggb_core_132;
  wire popcount23_fggb_core_133;
  wire popcount23_fggb_core_134;
  wire popcount23_fggb_core_135;
  wire popcount23_fggb_core_136;
  wire popcount23_fggb_core_137;
  wire popcount23_fggb_core_138;
  wire popcount23_fggb_core_139;
  wire popcount23_fggb_core_140;
  wire popcount23_fggb_core_141;
  wire popcount23_fggb_core_142;
  wire popcount23_fggb_core_145;
  wire popcount23_fggb_core_146;
  wire popcount23_fggb_core_147;
  wire popcount23_fggb_core_148;
  wire popcount23_fggb_core_149;
  wire popcount23_fggb_core_154;
  wire popcount23_fggb_core_156;
  wire popcount23_fggb_core_157;
  wire popcount23_fggb_core_158;
  wire popcount23_fggb_core_160;
  wire popcount23_fggb_core_161;
  wire popcount23_fggb_core_163;
  wire popcount23_fggb_core_164;
  wire popcount23_fggb_core_165;
  wire popcount23_fggb_core_168;
  wire popcount23_fggb_core_169;

  assign popcount23_fggb_core_026 = input_a[19] | input_a[8];
  assign popcount23_fggb_core_027 = input_a[13] | input_a[15];
  assign popcount23_fggb_core_029 = ~input_a[5];
  assign popcount23_fggb_core_031 = input_a[15] & input_a[8];
  assign popcount23_fggb_core_033 = ~(input_a[20] & input_a[2]);
  assign popcount23_fggb_core_034 = input_a[6] & input_a[15];
  assign popcount23_fggb_core_036 = ~(input_a[0] & input_a[4]);
  assign popcount23_fggb_core_037 = input_a[21] | input_a[14];
  assign popcount23_fggb_core_038 = ~(input_a[10] & input_a[22]);
  assign popcount23_fggb_core_040 = input_a[20] | input_a[0];
  assign popcount23_fggb_core_041 = ~(input_a[14] | input_a[1]);
  assign popcount23_fggb_core_043 = ~(input_a[4] & input_a[17]);
  assign popcount23_fggb_core_044 = ~(input_a[19] ^ input_a[22]);
  assign popcount23_fggb_core_045 = ~(input_a[1] ^ input_a[7]);
  assign popcount23_fggb_core_046 = ~(input_a[1] ^ input_a[0]);
  assign popcount23_fggb_core_048 = input_a[6] & input_a[5];
  assign popcount23_fggb_core_049 = ~(input_a[10] ^ input_a[17]);
  assign popcount23_fggb_core_050 = ~(input_a[17] | input_a[22]);
  assign popcount23_fggb_core_052 = input_a[4] ^ input_a[7];
  assign popcount23_fggb_core_053 = ~(input_a[11] | input_a[21]);
  assign popcount23_fggb_core_055 = input_a[14] | input_a[3];
  assign popcount23_fggb_core_059 = ~input_a[2];
  assign popcount23_fggb_core_061 = input_a[1] | input_a[16];
  assign popcount23_fggb_core_063 = input_a[3] ^ input_a[15];
  assign popcount23_fggb_core_065 = input_a[13] | input_a[21];
  assign popcount23_fggb_core_067 = input_a[3] & input_a[13];
  assign popcount23_fggb_core_068 = ~(input_a[14] & input_a[13]);
  assign popcount23_fggb_core_069 = input_a[2] & input_a[9];
  assign popcount23_fggb_core_071 = ~input_a[21];
  assign popcount23_fggb_core_078 = input_a[11] ^ input_a[8];
  assign popcount23_fggb_core_079 = ~input_a[19];
  assign popcount23_fggb_core_080 = ~input_a[2];
  assign popcount23_fggb_core_081 = input_a[13] | input_a[6];
  assign popcount23_fggb_core_082 = ~(input_a[13] & input_a[18]);
  assign popcount23_fggb_core_084 = input_a[18] ^ input_a[9];
  assign popcount23_fggb_core_085 = ~(input_a[10] | input_a[10]);
  assign popcount23_fggb_core_086 = input_a[5] | input_a[13];
  assign popcount23_fggb_core_087 = ~(input_a[21] | input_a[8]);
  assign popcount23_fggb_core_088 = input_a[4] & input_a[21];
  assign popcount23_fggb_core_089 = ~(input_a[9] ^ input_a[4]);
  assign popcount23_fggb_core_090 = ~(input_a[7] ^ input_a[1]);
  assign popcount23_fggb_core_093 = ~(input_a[9] | input_a[11]);
  assign popcount23_fggb_core_094 = ~(input_a[22] | input_a[4]);
  assign popcount23_fggb_core_095_not = ~input_a[11];
  assign popcount23_fggb_core_096 = ~(input_a[10] ^ input_a[0]);
  assign popcount23_fggb_core_097 = input_a[8] | input_a[11];
  assign popcount23_fggb_core_099 = input_a[22] ^ input_a[11];
  assign popcount23_fggb_core_100_not = ~input_a[10];
  assign popcount23_fggb_core_101 = ~(input_a[5] & input_a[13]);
  assign popcount23_fggb_core_103 = ~(input_a[12] ^ input_a[20]);
  assign popcount23_fggb_core_106 = ~(input_a[7] & input_a[2]);
  assign popcount23_fggb_core_107 = input_a[2] | input_a[2];
  assign popcount23_fggb_core_109 = ~(input_a[6] & input_a[22]);
  assign popcount23_fggb_core_110 = ~(input_a[0] | input_a[15]);
  assign popcount23_fggb_core_111 = ~(input_a[19] ^ input_a[21]);
  assign popcount23_fggb_core_112_not = ~input_a[22];
  assign popcount23_fggb_core_115 = ~(input_a[3] ^ input_a[16]);
  assign popcount23_fggb_core_116 = input_a[8] | input_a[20];
  assign popcount23_fggb_core_118 = input_a[22] & input_a[2];
  assign popcount23_fggb_core_119 = ~(input_a[4] | input_a[6]);
  assign popcount23_fggb_core_121 = input_a[16] | input_a[18];
  assign popcount23_fggb_core_122 = input_a[9] | input_a[19];
  assign popcount23_fggb_core_124 = ~(input_a[8] | input_a[0]);
  assign popcount23_fggb_core_126 = input_a[6] & input_a[4];
  assign popcount23_fggb_core_127 = ~(input_a[9] ^ input_a[14]);
  assign popcount23_fggb_core_128 = input_a[19] & input_a[1];
  assign popcount23_fggb_core_132 = ~(input_a[14] & input_a[17]);
  assign popcount23_fggb_core_133 = input_a[8] & input_a[2];
  assign popcount23_fggb_core_134 = ~(input_a[20] | input_a[9]);
  assign popcount23_fggb_core_135 = input_a[8] & input_a[4];
  assign popcount23_fggb_core_136 = input_a[21] & input_a[12];
  assign popcount23_fggb_core_137 = input_a[14] ^ input_a[3];
  assign popcount23_fggb_core_138 = input_a[13] ^ input_a[14];
  assign popcount23_fggb_core_139 = ~input_a[3];
  assign popcount23_fggb_core_140 = input_a[4] | input_a[6];
  assign popcount23_fggb_core_141 = input_a[0] | input_a[18];
  assign popcount23_fggb_core_142 = input_a[4] & input_a[18];
  assign popcount23_fggb_core_145 = ~(input_a[11] & input_a[7]);
  assign popcount23_fggb_core_146 = ~(input_a[15] | input_a[2]);
  assign popcount23_fggb_core_147 = ~(input_a[1] | input_a[17]);
  assign popcount23_fggb_core_148 = ~(input_a[6] & input_a[8]);
  assign popcount23_fggb_core_149 = input_a[13] & input_a[18];
  assign popcount23_fggb_core_154 = input_a[14] & input_a[7];
  assign popcount23_fggb_core_156 = ~(input_a[17] & input_a[9]);
  assign popcount23_fggb_core_157 = input_a[5] & input_a[16];
  assign popcount23_fggb_core_158 = input_a[14] ^ input_a[0];
  assign popcount23_fggb_core_160 = input_a[6] | input_a[12];
  assign popcount23_fggb_core_161 = input_a[19] | input_a[15];
  assign popcount23_fggb_core_163 = ~(input_a[21] | input_a[13]);
  assign popcount23_fggb_core_164 = ~(input_a[14] & input_a[17]);
  assign popcount23_fggb_core_165 = ~(input_a[10] ^ input_a[19]);
  assign popcount23_fggb_core_168 = ~(input_a[12] & input_a[15]);
  assign popcount23_fggb_core_169 = ~input_a[4];

  assign popcount23_fggb_out[0] = input_a[7];
  assign popcount23_fggb_out[1] = input_a[9];
  assign popcount23_fggb_out[2] = 1'b1;
  assign popcount23_fggb_out[3] = input_a[10];
  assign popcount23_fggb_out[4] = 1'b0;
endmodule