// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.70158
// WCE=19.0
// EP=0.884422%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_sqxy(input [33:0] input_a, output [5:0] popcount34_sqxy_out);
  wire popcount34_sqxy_core_038;
  wire popcount34_sqxy_core_039;
  wire popcount34_sqxy_core_040;
  wire popcount34_sqxy_core_041;
  wire popcount34_sqxy_core_042_not;
  wire popcount34_sqxy_core_043;
  wire popcount34_sqxy_core_047;
  wire popcount34_sqxy_core_049;
  wire popcount34_sqxy_core_050;
  wire popcount34_sqxy_core_052;
  wire popcount34_sqxy_core_055;
  wire popcount34_sqxy_core_056;
  wire popcount34_sqxy_core_057;
  wire popcount34_sqxy_core_060;
  wire popcount34_sqxy_core_062;
  wire popcount34_sqxy_core_063;
  wire popcount34_sqxy_core_065;
  wire popcount34_sqxy_core_067;
  wire popcount34_sqxy_core_068;
  wire popcount34_sqxy_core_070;
  wire popcount34_sqxy_core_073;
  wire popcount34_sqxy_core_074;
  wire popcount34_sqxy_core_075;
  wire popcount34_sqxy_core_076;
  wire popcount34_sqxy_core_077;
  wire popcount34_sqxy_core_082;
  wire popcount34_sqxy_core_083;
  wire popcount34_sqxy_core_084;
  wire popcount34_sqxy_core_085;
  wire popcount34_sqxy_core_086;
  wire popcount34_sqxy_core_087;
  wire popcount34_sqxy_core_088;
  wire popcount34_sqxy_core_089;
  wire popcount34_sqxy_core_090_not;
  wire popcount34_sqxy_core_091;
  wire popcount34_sqxy_core_094;
  wire popcount34_sqxy_core_096;
  wire popcount34_sqxy_core_099;
  wire popcount34_sqxy_core_101;
  wire popcount34_sqxy_core_102;
  wire popcount34_sqxy_core_105;
  wire popcount34_sqxy_core_107;
  wire popcount34_sqxy_core_108;
  wire popcount34_sqxy_core_110;
  wire popcount34_sqxy_core_111;
  wire popcount34_sqxy_core_112;
  wire popcount34_sqxy_core_113;
  wire popcount34_sqxy_core_114;
  wire popcount34_sqxy_core_115;
  wire popcount34_sqxy_core_117;
  wire popcount34_sqxy_core_120;
  wire popcount34_sqxy_core_121;
  wire popcount34_sqxy_core_123;
  wire popcount34_sqxy_core_124;
  wire popcount34_sqxy_core_125;
  wire popcount34_sqxy_core_126;
  wire popcount34_sqxy_core_128;
  wire popcount34_sqxy_core_130;
  wire popcount34_sqxy_core_131;
  wire popcount34_sqxy_core_132;
  wire popcount34_sqxy_core_133;
  wire popcount34_sqxy_core_134;
  wire popcount34_sqxy_core_135;
  wire popcount34_sqxy_core_136;
  wire popcount34_sqxy_core_137;
  wire popcount34_sqxy_core_139;
  wire popcount34_sqxy_core_141;
  wire popcount34_sqxy_core_142;
  wire popcount34_sqxy_core_143;
  wire popcount34_sqxy_core_144;
  wire popcount34_sqxy_core_146;
  wire popcount34_sqxy_core_147;
  wire popcount34_sqxy_core_149_not;
  wire popcount34_sqxy_core_150;
  wire popcount34_sqxy_core_151;
  wire popcount34_sqxy_core_153_not;
  wire popcount34_sqxy_core_154;
  wire popcount34_sqxy_core_155;
  wire popcount34_sqxy_core_156;
  wire popcount34_sqxy_core_159;
  wire popcount34_sqxy_core_161;
  wire popcount34_sqxy_core_163;
  wire popcount34_sqxy_core_166;
  wire popcount34_sqxy_core_167;
  wire popcount34_sqxy_core_168;
  wire popcount34_sqxy_core_170;
  wire popcount34_sqxy_core_171;
  wire popcount34_sqxy_core_172;
  wire popcount34_sqxy_core_174;
  wire popcount34_sqxy_core_176;
  wire popcount34_sqxy_core_177;
  wire popcount34_sqxy_core_179;
  wire popcount34_sqxy_core_183;
  wire popcount34_sqxy_core_184;
  wire popcount34_sqxy_core_186;
  wire popcount34_sqxy_core_187;
  wire popcount34_sqxy_core_189;
  wire popcount34_sqxy_core_190;
  wire popcount34_sqxy_core_193;
  wire popcount34_sqxy_core_194;
  wire popcount34_sqxy_core_195;
  wire popcount34_sqxy_core_196;
  wire popcount34_sqxy_core_197;
  wire popcount34_sqxy_core_200;
  wire popcount34_sqxy_core_201;
  wire popcount34_sqxy_core_202;
  wire popcount34_sqxy_core_203;
  wire popcount34_sqxy_core_204;
  wire popcount34_sqxy_core_205;
  wire popcount34_sqxy_core_206;
  wire popcount34_sqxy_core_207;
  wire popcount34_sqxy_core_209_not;
  wire popcount34_sqxy_core_210;
  wire popcount34_sqxy_core_212;
  wire popcount34_sqxy_core_213;
  wire popcount34_sqxy_core_214;
  wire popcount34_sqxy_core_218;
  wire popcount34_sqxy_core_219;
  wire popcount34_sqxy_core_220;
  wire popcount34_sqxy_core_221;
  wire popcount34_sqxy_core_222;
  wire popcount34_sqxy_core_227_not;
  wire popcount34_sqxy_core_229;
  wire popcount34_sqxy_core_230;
  wire popcount34_sqxy_core_231;
  wire popcount34_sqxy_core_232;
  wire popcount34_sqxy_core_233;
  wire popcount34_sqxy_core_234;
  wire popcount34_sqxy_core_235;
  wire popcount34_sqxy_core_237;
  wire popcount34_sqxy_core_238;
  wire popcount34_sqxy_core_239;
  wire popcount34_sqxy_core_241_not;
  wire popcount34_sqxy_core_242;
  wire popcount34_sqxy_core_243_not;
  wire popcount34_sqxy_core_249;
  wire popcount34_sqxy_core_250;
  wire popcount34_sqxy_core_251;
  wire popcount34_sqxy_core_252;

  assign popcount34_sqxy_core_038 = ~(input_a[13] & input_a[9]);
  assign popcount34_sqxy_core_039 = ~(input_a[13] | input_a[7]);
  assign popcount34_sqxy_core_040 = ~(input_a[10] & input_a[15]);
  assign popcount34_sqxy_core_041 = input_a[12] & input_a[11];
  assign popcount34_sqxy_core_042_not = ~input_a[18];
  assign popcount34_sqxy_core_043 = ~(input_a[28] | input_a[4]);
  assign popcount34_sqxy_core_047 = ~(input_a[22] | input_a[33]);
  assign popcount34_sqxy_core_049 = input_a[10] | input_a[26];
  assign popcount34_sqxy_core_050 = input_a[17] & input_a[16];
  assign popcount34_sqxy_core_052 = ~(input_a[23] ^ input_a[13]);
  assign popcount34_sqxy_core_055 = input_a[11] ^ input_a[20];
  assign popcount34_sqxy_core_056 = input_a[12] | input_a[12];
  assign popcount34_sqxy_core_057 = ~(input_a[16] & input_a[6]);
  assign popcount34_sqxy_core_060 = ~(input_a[13] ^ input_a[30]);
  assign popcount34_sqxy_core_062 = ~(input_a[2] & input_a[7]);
  assign popcount34_sqxy_core_063 = input_a[2] ^ input_a[14];
  assign popcount34_sqxy_core_065 = ~(input_a[1] ^ input_a[14]);
  assign popcount34_sqxy_core_067 = ~input_a[12];
  assign popcount34_sqxy_core_068 = ~(input_a[27] | input_a[26]);
  assign popcount34_sqxy_core_070 = ~(input_a[29] ^ input_a[19]);
  assign popcount34_sqxy_core_073 = ~(input_a[26] & input_a[26]);
  assign popcount34_sqxy_core_074 = ~input_a[7];
  assign popcount34_sqxy_core_075 = ~(input_a[18] ^ input_a[28]);
  assign popcount34_sqxy_core_076 = input_a[13] | input_a[24];
  assign popcount34_sqxy_core_077 = input_a[20] | input_a[12];
  assign popcount34_sqxy_core_082 = ~(input_a[7] ^ input_a[32]);
  assign popcount34_sqxy_core_083 = input_a[4] & input_a[9];
  assign popcount34_sqxy_core_084 = ~(input_a[14] | input_a[29]);
  assign popcount34_sqxy_core_085 = ~(input_a[31] ^ input_a[18]);
  assign popcount34_sqxy_core_086 = ~(input_a[25] & input_a[1]);
  assign popcount34_sqxy_core_087 = ~(input_a[15] ^ input_a[6]);
  assign popcount34_sqxy_core_088 = ~input_a[12];
  assign popcount34_sqxy_core_089 = input_a[3] ^ input_a[32];
  assign popcount34_sqxy_core_090_not = ~input_a[31];
  assign popcount34_sqxy_core_091 = input_a[7] | input_a[17];
  assign popcount34_sqxy_core_094 = ~input_a[31];
  assign popcount34_sqxy_core_096 = input_a[9] & input_a[6];
  assign popcount34_sqxy_core_099 = input_a[18] ^ input_a[17];
  assign popcount34_sqxy_core_101 = ~(input_a[28] & input_a[13]);
  assign popcount34_sqxy_core_102 = input_a[6] ^ input_a[33];
  assign popcount34_sqxy_core_105 = input_a[29] ^ input_a[32];
  assign popcount34_sqxy_core_107 = input_a[0] ^ input_a[2];
  assign popcount34_sqxy_core_108 = input_a[11] & input_a[12];
  assign popcount34_sqxy_core_110 = ~(input_a[32] ^ input_a[10]);
  assign popcount34_sqxy_core_111 = ~(input_a[30] & input_a[33]);
  assign popcount34_sqxy_core_112 = input_a[29] ^ input_a[31];
  assign popcount34_sqxy_core_113 = input_a[16] | input_a[5];
  assign popcount34_sqxy_core_114 = input_a[10] | input_a[13];
  assign popcount34_sqxy_core_115 = input_a[31] | input_a[5];
  assign popcount34_sqxy_core_117 = input_a[4] ^ input_a[13];
  assign popcount34_sqxy_core_120 = input_a[9] | input_a[29];
  assign popcount34_sqxy_core_121 = ~input_a[13];
  assign popcount34_sqxy_core_123 = input_a[0] ^ input_a[28];
  assign popcount34_sqxy_core_124 = ~(input_a[17] ^ input_a[25]);
  assign popcount34_sqxy_core_125 = input_a[30] | input_a[11];
  assign popcount34_sqxy_core_126 = ~(input_a[29] | input_a[3]);
  assign popcount34_sqxy_core_128 = ~(input_a[13] ^ input_a[13]);
  assign popcount34_sqxy_core_130 = input_a[1] & input_a[10];
  assign popcount34_sqxy_core_131 = input_a[5] ^ input_a[10];
  assign popcount34_sqxy_core_132 = input_a[6] | input_a[27];
  assign popcount34_sqxy_core_133 = ~(input_a[32] & input_a[32]);
  assign popcount34_sqxy_core_134 = ~(input_a[25] | input_a[28]);
  assign popcount34_sqxy_core_135 = ~(input_a[33] | input_a[17]);
  assign popcount34_sqxy_core_136 = ~(input_a[33] | input_a[17]);
  assign popcount34_sqxy_core_137 = input_a[17] ^ input_a[10];
  assign popcount34_sqxy_core_139 = ~(input_a[27] | input_a[23]);
  assign popcount34_sqxy_core_141 = ~(input_a[19] & input_a[1]);
  assign popcount34_sqxy_core_142 = ~input_a[20];
  assign popcount34_sqxy_core_143 = input_a[11] & input_a[13];
  assign popcount34_sqxy_core_144 = input_a[10] | input_a[18];
  assign popcount34_sqxy_core_146 = input_a[25] & input_a[28];
  assign popcount34_sqxy_core_147 = ~(input_a[6] ^ input_a[12]);
  assign popcount34_sqxy_core_149_not = ~input_a[19];
  assign popcount34_sqxy_core_150 = input_a[27] | input_a[2];
  assign popcount34_sqxy_core_151 = ~(input_a[3] ^ input_a[24]);
  assign popcount34_sqxy_core_153_not = ~input_a[27];
  assign popcount34_sqxy_core_154 = input_a[16] & input_a[26];
  assign popcount34_sqxy_core_155 = ~(input_a[30] | input_a[14]);
  assign popcount34_sqxy_core_156 = input_a[0] ^ input_a[16];
  assign popcount34_sqxy_core_159 = input_a[1] ^ input_a[1];
  assign popcount34_sqxy_core_161 = ~(input_a[13] & input_a[10]);
  assign popcount34_sqxy_core_163 = input_a[9] | input_a[12];
  assign popcount34_sqxy_core_166 = input_a[18] & input_a[6];
  assign popcount34_sqxy_core_167 = ~(input_a[32] & input_a[9]);
  assign popcount34_sqxy_core_168 = ~(input_a[29] | input_a[31]);
  assign popcount34_sqxy_core_170 = ~(input_a[10] & input_a[21]);
  assign popcount34_sqxy_core_171 = ~(input_a[0] | input_a[28]);
  assign popcount34_sqxy_core_172 = ~(input_a[18] & input_a[2]);
  assign popcount34_sqxy_core_174 = ~input_a[25];
  assign popcount34_sqxy_core_176 = ~input_a[27];
  assign popcount34_sqxy_core_177 = input_a[28] | input_a[2];
  assign popcount34_sqxy_core_179 = ~(input_a[30] | input_a[23]);
  assign popcount34_sqxy_core_183 = ~input_a[5];
  assign popcount34_sqxy_core_184 = ~input_a[10];
  assign popcount34_sqxy_core_186 = ~(input_a[25] | input_a[17]);
  assign popcount34_sqxy_core_187 = input_a[28] ^ input_a[14];
  assign popcount34_sqxy_core_189 = ~input_a[6];
  assign popcount34_sqxy_core_190 = input_a[13] | input_a[31];
  assign popcount34_sqxy_core_193 = input_a[9] & input_a[11];
  assign popcount34_sqxy_core_194 = input_a[3] | input_a[13];
  assign popcount34_sqxy_core_195 = input_a[19] ^ input_a[17];
  assign popcount34_sqxy_core_196 = input_a[14] | input_a[5];
  assign popcount34_sqxy_core_197 = ~(input_a[32] & input_a[6]);
  assign popcount34_sqxy_core_200 = input_a[11] ^ input_a[21];
  assign popcount34_sqxy_core_201 = input_a[28] ^ input_a[16];
  assign popcount34_sqxy_core_202 = ~(input_a[2] & input_a[2]);
  assign popcount34_sqxy_core_203 = ~(input_a[26] & input_a[33]);
  assign popcount34_sqxy_core_204 = ~input_a[8];
  assign popcount34_sqxy_core_205 = ~(input_a[26] & input_a[0]);
  assign popcount34_sqxy_core_206 = ~input_a[6];
  assign popcount34_sqxy_core_207 = input_a[4] | input_a[7];
  assign popcount34_sqxy_core_209_not = ~input_a[2];
  assign popcount34_sqxy_core_210 = input_a[18] ^ input_a[15];
  assign popcount34_sqxy_core_212 = ~(input_a[11] ^ input_a[5]);
  assign popcount34_sqxy_core_213 = input_a[19] | input_a[18];
  assign popcount34_sqxy_core_214 = input_a[3] & input_a[23];
  assign popcount34_sqxy_core_218 = ~(input_a[32] | input_a[6]);
  assign popcount34_sqxy_core_219 = ~(input_a[4] & input_a[1]);
  assign popcount34_sqxy_core_220 = ~(input_a[15] ^ input_a[19]);
  assign popcount34_sqxy_core_221 = ~(input_a[32] & input_a[18]);
  assign popcount34_sqxy_core_222 = ~(input_a[7] & input_a[2]);
  assign popcount34_sqxy_core_227_not = ~input_a[19];
  assign popcount34_sqxy_core_229 = input_a[29] | input_a[17];
  assign popcount34_sqxy_core_230 = ~input_a[22];
  assign popcount34_sqxy_core_231 = input_a[14] ^ input_a[18];
  assign popcount34_sqxy_core_232 = input_a[26] & input_a[26];
  assign popcount34_sqxy_core_233 = ~(input_a[2] ^ input_a[21]);
  assign popcount34_sqxy_core_234 = ~(input_a[14] & input_a[26]);
  assign popcount34_sqxy_core_235 = ~input_a[15];
  assign popcount34_sqxy_core_237 = ~(input_a[21] | input_a[33]);
  assign popcount34_sqxy_core_238 = ~(input_a[30] & input_a[33]);
  assign popcount34_sqxy_core_239 = input_a[23] ^ input_a[32];
  assign popcount34_sqxy_core_241_not = ~input_a[1];
  assign popcount34_sqxy_core_242 = ~input_a[1];
  assign popcount34_sqxy_core_243_not = ~input_a[1];
  assign popcount34_sqxy_core_249 = ~(input_a[0] ^ input_a[17]);
  assign popcount34_sqxy_core_250 = ~(input_a[4] | input_a[13]);
  assign popcount34_sqxy_core_251 = ~(input_a[2] | input_a[1]);
  assign popcount34_sqxy_core_252 = ~(input_a[12] & input_a[26]);

  assign popcount34_sqxy_out[0] = 1'b0;
  assign popcount34_sqxy_out[1] = 1'b0;
  assign popcount34_sqxy_out[2] = input_a[6];
  assign popcount34_sqxy_out[3] = 1'b0;
  assign popcount34_sqxy_out[4] = 1'b1;
  assign popcount34_sqxy_out[5] = 1'b0;
endmodule