// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.85013
// WCE=22.0
// EP=0.945404%
// Printed PDK parameters:
//  Area=33604206.0
//  Delay=62162432.0
//  Power=1195300.0

module popcount43_zk3b(input [42:0] input_a, output [5:0] popcount43_zk3b_out);
  wire popcount43_zk3b_core_045;
  wire popcount43_zk3b_core_046;
  wire popcount43_zk3b_core_047;
  wire popcount43_zk3b_core_048;
  wire popcount43_zk3b_core_049;
  wire popcount43_zk3b_core_056;
  wire popcount43_zk3b_core_058;
  wire popcount43_zk3b_core_062;
  wire popcount43_zk3b_core_063;
  wire popcount43_zk3b_core_065;
  wire popcount43_zk3b_core_066;
  wire popcount43_zk3b_core_067;
  wire popcount43_zk3b_core_068;
  wire popcount43_zk3b_core_072;
  wire popcount43_zk3b_core_073;
  wire popcount43_zk3b_core_077;
  wire popcount43_zk3b_core_078;
  wire popcount43_zk3b_core_080;
  wire popcount43_zk3b_core_082_not;
  wire popcount43_zk3b_core_086;
  wire popcount43_zk3b_core_087;
  wire popcount43_zk3b_core_089;
  wire popcount43_zk3b_core_091;
  wire popcount43_zk3b_core_093;
  wire popcount43_zk3b_core_094;
  wire popcount43_zk3b_core_095;
  wire popcount43_zk3b_core_097;
  wire popcount43_zk3b_core_098;
  wire popcount43_zk3b_core_099;
  wire popcount43_zk3b_core_100;
  wire popcount43_zk3b_core_106;
  wire popcount43_zk3b_core_107;
  wire popcount43_zk3b_core_113;
  wire popcount43_zk3b_core_114;
  wire popcount43_zk3b_core_115;
  wire popcount43_zk3b_core_116;
  wire popcount43_zk3b_core_117;
  wire popcount43_zk3b_core_118;
  wire popcount43_zk3b_core_119;
  wire popcount43_zk3b_core_120;
  wire popcount43_zk3b_core_121;
  wire popcount43_zk3b_core_122;
  wire popcount43_zk3b_core_123;
  wire popcount43_zk3b_core_124;
  wire popcount43_zk3b_core_125;
  wire popcount43_zk3b_core_126;
  wire popcount43_zk3b_core_127;
  wire popcount43_zk3b_core_128;
  wire popcount43_zk3b_core_129;
  wire popcount43_zk3b_core_130;
  wire popcount43_zk3b_core_131;
  wire popcount43_zk3b_core_133;
  wire popcount43_zk3b_core_135;
  wire popcount43_zk3b_core_142;
  wire popcount43_zk3b_core_144;
  wire popcount43_zk3b_core_145;
  wire popcount43_zk3b_core_152;
  wire popcount43_zk3b_core_153;
  wire popcount43_zk3b_core_154;
  wire popcount43_zk3b_core_155;
  wire popcount43_zk3b_core_157;
  wire popcount43_zk3b_core_158;
  wire popcount43_zk3b_core_159;
  wire popcount43_zk3b_core_160;
  wire popcount43_zk3b_core_161;
  wire popcount43_zk3b_core_162;
  wire popcount43_zk3b_core_163;
  wire popcount43_zk3b_core_164;
  wire popcount43_zk3b_core_165;
  wire popcount43_zk3b_core_166;
  wire popcount43_zk3b_core_167;
  wire popcount43_zk3b_core_168;
  wire popcount43_zk3b_core_169;
  wire popcount43_zk3b_core_170;
  wire popcount43_zk3b_core_172;
  wire popcount43_zk3b_core_175;
  wire popcount43_zk3b_core_179;
  wire popcount43_zk3b_core_183;
  wire popcount43_zk3b_core_185;
  wire popcount43_zk3b_core_186;
  wire popcount43_zk3b_core_187;
  wire popcount43_zk3b_core_188;
  wire popcount43_zk3b_core_190;
  wire popcount43_zk3b_core_193;
  wire popcount43_zk3b_core_194;
  wire popcount43_zk3b_core_195;
  wire popcount43_zk3b_core_196;
  wire popcount43_zk3b_core_197;
  wire popcount43_zk3b_core_198;
  wire popcount43_zk3b_core_199;
  wire popcount43_zk3b_core_201;
  wire popcount43_zk3b_core_202;
  wire popcount43_zk3b_core_204;
  wire popcount43_zk3b_core_205;
  wire popcount43_zk3b_core_206;
  wire popcount43_zk3b_core_207;
  wire popcount43_zk3b_core_208;
  wire popcount43_zk3b_core_209;
  wire popcount43_zk3b_core_210;
  wire popcount43_zk3b_core_211;
  wire popcount43_zk3b_core_212;
  wire popcount43_zk3b_core_213;
  wire popcount43_zk3b_core_214;
  wire popcount43_zk3b_core_215;
  wire popcount43_zk3b_core_217;
  wire popcount43_zk3b_core_218;
  wire popcount43_zk3b_core_220;
  wire popcount43_zk3b_core_221;
  wire popcount43_zk3b_core_226;
  wire popcount43_zk3b_core_227;
  wire popcount43_zk3b_core_228;
  wire popcount43_zk3b_core_234;
  wire popcount43_zk3b_core_235;
  wire popcount43_zk3b_core_236;
  wire popcount43_zk3b_core_240;
  wire popcount43_zk3b_core_242;
  wire popcount43_zk3b_core_244;
  wire popcount43_zk3b_core_245;
  wire popcount43_zk3b_core_246;
  wire popcount43_zk3b_core_247;
  wire popcount43_zk3b_core_248;
  wire popcount43_zk3b_core_250;
  wire popcount43_zk3b_core_251;
  wire popcount43_zk3b_core_256;
  wire popcount43_zk3b_core_257;
  wire popcount43_zk3b_core_258;
  wire popcount43_zk3b_core_260;
  wire popcount43_zk3b_core_265;
  wire popcount43_zk3b_core_266;
  wire popcount43_zk3b_core_267;
  wire popcount43_zk3b_core_269;
  wire popcount43_zk3b_core_270;
  wire popcount43_zk3b_core_271_not;
  wire popcount43_zk3b_core_272;
  wire popcount43_zk3b_core_274;
  wire popcount43_zk3b_core_275;
  wire popcount43_zk3b_core_277;
  wire popcount43_zk3b_core_278;
  wire popcount43_zk3b_core_279;
  wire popcount43_zk3b_core_280;
  wire popcount43_zk3b_core_283;
  wire popcount43_zk3b_core_284;
  wire popcount43_zk3b_core_285;
  wire popcount43_zk3b_core_286;
  wire popcount43_zk3b_core_288;
  wire popcount43_zk3b_core_290;
  wire popcount43_zk3b_core_293;
  wire popcount43_zk3b_core_294;
  wire popcount43_zk3b_core_296;
  wire popcount43_zk3b_core_297;
  wire popcount43_zk3b_core_298;
  wire popcount43_zk3b_core_299;
  wire popcount43_zk3b_core_301;
  wire popcount43_zk3b_core_306;
  wire popcount43_zk3b_core_317;
  wire popcount43_zk3b_core_319;
  wire popcount43_zk3b_core_322;
  wire popcount43_zk3b_core_323;
  wire popcount43_zk3b_core_324;
  wire popcount43_zk3b_core_325;
  wire popcount43_zk3b_core_326;
  wire popcount43_zk3b_core_327;
  wire popcount43_zk3b_core_328;
  wire popcount43_zk3b_core_329;
  wire popcount43_zk3b_core_330;
  wire popcount43_zk3b_core_331;
  wire popcount43_zk3b_core_332;
  wire popcount43_zk3b_core_333;
  wire popcount43_zk3b_core_334;
  wire popcount43_zk3b_core_335;
  wire popcount43_zk3b_core_337;
  wire popcount43_zk3b_core_339;
  wire popcount43_zk3b_core_340;

  assign popcount43_zk3b_core_045 = ~(input_a[0] | input_a[3]);
  assign popcount43_zk3b_core_046 = input_a[0] & input_a[41];
  assign popcount43_zk3b_core_047 = input_a[42] & input_a[37];
  assign popcount43_zk3b_core_048 = input_a[3] & input_a[4];
  assign popcount43_zk3b_core_049 = input_a[2] | input_a[8];
  assign popcount43_zk3b_core_056 = popcount43_zk3b_core_046 & popcount43_zk3b_core_048;
  assign popcount43_zk3b_core_058 = input_a[34] & input_a[27];
  assign popcount43_zk3b_core_062 = ~(input_a[34] & input_a[6]);
  assign popcount43_zk3b_core_063 = input_a[23] & input_a[11];
  assign popcount43_zk3b_core_065 = input_a[2] & input_a[38];
  assign popcount43_zk3b_core_066 = input_a[8] & input_a[5];
  assign popcount43_zk3b_core_067 = ~(input_a[29] & input_a[32]);
  assign popcount43_zk3b_core_068 = ~popcount43_zk3b_core_065;
  assign popcount43_zk3b_core_072 = popcount43_zk3b_core_063 ^ popcount43_zk3b_core_068;
  assign popcount43_zk3b_core_073 = popcount43_zk3b_core_063 & popcount43_zk3b_core_068;
  assign popcount43_zk3b_core_077 = popcount43_zk3b_core_065 | popcount43_zk3b_core_073;
  assign popcount43_zk3b_core_078 = popcount43_zk3b_core_065 & popcount43_zk3b_core_073;
  assign popcount43_zk3b_core_080 = ~(input_a[4] & input_a[39]);
  assign popcount43_zk3b_core_082_not = ~input_a[23];
  assign popcount43_zk3b_core_086 = popcount43_zk3b_core_056 ^ popcount43_zk3b_core_077;
  assign popcount43_zk3b_core_087 = popcount43_zk3b_core_056 & popcount43_zk3b_core_077;
  assign popcount43_zk3b_core_089 = ~(input_a[40] ^ input_a[21]);
  assign popcount43_zk3b_core_091 = input_a[6] & popcount43_zk3b_core_078;
  assign popcount43_zk3b_core_093 = popcount43_zk3b_core_091 | popcount43_zk3b_core_087;
  assign popcount43_zk3b_core_094 = input_a[4] ^ input_a[6];
  assign popcount43_zk3b_core_095 = ~(input_a[41] & input_a[26]);
  assign popcount43_zk3b_core_097 = input_a[32] & input_a[5];
  assign popcount43_zk3b_core_098 = ~(input_a[26] ^ input_a[14]);
  assign popcount43_zk3b_core_099 = input_a[13] & input_a[14];
  assign popcount43_zk3b_core_100 = ~input_a[7];
  assign popcount43_zk3b_core_106 = input_a[27] ^ input_a[18];
  assign popcount43_zk3b_core_107 = popcount43_zk3b_core_097 & popcount43_zk3b_core_099;
  assign popcount43_zk3b_core_113 = input_a[16] ^ input_a[17];
  assign popcount43_zk3b_core_114 = input_a[16] & input_a[17];
  assign popcount43_zk3b_core_115 = input_a[15] ^ popcount43_zk3b_core_113;
  assign popcount43_zk3b_core_116 = input_a[15] & popcount43_zk3b_core_113;
  assign popcount43_zk3b_core_117 = popcount43_zk3b_core_114 | popcount43_zk3b_core_116;
  assign popcount43_zk3b_core_118 = ~(input_a[9] | input_a[33]);
  assign popcount43_zk3b_core_119 = input_a[19] | input_a[25];
  assign popcount43_zk3b_core_120 = input_a[19] & input_a[20];
  assign popcount43_zk3b_core_121 = ~(input_a[14] ^ popcount43_zk3b_core_119);
  assign popcount43_zk3b_core_122 = input_a[18] & popcount43_zk3b_core_119;
  assign popcount43_zk3b_core_123 = popcount43_zk3b_core_120 | popcount43_zk3b_core_122;
  assign popcount43_zk3b_core_124 = ~(input_a[28] ^ input_a[9]);
  assign popcount43_zk3b_core_125 = input_a[32] ^ input_a[1];
  assign popcount43_zk3b_core_126 = popcount43_zk3b_core_115 & input_a[27];
  assign popcount43_zk3b_core_127 = popcount43_zk3b_core_117 ^ popcount43_zk3b_core_123;
  assign popcount43_zk3b_core_128 = popcount43_zk3b_core_117 & popcount43_zk3b_core_123;
  assign popcount43_zk3b_core_129 = popcount43_zk3b_core_127 ^ popcount43_zk3b_core_126;
  assign popcount43_zk3b_core_130 = popcount43_zk3b_core_127 & popcount43_zk3b_core_126;
  assign popcount43_zk3b_core_131 = popcount43_zk3b_core_128 | popcount43_zk3b_core_130;
  assign popcount43_zk3b_core_133 = ~input_a[0];
  assign popcount43_zk3b_core_135 = ~(input_a[19] & input_a[35]);
  assign popcount43_zk3b_core_142 = input_a[21] ^ input_a[31];
  assign popcount43_zk3b_core_144 = popcount43_zk3b_core_107 ^ popcount43_zk3b_core_131;
  assign popcount43_zk3b_core_145 = popcount43_zk3b_core_107 & popcount43_zk3b_core_131;
  assign popcount43_zk3b_core_152 = input_a[19] & input_a[16];
  assign popcount43_zk3b_core_153 = input_a[29] ^ input_a[32];
  assign popcount43_zk3b_core_154 = ~(input_a[38] | input_a[10]);
  assign popcount43_zk3b_core_155 = input_a[39] & input_a[26];
  assign popcount43_zk3b_core_157 = popcount43_zk3b_core_072 & popcount43_zk3b_core_129;
  assign popcount43_zk3b_core_158 = input_a[7] ^ input_a[37];
  assign popcount43_zk3b_core_159 = popcount43_zk3b_core_072 & popcount43_zk3b_core_155;
  assign popcount43_zk3b_core_160 = popcount43_zk3b_core_157 | popcount43_zk3b_core_159;
  assign popcount43_zk3b_core_161 = popcount43_zk3b_core_086 ^ popcount43_zk3b_core_144;
  assign popcount43_zk3b_core_162 = popcount43_zk3b_core_086 & popcount43_zk3b_core_144;
  assign popcount43_zk3b_core_163 = popcount43_zk3b_core_161 ^ popcount43_zk3b_core_160;
  assign popcount43_zk3b_core_164 = popcount43_zk3b_core_161 & popcount43_zk3b_core_160;
  assign popcount43_zk3b_core_165 = popcount43_zk3b_core_162 | popcount43_zk3b_core_164;
  assign popcount43_zk3b_core_166 = popcount43_zk3b_core_093 ^ popcount43_zk3b_core_145;
  assign popcount43_zk3b_core_167 = popcount43_zk3b_core_093 & popcount43_zk3b_core_145;
  assign popcount43_zk3b_core_168 = popcount43_zk3b_core_166 ^ popcount43_zk3b_core_165;
  assign popcount43_zk3b_core_169 = popcount43_zk3b_core_166 & popcount43_zk3b_core_165;
  assign popcount43_zk3b_core_170 = popcount43_zk3b_core_167 | popcount43_zk3b_core_169;
  assign popcount43_zk3b_core_172 = input_a[39] | input_a[37];
  assign popcount43_zk3b_core_175 = input_a[9] | input_a[36];
  assign popcount43_zk3b_core_179 = input_a[1] & input_a[12];
  assign popcount43_zk3b_core_183 = ~input_a[14];
  assign popcount43_zk3b_core_185 = ~(input_a[8] | input_a[5]);
  assign popcount43_zk3b_core_186 = ~(input_a[38] ^ input_a[14]);
  assign popcount43_zk3b_core_187 = ~input_a[4];
  assign popcount43_zk3b_core_188 = input_a[0] & input_a[23];
  assign popcount43_zk3b_core_190 = input_a[4] & input_a[15];
  assign popcount43_zk3b_core_193 = ~(input_a[35] ^ input_a[6]);
  assign popcount43_zk3b_core_194 = ~input_a[21];
  assign popcount43_zk3b_core_195 = input_a[1] ^ input_a[9];
  assign popcount43_zk3b_core_196 = ~input_a[35];
  assign popcount43_zk3b_core_197 = input_a[19] & input_a[11];
  assign popcount43_zk3b_core_198 = ~(input_a[5] | input_a[3]);
  assign popcount43_zk3b_core_199 = ~(input_a[41] & input_a[12]);
  assign popcount43_zk3b_core_201 = ~input_a[28];
  assign popcount43_zk3b_core_202 = input_a[10] ^ input_a[13];
  assign popcount43_zk3b_core_204 = ~(input_a[9] ^ input_a[13]);
  assign popcount43_zk3b_core_205 = input_a[15] ^ input_a[24];
  assign popcount43_zk3b_core_206 = ~(input_a[8] & input_a[9]);
  assign popcount43_zk3b_core_207 = ~(input_a[3] ^ input_a[2]);
  assign popcount43_zk3b_core_208 = ~input_a[23];
  assign popcount43_zk3b_core_209 = input_a[15] & input_a[16];
  assign popcount43_zk3b_core_210 = ~input_a[35];
  assign popcount43_zk3b_core_211 = input_a[20] & input_a[40];
  assign popcount43_zk3b_core_212 = ~input_a[31];
  assign popcount43_zk3b_core_213 = ~(input_a[38] & input_a[34]);
  assign popcount43_zk3b_core_214 = ~(input_a[22] | input_a[9]);
  assign popcount43_zk3b_core_215 = input_a[31] & input_a[11];
  assign popcount43_zk3b_core_217 = ~input_a[32];
  assign popcount43_zk3b_core_218 = input_a[6] ^ input_a[40];
  assign popcount43_zk3b_core_220 = ~(input_a[2] ^ input_a[17]);
  assign popcount43_zk3b_core_221 = ~(input_a[14] | input_a[5]);
  assign popcount43_zk3b_core_226 = input_a[17] | input_a[35];
  assign popcount43_zk3b_core_227 = ~(input_a[18] ^ input_a[5]);
  assign popcount43_zk3b_core_228 = input_a[42] & input_a[22];
  assign popcount43_zk3b_core_234 = input_a[30] | input_a[23];
  assign popcount43_zk3b_core_235 = input_a[13] & input_a[37];
  assign popcount43_zk3b_core_236 = input_a[24] & input_a[32];
  assign popcount43_zk3b_core_240 = input_a[4] ^ input_a[42];
  assign popcount43_zk3b_core_242 = ~input_a[13];
  assign popcount43_zk3b_core_244 = ~(input_a[22] | input_a[20]);
  assign popcount43_zk3b_core_245 = input_a[35] & input_a[1];
  assign popcount43_zk3b_core_246 = ~input_a[6];
  assign popcount43_zk3b_core_247 = input_a[24] & input_a[9];
  assign popcount43_zk3b_core_248 = popcount43_zk3b_core_245 | popcount43_zk3b_core_247;
  assign popcount43_zk3b_core_250 = ~(input_a[39] ^ input_a[17]);
  assign popcount43_zk3b_core_251 = ~(input_a[13] ^ input_a[10]);
  assign popcount43_zk3b_core_256 = ~input_a[13];
  assign popcount43_zk3b_core_257 = ~(input_a[31] | input_a[6]);
  assign popcount43_zk3b_core_258 = input_a[38] & input_a[35];
  assign popcount43_zk3b_core_260 = ~(input_a[9] | input_a[2]);
  assign popcount43_zk3b_core_265 = ~(input_a[15] | input_a[15]);
  assign popcount43_zk3b_core_266 = ~(input_a[1] ^ input_a[19]);
  assign popcount43_zk3b_core_267 = ~(input_a[34] & input_a[1]);
  assign popcount43_zk3b_core_269 = ~(input_a[29] | input_a[13]);
  assign popcount43_zk3b_core_270 = ~(input_a[37] ^ input_a[6]);
  assign popcount43_zk3b_core_271_not = ~popcount43_zk3b_core_256;
  assign popcount43_zk3b_core_272 = ~(input_a[36] ^ input_a[18]);
  assign popcount43_zk3b_core_274 = ~(input_a[22] & input_a[9]);
  assign popcount43_zk3b_core_275 = ~(input_a[16] & input_a[19]);
  assign popcount43_zk3b_core_277 = ~(input_a[6] ^ input_a[31]);
  assign popcount43_zk3b_core_278 = ~(input_a[1] ^ input_a[12]);
  assign popcount43_zk3b_core_279 = input_a[32] & input_a[33];
  assign popcount43_zk3b_core_280 = ~(input_a[42] | input_a[11]);
  assign popcount43_zk3b_core_283 = popcount43_zk3b_core_248 & input_a[31];
  assign popcount43_zk3b_core_284 = input_a[0] | input_a[16];
  assign popcount43_zk3b_core_285 = popcount43_zk3b_core_248 & input_a[22];
  assign popcount43_zk3b_core_286 = popcount43_zk3b_core_283 | popcount43_zk3b_core_285;
  assign popcount43_zk3b_core_288 = input_a[36] & input_a[13];
  assign popcount43_zk3b_core_290 = ~(input_a[8] & input_a[10]);
  assign popcount43_zk3b_core_293 = ~(input_a[2] & input_a[34]);
  assign popcount43_zk3b_core_294 = ~(input_a[3] & input_a[37]);
  assign popcount43_zk3b_core_296 = input_a[41] | input_a[20];
  assign popcount43_zk3b_core_297 = ~(input_a[42] | input_a[27]);
  assign popcount43_zk3b_core_298 = input_a[42] | input_a[12];
  assign popcount43_zk3b_core_299 = input_a[17] & input_a[8];
  assign popcount43_zk3b_core_301 = input_a[1] & input_a[36];
  assign popcount43_zk3b_core_306 = ~popcount43_zk3b_core_286;
  assign popcount43_zk3b_core_317 = input_a[5] & input_a[37];
  assign popcount43_zk3b_core_319 = input_a[13] & input_a[36];
  assign popcount43_zk3b_core_322 = popcount43_zk3b_core_163 & input_a[21];
  assign popcount43_zk3b_core_323 = input_a[7] ^ input_a[30];
  assign popcount43_zk3b_core_324 = input_a[7] & input_a[30];
  assign popcount43_zk3b_core_325 = popcount43_zk3b_core_322 | popcount43_zk3b_core_324;
  assign popcount43_zk3b_core_326 = popcount43_zk3b_core_168 | popcount43_zk3b_core_306;
  assign popcount43_zk3b_core_327 = popcount43_zk3b_core_168 & popcount43_zk3b_core_306;
  assign popcount43_zk3b_core_328 = popcount43_zk3b_core_326 ^ popcount43_zk3b_core_325;
  assign popcount43_zk3b_core_329 = popcount43_zk3b_core_326 & popcount43_zk3b_core_325;
  assign popcount43_zk3b_core_330 = popcount43_zk3b_core_327 | popcount43_zk3b_core_329;
  assign popcount43_zk3b_core_331 = popcount43_zk3b_core_170 ^ popcount43_zk3b_core_286;
  assign popcount43_zk3b_core_332 = popcount43_zk3b_core_170 & popcount43_zk3b_core_286;
  assign popcount43_zk3b_core_333 = popcount43_zk3b_core_331 ^ popcount43_zk3b_core_330;
  assign popcount43_zk3b_core_334 = popcount43_zk3b_core_331 & popcount43_zk3b_core_330;
  assign popcount43_zk3b_core_335 = popcount43_zk3b_core_332 | popcount43_zk3b_core_334;
  assign popcount43_zk3b_core_337 = input_a[1] | input_a[11];
  assign popcount43_zk3b_core_339 = ~(input_a[23] | input_a[21]);
  assign popcount43_zk3b_core_340 = input_a[2] & input_a[13];

  assign popcount43_zk3b_out[0] = input_a[37];
  assign popcount43_zk3b_out[1] = input_a[42];
  assign popcount43_zk3b_out[2] = popcount43_zk3b_core_323;
  assign popcount43_zk3b_out[3] = popcount43_zk3b_core_328;
  assign popcount43_zk3b_out[4] = popcount43_zk3b_core_333;
  assign popcount43_zk3b_out[5] = popcount43_zk3b_core_335;
endmodule