// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.75792
// WCE=20.0
// EP=0.921718%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_s0xx(input [26:0] input_a, output [4:0] popcount27_s0xx_out);
  wire popcount27_s0xx_core_032;
  wire popcount27_s0xx_core_033;
  wire popcount27_s0xx_core_034;
  wire popcount27_s0xx_core_038_not;
  wire popcount27_s0xx_core_039;
  wire popcount27_s0xx_core_040;
  wire popcount27_s0xx_core_042;
  wire popcount27_s0xx_core_043;
  wire popcount27_s0xx_core_046;
  wire popcount27_s0xx_core_047;
  wire popcount27_s0xx_core_048_not;
  wire popcount27_s0xx_core_050;
  wire popcount27_s0xx_core_052;
  wire popcount27_s0xx_core_053;
  wire popcount27_s0xx_core_054;
  wire popcount27_s0xx_core_055;
  wire popcount27_s0xx_core_056;
  wire popcount27_s0xx_core_057;
  wire popcount27_s0xx_core_058;
  wire popcount27_s0xx_core_059;
  wire popcount27_s0xx_core_060;
  wire popcount27_s0xx_core_061;
  wire popcount27_s0xx_core_062;
  wire popcount27_s0xx_core_063;
  wire popcount27_s0xx_core_064;
  wire popcount27_s0xx_core_067;
  wire popcount27_s0xx_core_068;
  wire popcount27_s0xx_core_069;
  wire popcount27_s0xx_core_070;
  wire popcount27_s0xx_core_071;
  wire popcount27_s0xx_core_072;
  wire popcount27_s0xx_core_073;
  wire popcount27_s0xx_core_075;
  wire popcount27_s0xx_core_076;
  wire popcount27_s0xx_core_077;
  wire popcount27_s0xx_core_078;
  wire popcount27_s0xx_core_079;
  wire popcount27_s0xx_core_080;
  wire popcount27_s0xx_core_081;
  wire popcount27_s0xx_core_082;
  wire popcount27_s0xx_core_083;
  wire popcount27_s0xx_core_084;
  wire popcount27_s0xx_core_086;
  wire popcount27_s0xx_core_087;
  wire popcount27_s0xx_core_089;
  wire popcount27_s0xx_core_091;
  wire popcount27_s0xx_core_094;
  wire popcount27_s0xx_core_095;
  wire popcount27_s0xx_core_096;
  wire popcount27_s0xx_core_097;
  wire popcount27_s0xx_core_099;
  wire popcount27_s0xx_core_101;
  wire popcount27_s0xx_core_102;
  wire popcount27_s0xx_core_103;
  wire popcount27_s0xx_core_104;
  wire popcount27_s0xx_core_105;
  wire popcount27_s0xx_core_106;
  wire popcount27_s0xx_core_108_not;
  wire popcount27_s0xx_core_110;
  wire popcount27_s0xx_core_112;
  wire popcount27_s0xx_core_115_not;
  wire popcount27_s0xx_core_116;
  wire popcount27_s0xx_core_119;
  wire popcount27_s0xx_core_120;
  wire popcount27_s0xx_core_121;
  wire popcount27_s0xx_core_123;
  wire popcount27_s0xx_core_126;
  wire popcount27_s0xx_core_127;
  wire popcount27_s0xx_core_130;
  wire popcount27_s0xx_core_132;
  wire popcount27_s0xx_core_133;
  wire popcount27_s0xx_core_134;
  wire popcount27_s0xx_core_136_not;
  wire popcount27_s0xx_core_138;
  wire popcount27_s0xx_core_139;
  wire popcount27_s0xx_core_143;
  wire popcount27_s0xx_core_144;
  wire popcount27_s0xx_core_146;
  wire popcount27_s0xx_core_149;
  wire popcount27_s0xx_core_150;
  wire popcount27_s0xx_core_151;
  wire popcount27_s0xx_core_154;
  wire popcount27_s0xx_core_155;
  wire popcount27_s0xx_core_156;
  wire popcount27_s0xx_core_158;
  wire popcount27_s0xx_core_163;
  wire popcount27_s0xx_core_164;
  wire popcount27_s0xx_core_165;
  wire popcount27_s0xx_core_166;
  wire popcount27_s0xx_core_171;
  wire popcount27_s0xx_core_173;
  wire popcount27_s0xx_core_174;
  wire popcount27_s0xx_core_175;
  wire popcount27_s0xx_core_176;
  wire popcount27_s0xx_core_177;
  wire popcount27_s0xx_core_178;
  wire popcount27_s0xx_core_179;
  wire popcount27_s0xx_core_182;
  wire popcount27_s0xx_core_187;
  wire popcount27_s0xx_core_188;
  wire popcount27_s0xx_core_189;
  wire popcount27_s0xx_core_191;
  wire popcount27_s0xx_core_192;
  wire popcount27_s0xx_core_195;

  assign popcount27_s0xx_core_032 = ~(input_a[21] & input_a[20]);
  assign popcount27_s0xx_core_033 = input_a[7] | input_a[15];
  assign popcount27_s0xx_core_034 = input_a[18] & input_a[9];
  assign popcount27_s0xx_core_038_not = ~input_a[13];
  assign popcount27_s0xx_core_039 = ~(input_a[17] & input_a[26]);
  assign popcount27_s0xx_core_040 = ~(input_a[12] | input_a[15]);
  assign popcount27_s0xx_core_042 = input_a[15] ^ input_a[5];
  assign popcount27_s0xx_core_043 = ~(input_a[17] ^ input_a[15]);
  assign popcount27_s0xx_core_046 = ~(input_a[0] ^ input_a[3]);
  assign popcount27_s0xx_core_047 = ~(input_a[6] | input_a[25]);
  assign popcount27_s0xx_core_048_not = ~input_a[13];
  assign popcount27_s0xx_core_050 = input_a[13] ^ input_a[23];
  assign popcount27_s0xx_core_052 = ~(input_a[2] ^ input_a[16]);
  assign popcount27_s0xx_core_053 = ~(input_a[11] & input_a[24]);
  assign popcount27_s0xx_core_054 = input_a[9] ^ input_a[8];
  assign popcount27_s0xx_core_055 = input_a[26] | input_a[20];
  assign popcount27_s0xx_core_056 = input_a[21] & input_a[15];
  assign popcount27_s0xx_core_057 = ~(input_a[12] & input_a[2]);
  assign popcount27_s0xx_core_058 = ~(input_a[21] ^ input_a[12]);
  assign popcount27_s0xx_core_059 = input_a[10] & input_a[18];
  assign popcount27_s0xx_core_060 = ~(input_a[20] | input_a[26]);
  assign popcount27_s0xx_core_061 = ~(input_a[10] & input_a[3]);
  assign popcount27_s0xx_core_062 = ~(input_a[5] ^ input_a[6]);
  assign popcount27_s0xx_core_063 = input_a[10] & input_a[13];
  assign popcount27_s0xx_core_064 = input_a[20] & input_a[13];
  assign popcount27_s0xx_core_067 = input_a[14] ^ input_a[6];
  assign popcount27_s0xx_core_068 = ~(input_a[4] | input_a[16]);
  assign popcount27_s0xx_core_069 = ~(input_a[17] & input_a[13]);
  assign popcount27_s0xx_core_070 = ~(input_a[17] ^ input_a[26]);
  assign popcount27_s0xx_core_071 = ~(input_a[1] & input_a[25]);
  assign popcount27_s0xx_core_072 = ~input_a[16];
  assign popcount27_s0xx_core_073 = ~(input_a[6] | input_a[20]);
  assign popcount27_s0xx_core_075 = input_a[0] | input_a[18];
  assign popcount27_s0xx_core_076 = ~(input_a[10] | input_a[17]);
  assign popcount27_s0xx_core_077 = input_a[15] ^ input_a[2];
  assign popcount27_s0xx_core_078 = input_a[1] | input_a[10];
  assign popcount27_s0xx_core_079 = input_a[5] ^ input_a[26];
  assign popcount27_s0xx_core_080 = input_a[11] | input_a[13];
  assign popcount27_s0xx_core_081 = ~(input_a[6] & input_a[6]);
  assign popcount27_s0xx_core_082 = ~input_a[20];
  assign popcount27_s0xx_core_083 = ~input_a[18];
  assign popcount27_s0xx_core_084 = ~(input_a[6] | input_a[20]);
  assign popcount27_s0xx_core_086 = input_a[4] | input_a[20];
  assign popcount27_s0xx_core_087 = input_a[1] | input_a[5];
  assign popcount27_s0xx_core_089 = input_a[4] ^ input_a[22];
  assign popcount27_s0xx_core_091 = input_a[18] & input_a[18];
  assign popcount27_s0xx_core_094 = ~(input_a[3] ^ input_a[18]);
  assign popcount27_s0xx_core_095 = input_a[20] & input_a[0];
  assign popcount27_s0xx_core_096 = input_a[9] | input_a[16];
  assign popcount27_s0xx_core_097 = ~(input_a[24] & input_a[15]);
  assign popcount27_s0xx_core_099 = input_a[6] | input_a[4];
  assign popcount27_s0xx_core_101 = input_a[16] | input_a[7];
  assign popcount27_s0xx_core_102 = ~input_a[4];
  assign popcount27_s0xx_core_103 = ~(input_a[6] & input_a[21]);
  assign popcount27_s0xx_core_104 = input_a[24] | input_a[12];
  assign popcount27_s0xx_core_105 = input_a[5] | input_a[0];
  assign popcount27_s0xx_core_106 = input_a[3] | input_a[7];
  assign popcount27_s0xx_core_108_not = ~input_a[14];
  assign popcount27_s0xx_core_110 = ~input_a[22];
  assign popcount27_s0xx_core_112 = ~(input_a[20] ^ input_a[13]);
  assign popcount27_s0xx_core_115_not = ~input_a[20];
  assign popcount27_s0xx_core_116 = input_a[18] & input_a[23];
  assign popcount27_s0xx_core_119 = ~input_a[24];
  assign popcount27_s0xx_core_120 = input_a[9] ^ input_a[12];
  assign popcount27_s0xx_core_121 = ~(input_a[8] ^ input_a[18]);
  assign popcount27_s0xx_core_123 = input_a[4] | input_a[25];
  assign popcount27_s0xx_core_126 = ~(input_a[5] & input_a[20]);
  assign popcount27_s0xx_core_127 = input_a[16] ^ input_a[4];
  assign popcount27_s0xx_core_130 = ~input_a[18];
  assign popcount27_s0xx_core_132 = ~(input_a[11] & input_a[7]);
  assign popcount27_s0xx_core_133 = ~input_a[20];
  assign popcount27_s0xx_core_134 = input_a[21] | input_a[18];
  assign popcount27_s0xx_core_136_not = ~input_a[7];
  assign popcount27_s0xx_core_138 = input_a[25] & input_a[10];
  assign popcount27_s0xx_core_139 = ~(input_a[0] ^ input_a[26]);
  assign popcount27_s0xx_core_143 = ~(input_a[17] & input_a[21]);
  assign popcount27_s0xx_core_144 = input_a[8] & input_a[22];
  assign popcount27_s0xx_core_146 = input_a[25] ^ input_a[15];
  assign popcount27_s0xx_core_149 = ~input_a[6];
  assign popcount27_s0xx_core_150 = input_a[3] | input_a[23];
  assign popcount27_s0xx_core_151 = ~(input_a[16] & input_a[26]);
  assign popcount27_s0xx_core_154 = ~input_a[8];
  assign popcount27_s0xx_core_155 = input_a[18] | input_a[4];
  assign popcount27_s0xx_core_156 = ~(input_a[15] | input_a[4]);
  assign popcount27_s0xx_core_158 = input_a[4] ^ input_a[13];
  assign popcount27_s0xx_core_163 = input_a[1] & input_a[23];
  assign popcount27_s0xx_core_164 = input_a[1] ^ input_a[12];
  assign popcount27_s0xx_core_165 = input_a[9] & input_a[11];
  assign popcount27_s0xx_core_166 = ~(input_a[2] & input_a[0]);
  assign popcount27_s0xx_core_171 = ~(input_a[25] & input_a[5]);
  assign popcount27_s0xx_core_173 = input_a[15] & input_a[15];
  assign popcount27_s0xx_core_174 = input_a[2] & input_a[3];
  assign popcount27_s0xx_core_175 = ~(input_a[6] | input_a[0]);
  assign popcount27_s0xx_core_176 = ~(input_a[0] ^ input_a[21]);
  assign popcount27_s0xx_core_177 = ~input_a[11];
  assign popcount27_s0xx_core_178 = ~(input_a[3] | input_a[25]);
  assign popcount27_s0xx_core_179 = input_a[23] & input_a[18];
  assign popcount27_s0xx_core_182 = ~input_a[0];
  assign popcount27_s0xx_core_187 = ~(input_a[10] | input_a[5]);
  assign popcount27_s0xx_core_188 = ~(input_a[2] | input_a[8]);
  assign popcount27_s0xx_core_189 = input_a[13] ^ input_a[9];
  assign popcount27_s0xx_core_191 = input_a[20] & input_a[20];
  assign popcount27_s0xx_core_192 = input_a[3] ^ input_a[12];
  assign popcount27_s0xx_core_195 = input_a[26] & input_a[8];

  assign popcount27_s0xx_out[0] = input_a[3];
  assign popcount27_s0xx_out[1] = input_a[0];
  assign popcount27_s0xx_out[2] = 1'b1;
  assign popcount27_s0xx_out[3] = input_a[10];
  assign popcount27_s0xx_out[4] = 1'b0;
endmodule