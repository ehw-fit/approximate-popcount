// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.69417
// WCE=21.0
// EP=0.953061%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_35id(input [31:0] input_a, output [5:0] popcount32_35id_out);
  wire popcount32_35id_core_034_not;
  wire popcount32_35id_core_035;
  wire popcount32_35id_core_036;
  wire popcount32_35id_core_037;
  wire popcount32_35id_core_038;
  wire popcount32_35id_core_040;
  wire popcount32_35id_core_041;
  wire popcount32_35id_core_042;
  wire popcount32_35id_core_043;
  wire popcount32_35id_core_047;
  wire popcount32_35id_core_048;
  wire popcount32_35id_core_049;
  wire popcount32_35id_core_050;
  wire popcount32_35id_core_052_not;
  wire popcount32_35id_core_055;
  wire popcount32_35id_core_056;
  wire popcount32_35id_core_057;
  wire popcount32_35id_core_059;
  wire popcount32_35id_core_060;
  wire popcount32_35id_core_062;
  wire popcount32_35id_core_064;
  wire popcount32_35id_core_065;
  wire popcount32_35id_core_068;
  wire popcount32_35id_core_069;
  wire popcount32_35id_core_070;
  wire popcount32_35id_core_071;
  wire popcount32_35id_core_072;
  wire popcount32_35id_core_073;
  wire popcount32_35id_core_074;
  wire popcount32_35id_core_076;
  wire popcount32_35id_core_077;
  wire popcount32_35id_core_080;
  wire popcount32_35id_core_081;
  wire popcount32_35id_core_082;
  wire popcount32_35id_core_083;
  wire popcount32_35id_core_085;
  wire popcount32_35id_core_087;
  wire popcount32_35id_core_088;
  wire popcount32_35id_core_090;
  wire popcount32_35id_core_091;
  wire popcount32_35id_core_092;
  wire popcount32_35id_core_093;
  wire popcount32_35id_core_094;
  wire popcount32_35id_core_096;
  wire popcount32_35id_core_099;
  wire popcount32_35id_core_100_not;
  wire popcount32_35id_core_104;
  wire popcount32_35id_core_105;
  wire popcount32_35id_core_106;
  wire popcount32_35id_core_107;
  wire popcount32_35id_core_109;
  wire popcount32_35id_core_110;
  wire popcount32_35id_core_111;
  wire popcount32_35id_core_114;
  wire popcount32_35id_core_115;
  wire popcount32_35id_core_116;
  wire popcount32_35id_core_117;
  wire popcount32_35id_core_118;
  wire popcount32_35id_core_119;
  wire popcount32_35id_core_120;
  wire popcount32_35id_core_121;
  wire popcount32_35id_core_125;
  wire popcount32_35id_core_127;
  wire popcount32_35id_core_128;
  wire popcount32_35id_core_129;
  wire popcount32_35id_core_132_not;
  wire popcount32_35id_core_133;
  wire popcount32_35id_core_134;
  wire popcount32_35id_core_135;
  wire popcount32_35id_core_136;
  wire popcount32_35id_core_137;
  wire popcount32_35id_core_138;
  wire popcount32_35id_core_141;
  wire popcount32_35id_core_142;
  wire popcount32_35id_core_144;
  wire popcount32_35id_core_145;
  wire popcount32_35id_core_146;
  wire popcount32_35id_core_147;
  wire popcount32_35id_core_148;
  wire popcount32_35id_core_149;
  wire popcount32_35id_core_151;
  wire popcount32_35id_core_152;
  wire popcount32_35id_core_154;
  wire popcount32_35id_core_155;
  wire popcount32_35id_core_156;
  wire popcount32_35id_core_158;
  wire popcount32_35id_core_160;
  wire popcount32_35id_core_161;
  wire popcount32_35id_core_163;
  wire popcount32_35id_core_164;
  wire popcount32_35id_core_165;
  wire popcount32_35id_core_166;
  wire popcount32_35id_core_167;
  wire popcount32_35id_core_168;
  wire popcount32_35id_core_169;
  wire popcount32_35id_core_172;
  wire popcount32_35id_core_173;
  wire popcount32_35id_core_174;
  wire popcount32_35id_core_176;
  wire popcount32_35id_core_177;
  wire popcount32_35id_core_178;
  wire popcount32_35id_core_180;
  wire popcount32_35id_core_182;
  wire popcount32_35id_core_183;
  wire popcount32_35id_core_184_not;
  wire popcount32_35id_core_185;
  wire popcount32_35id_core_186;
  wire popcount32_35id_core_187;
  wire popcount32_35id_core_188;
  wire popcount32_35id_core_190;
  wire popcount32_35id_core_191;
  wire popcount32_35id_core_192;
  wire popcount32_35id_core_194;
  wire popcount32_35id_core_196;
  wire popcount32_35id_core_197;
  wire popcount32_35id_core_199;
  wire popcount32_35id_core_200;
  wire popcount32_35id_core_201;
  wire popcount32_35id_core_202;
  wire popcount32_35id_core_205;
  wire popcount32_35id_core_208;
  wire popcount32_35id_core_209;
  wire popcount32_35id_core_212;
  wire popcount32_35id_core_213;
  wire popcount32_35id_core_214;
  wire popcount32_35id_core_216;
  wire popcount32_35id_core_217;
  wire popcount32_35id_core_218;
  wire popcount32_35id_core_219;
  wire popcount32_35id_core_220;
  wire popcount32_35id_core_221;
  wire popcount32_35id_core_222;
  wire popcount32_35id_core_223;
  wire popcount32_35id_core_224;
  wire popcount32_35id_core_225;

  assign popcount32_35id_core_034_not = ~input_a[28];
  assign popcount32_35id_core_035 = input_a[1] & input_a[6];
  assign popcount32_35id_core_036 = ~input_a[7];
  assign popcount32_35id_core_037 = ~(input_a[3] | input_a[9]);
  assign popcount32_35id_core_038 = input_a[22] & input_a[26];
  assign popcount32_35id_core_040 = ~(input_a[30] | input_a[17]);
  assign popcount32_35id_core_041 = ~(input_a[21] | input_a[7]);
  assign popcount32_35id_core_042 = input_a[5] & input_a[16];
  assign popcount32_35id_core_043 = input_a[1] | input_a[28];
  assign popcount32_35id_core_047 = ~(input_a[11] ^ input_a[6]);
  assign popcount32_35id_core_048 = ~(input_a[3] & input_a[6]);
  assign popcount32_35id_core_049 = ~(input_a[6] & input_a[12]);
  assign popcount32_35id_core_050 = ~(input_a[31] ^ input_a[31]);
  assign popcount32_35id_core_052_not = ~input_a[7];
  assign popcount32_35id_core_055 = ~(input_a[4] & input_a[22]);
  assign popcount32_35id_core_056 = ~input_a[30];
  assign popcount32_35id_core_057 = input_a[22] & input_a[15];
  assign popcount32_35id_core_059 = ~(input_a[25] ^ input_a[25]);
  assign popcount32_35id_core_060 = ~input_a[22];
  assign popcount32_35id_core_062 = ~(input_a[10] ^ input_a[21]);
  assign popcount32_35id_core_064 = ~(input_a[27] | input_a[3]);
  assign popcount32_35id_core_065 = input_a[14] & input_a[23];
  assign popcount32_35id_core_068 = ~(input_a[27] ^ input_a[19]);
  assign popcount32_35id_core_069 = input_a[22] & input_a[17];
  assign popcount32_35id_core_070 = ~(input_a[11] ^ input_a[4]);
  assign popcount32_35id_core_071 = ~(input_a[12] ^ input_a[16]);
  assign popcount32_35id_core_072 = input_a[25] | input_a[4];
  assign popcount32_35id_core_073 = ~(input_a[17] ^ input_a[8]);
  assign popcount32_35id_core_074 = input_a[5] ^ input_a[3];
  assign popcount32_35id_core_076 = input_a[27] & input_a[29];
  assign popcount32_35id_core_077 = input_a[24] & input_a[1];
  assign popcount32_35id_core_080 = ~(input_a[9] & input_a[24]);
  assign popcount32_35id_core_081 = ~(input_a[9] | input_a[6]);
  assign popcount32_35id_core_082 = ~input_a[7];
  assign popcount32_35id_core_083 = input_a[5] & input_a[0];
  assign popcount32_35id_core_085 = input_a[6] ^ input_a[20];
  assign popcount32_35id_core_087 = input_a[4] ^ input_a[30];
  assign popcount32_35id_core_088 = ~input_a[25];
  assign popcount32_35id_core_090 = input_a[3] | input_a[23];
  assign popcount32_35id_core_091 = ~(input_a[9] | input_a[27]);
  assign popcount32_35id_core_092 = ~(input_a[24] & input_a[14]);
  assign popcount32_35id_core_093 = input_a[7] | input_a[26];
  assign popcount32_35id_core_094 = ~(input_a[7] | input_a[25]);
  assign popcount32_35id_core_096 = ~(input_a[27] ^ input_a[0]);
  assign popcount32_35id_core_099 = ~(input_a[10] ^ input_a[17]);
  assign popcount32_35id_core_100_not = ~input_a[31];
  assign popcount32_35id_core_104 = input_a[30] | input_a[10];
  assign popcount32_35id_core_105 = input_a[23] | input_a[2];
  assign popcount32_35id_core_106 = input_a[22] | input_a[9];
  assign popcount32_35id_core_107 = ~input_a[2];
  assign popcount32_35id_core_109 = ~input_a[7];
  assign popcount32_35id_core_110 = input_a[23] | input_a[12];
  assign popcount32_35id_core_111 = input_a[15] & input_a[3];
  assign popcount32_35id_core_114 = input_a[23] | input_a[1];
  assign popcount32_35id_core_115 = ~input_a[9];
  assign popcount32_35id_core_116 = input_a[6] & input_a[18];
  assign popcount32_35id_core_117 = ~(input_a[30] | input_a[7]);
  assign popcount32_35id_core_118 = ~(input_a[9] | input_a[21]);
  assign popcount32_35id_core_119 = ~(input_a[21] & input_a[23]);
  assign popcount32_35id_core_120 = ~(input_a[17] | input_a[30]);
  assign popcount32_35id_core_121 = input_a[3] & input_a[16];
  assign popcount32_35id_core_125 = ~(input_a[12] ^ input_a[18]);
  assign popcount32_35id_core_127 = ~(input_a[13] & input_a[24]);
  assign popcount32_35id_core_128 = ~(input_a[29] | input_a[6]);
  assign popcount32_35id_core_129 = input_a[9] | input_a[3];
  assign popcount32_35id_core_132_not = ~input_a[31];
  assign popcount32_35id_core_133 = ~(input_a[7] ^ input_a[21]);
  assign popcount32_35id_core_134 = ~input_a[23];
  assign popcount32_35id_core_135 = ~(input_a[11] & input_a[13]);
  assign popcount32_35id_core_136 = ~(input_a[27] | input_a[13]);
  assign popcount32_35id_core_137 = ~input_a[0];
  assign popcount32_35id_core_138 = input_a[23] ^ input_a[19];
  assign popcount32_35id_core_141 = input_a[18] ^ input_a[20];
  assign popcount32_35id_core_142 = input_a[21] | input_a[7];
  assign popcount32_35id_core_144 = ~(input_a[18] ^ input_a[23]);
  assign popcount32_35id_core_145 = ~(input_a[6] | input_a[9]);
  assign popcount32_35id_core_146 = ~(input_a[22] & input_a[24]);
  assign popcount32_35id_core_147 = input_a[25] & input_a[13];
  assign popcount32_35id_core_148 = input_a[6] ^ input_a[20];
  assign popcount32_35id_core_149 = input_a[6] & input_a[30];
  assign popcount32_35id_core_151 = input_a[15] & input_a[19];
  assign popcount32_35id_core_152 = input_a[2] & input_a[17];
  assign popcount32_35id_core_154 = ~(input_a[25] | input_a[11]);
  assign popcount32_35id_core_155 = ~(input_a[19] | input_a[12]);
  assign popcount32_35id_core_156 = ~(input_a[15] ^ input_a[4]);
  assign popcount32_35id_core_158 = ~(input_a[1] & input_a[26]);
  assign popcount32_35id_core_160 = input_a[10] | input_a[5];
  assign popcount32_35id_core_161 = ~input_a[22];
  assign popcount32_35id_core_163 = input_a[8] | input_a[30];
  assign popcount32_35id_core_164 = input_a[13] & input_a[16];
  assign popcount32_35id_core_165 = ~input_a[8];
  assign popcount32_35id_core_166 = ~(input_a[11] | input_a[26]);
  assign popcount32_35id_core_167 = ~(input_a[19] | input_a[30]);
  assign popcount32_35id_core_168 = input_a[12] | input_a[15];
  assign popcount32_35id_core_169 = ~(input_a[29] & input_a[21]);
  assign popcount32_35id_core_172 = ~(input_a[25] | input_a[27]);
  assign popcount32_35id_core_173 = ~(input_a[30] ^ input_a[4]);
  assign popcount32_35id_core_174 = input_a[11] ^ input_a[27];
  assign popcount32_35id_core_176 = ~(input_a[19] & input_a[7]);
  assign popcount32_35id_core_177 = ~input_a[20];
  assign popcount32_35id_core_178 = input_a[28] & input_a[18];
  assign popcount32_35id_core_180 = ~(input_a[25] & input_a[2]);
  assign popcount32_35id_core_182 = input_a[19] ^ input_a[13];
  assign popcount32_35id_core_183 = ~(input_a[28] | input_a[19]);
  assign popcount32_35id_core_184_not = ~input_a[30];
  assign popcount32_35id_core_185 = input_a[11] ^ input_a[26];
  assign popcount32_35id_core_186 = ~(input_a[28] & input_a[0]);
  assign popcount32_35id_core_187 = ~(input_a[26] | input_a[24]);
  assign popcount32_35id_core_188 = input_a[7] | input_a[3];
  assign popcount32_35id_core_190 = ~(input_a[30] ^ input_a[6]);
  assign popcount32_35id_core_191 = ~(input_a[11] ^ input_a[20]);
  assign popcount32_35id_core_192 = ~(input_a[24] ^ input_a[7]);
  assign popcount32_35id_core_194 = ~input_a[26];
  assign popcount32_35id_core_196 = input_a[26] | input_a[30];
  assign popcount32_35id_core_197 = input_a[18] ^ input_a[19];
  assign popcount32_35id_core_199 = ~(input_a[10] ^ input_a[1]);
  assign popcount32_35id_core_200 = ~input_a[26];
  assign popcount32_35id_core_201 = input_a[17] & input_a[1];
  assign popcount32_35id_core_202 = ~(input_a[1] | input_a[21]);
  assign popcount32_35id_core_205 = ~input_a[13];
  assign popcount32_35id_core_208 = ~(input_a[28] | input_a[9]);
  assign popcount32_35id_core_209 = ~(input_a[27] & input_a[13]);
  assign popcount32_35id_core_212 = input_a[9] & input_a[10];
  assign popcount32_35id_core_213 = ~(input_a[15] ^ input_a[22]);
  assign popcount32_35id_core_214 = ~(input_a[12] ^ input_a[24]);
  assign popcount32_35id_core_216 = input_a[12] ^ input_a[14];
  assign popcount32_35id_core_217 = ~(input_a[25] | input_a[13]);
  assign popcount32_35id_core_218 = ~(input_a[12] & input_a[21]);
  assign popcount32_35id_core_219 = ~(input_a[22] | input_a[9]);
  assign popcount32_35id_core_220 = ~(input_a[11] | input_a[26]);
  assign popcount32_35id_core_221 = ~(input_a[22] | input_a[6]);
  assign popcount32_35id_core_222 = input_a[25] | input_a[16];
  assign popcount32_35id_core_223 = ~(input_a[7] | input_a[29]);
  assign popcount32_35id_core_224 = input_a[27] | input_a[29];
  assign popcount32_35id_core_225 = ~input_a[13];

  assign popcount32_35id_out[0] = input_a[21];
  assign popcount32_35id_out[1] = input_a[31];
  assign popcount32_35id_out[2] = input_a[23];
  assign popcount32_35id_out[3] = 1'b1;
  assign popcount32_35id_out[4] = 1'b0;
  assign popcount32_35id_out[5] = 1'b0;
endmodule