// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.41218
// WCE=17.0
// EP=0.994043%
// Printed PDK parameters:
//  Area=28944668.0
//  Delay=44634204.0
//  Power=1472400.0

module popcount33_w6o5(input [32:0] input_a, output [5:0] popcount33_w6o5_out);
  wire popcount33_w6o5_core_035;
  wire popcount33_w6o5_core_036;
  wire popcount33_w6o5_core_037;
  wire popcount33_w6o5_core_038;
  wire popcount33_w6o5_core_040;
  wire popcount33_w6o5_core_041;
  wire popcount33_w6o5_core_042;
  wire popcount33_w6o5_core_043;
  wire popcount33_w6o5_core_044;
  wire popcount33_w6o5_core_046;
  wire popcount33_w6o5_core_047;
  wire popcount33_w6o5_core_048;
  wire popcount33_w6o5_core_049;
  wire popcount33_w6o5_core_050;
  wire popcount33_w6o5_core_051;
  wire popcount33_w6o5_core_052;
  wire popcount33_w6o5_core_053;
  wire popcount33_w6o5_core_054;
  wire popcount33_w6o5_core_057;
  wire popcount33_w6o5_core_058;
  wire popcount33_w6o5_core_059;
  wire popcount33_w6o5_core_060;
  wire popcount33_w6o5_core_062;
  wire popcount33_w6o5_core_064;
  wire popcount33_w6o5_core_065;
  wire popcount33_w6o5_core_066;
  wire popcount33_w6o5_core_067;
  wire popcount33_w6o5_core_069;
  wire popcount33_w6o5_core_070;
  wire popcount33_w6o5_core_071;
  wire popcount33_w6o5_core_072;
  wire popcount33_w6o5_core_073;
  wire popcount33_w6o5_core_074;
  wire popcount33_w6o5_core_075;
  wire popcount33_w6o5_core_076;
  wire popcount33_w6o5_core_077;
  wire popcount33_w6o5_core_078;
  wire popcount33_w6o5_core_080;
  wire popcount33_w6o5_core_081;
  wire popcount33_w6o5_core_083;
  wire popcount33_w6o5_core_084;
  wire popcount33_w6o5_core_085;
  wire popcount33_w6o5_core_087;
  wire popcount33_w6o5_core_089;
  wire popcount33_w6o5_core_090;
  wire popcount33_w6o5_core_091;
  wire popcount33_w6o5_core_092;
  wire popcount33_w6o5_core_093;
  wire popcount33_w6o5_core_094;
  wire popcount33_w6o5_core_095;
  wire popcount33_w6o5_core_096;
  wire popcount33_w6o5_core_097;
  wire popcount33_w6o5_core_099;
  wire popcount33_w6o5_core_100;
  wire popcount33_w6o5_core_103;
  wire popcount33_w6o5_core_104;
  wire popcount33_w6o5_core_105;
  wire popcount33_w6o5_core_106;
  wire popcount33_w6o5_core_108;
  wire popcount33_w6o5_core_110;
  wire popcount33_w6o5_core_111;
  wire popcount33_w6o5_core_112;
  wire popcount33_w6o5_core_113;
  wire popcount33_w6o5_core_114;
  wire popcount33_w6o5_core_116;
  wire popcount33_w6o5_core_117;
  wire popcount33_w6o5_core_121;
  wire popcount33_w6o5_core_122;
  wire popcount33_w6o5_core_124;
  wire popcount33_w6o5_core_125;
  wire popcount33_w6o5_core_128;
  wire popcount33_w6o5_core_129;
  wire popcount33_w6o5_core_131;
  wire popcount33_w6o5_core_132;
  wire popcount33_w6o5_core_133;
  wire popcount33_w6o5_core_134;
  wire popcount33_w6o5_core_135;
  wire popcount33_w6o5_core_137;
  wire popcount33_w6o5_core_138;
  wire popcount33_w6o5_core_141;
  wire popcount33_w6o5_core_142_not;
  wire popcount33_w6o5_core_145;
  wire popcount33_w6o5_core_149;
  wire popcount33_w6o5_core_150;
  wire popcount33_w6o5_core_152;
  wire popcount33_w6o5_core_153;
  wire popcount33_w6o5_core_154;
  wire popcount33_w6o5_core_156;
  wire popcount33_w6o5_core_157;
  wire popcount33_w6o5_core_158;
  wire popcount33_w6o5_core_159;
  wire popcount33_w6o5_core_160;
  wire popcount33_w6o5_core_161;
  wire popcount33_w6o5_core_163;
  wire popcount33_w6o5_core_165;
  wire popcount33_w6o5_core_168;
  wire popcount33_w6o5_core_169;
  wire popcount33_w6o5_core_170;
  wire popcount33_w6o5_core_171;
  wire popcount33_w6o5_core_172;
  wire popcount33_w6o5_core_173;
  wire popcount33_w6o5_core_174;
  wire popcount33_w6o5_core_176;
  wire popcount33_w6o5_core_178;
  wire popcount33_w6o5_core_179;
  wire popcount33_w6o5_core_181;
  wire popcount33_w6o5_core_183;
  wire popcount33_w6o5_core_184;
  wire popcount33_w6o5_core_185;
  wire popcount33_w6o5_core_188;
  wire popcount33_w6o5_core_189;
  wire popcount33_w6o5_core_190;
  wire popcount33_w6o5_core_191;
  wire popcount33_w6o5_core_192;
  wire popcount33_w6o5_core_193;
  wire popcount33_w6o5_core_195;
  wire popcount33_w6o5_core_196;
  wire popcount33_w6o5_core_197;
  wire popcount33_w6o5_core_198;
  wire popcount33_w6o5_core_199;
  wire popcount33_w6o5_core_200;
  wire popcount33_w6o5_core_201;
  wire popcount33_w6o5_core_202;
  wire popcount33_w6o5_core_203;
  wire popcount33_w6o5_core_204_not;
  wire popcount33_w6o5_core_205;
  wire popcount33_w6o5_core_206;
  wire popcount33_w6o5_core_207;
  wire popcount33_w6o5_core_210;
  wire popcount33_w6o5_core_211;
  wire popcount33_w6o5_core_212;
  wire popcount33_w6o5_core_214;
  wire popcount33_w6o5_core_215;
  wire popcount33_w6o5_core_216;
  wire popcount33_w6o5_core_217;
  wire popcount33_w6o5_core_220;
  wire popcount33_w6o5_core_224;
  wire popcount33_w6o5_core_225;
  wire popcount33_w6o5_core_229;
  wire popcount33_w6o5_core_230;
  wire popcount33_w6o5_core_232;
  wire popcount33_w6o5_core_233;
  wire popcount33_w6o5_core_234;
  wire popcount33_w6o5_core_235;
  wire popcount33_w6o5_core_236;
  wire popcount33_w6o5_core_238;

  assign popcount33_w6o5_core_035 = input_a[25] | input_a[1];
  assign popcount33_w6o5_core_036 = input_a[26] & input_a[22];
  assign popcount33_w6o5_core_037 = input_a[2] ^ input_a[3];
  assign popcount33_w6o5_core_038 = input_a[2] & input_a[3];
  assign popcount33_w6o5_core_040 = input_a[30] & popcount33_w6o5_core_037;
  assign popcount33_w6o5_core_041 = popcount33_w6o5_core_036 ^ popcount33_w6o5_core_038;
  assign popcount33_w6o5_core_042 = popcount33_w6o5_core_036 & popcount33_w6o5_core_038;
  assign popcount33_w6o5_core_043 = popcount33_w6o5_core_041 | popcount33_w6o5_core_040;
  assign popcount33_w6o5_core_044 = input_a[4] & input_a[18];
  assign popcount33_w6o5_core_046 = input_a[15] & input_a[8];
  assign popcount33_w6o5_core_047 = input_a[25] & input_a[14];
  assign popcount33_w6o5_core_048 = input_a[6] ^ input_a[7];
  assign popcount33_w6o5_core_049 = input_a[6] & input_a[7];
  assign popcount33_w6o5_core_050 = input_a[4] ^ input_a[29];
  assign popcount33_w6o5_core_051 = input_a[28] & popcount33_w6o5_core_048;
  assign popcount33_w6o5_core_052 = popcount33_w6o5_core_047 ^ popcount33_w6o5_core_049;
  assign popcount33_w6o5_core_053 = popcount33_w6o5_core_047 & popcount33_w6o5_core_049;
  assign popcount33_w6o5_core_054 = popcount33_w6o5_core_052 | popcount33_w6o5_core_051;
  assign popcount33_w6o5_core_057 = ~(input_a[18] | input_a[5]);
  assign popcount33_w6o5_core_058 = ~(input_a[22] ^ input_a[16]);
  assign popcount33_w6o5_core_059 = popcount33_w6o5_core_043 ^ popcount33_w6o5_core_054;
  assign popcount33_w6o5_core_060 = popcount33_w6o5_core_043 & popcount33_w6o5_core_054;
  assign popcount33_w6o5_core_062 = ~(input_a[23] & input_a[31]);
  assign popcount33_w6o5_core_064 = popcount33_w6o5_core_042 ^ popcount33_w6o5_core_053;
  assign popcount33_w6o5_core_065 = popcount33_w6o5_core_042 & popcount33_w6o5_core_053;
  assign popcount33_w6o5_core_066 = popcount33_w6o5_core_064 | popcount33_w6o5_core_060;
  assign popcount33_w6o5_core_067 = input_a[29] & input_a[3];
  assign popcount33_w6o5_core_069 = input_a[8] ^ input_a[9];
  assign popcount33_w6o5_core_070 = input_a[8] & input_a[9];
  assign popcount33_w6o5_core_071 = input_a[10] ^ input_a[11];
  assign popcount33_w6o5_core_072 = input_a[10] & input_a[11];
  assign popcount33_w6o5_core_073 = popcount33_w6o5_core_069 ^ popcount33_w6o5_core_071;
  assign popcount33_w6o5_core_074 = popcount33_w6o5_core_069 & popcount33_w6o5_core_071;
  assign popcount33_w6o5_core_075 = popcount33_w6o5_core_070 ^ popcount33_w6o5_core_072;
  assign popcount33_w6o5_core_076 = popcount33_w6o5_core_070 & popcount33_w6o5_core_072;
  assign popcount33_w6o5_core_077 = popcount33_w6o5_core_075 | popcount33_w6o5_core_074;
  assign popcount33_w6o5_core_078 = ~input_a[17];
  assign popcount33_w6o5_core_080 = ~(input_a[24] & input_a[26]);
  assign popcount33_w6o5_core_081 = input_a[19] & input_a[5];
  assign popcount33_w6o5_core_083 = input_a[18] | input_a[21];
  assign popcount33_w6o5_core_084 = ~input_a[11];
  assign popcount33_w6o5_core_085 = input_a[26] | input_a[22];
  assign popcount33_w6o5_core_087 = ~(input_a[0] ^ input_a[7]);
  assign popcount33_w6o5_core_089 = ~input_a[5];
  assign popcount33_w6o5_core_090 = ~(input_a[16] ^ input_a[14]);
  assign popcount33_w6o5_core_091 = ~(input_a[9] ^ input_a[21]);
  assign popcount33_w6o5_core_092 = popcount33_w6o5_core_073 & input_a[16];
  assign popcount33_w6o5_core_093 = popcount33_w6o5_core_077 ^ popcount33_w6o5_core_081;
  assign popcount33_w6o5_core_094 = popcount33_w6o5_core_077 & popcount33_w6o5_core_081;
  assign popcount33_w6o5_core_095 = popcount33_w6o5_core_093 ^ popcount33_w6o5_core_092;
  assign popcount33_w6o5_core_096 = popcount33_w6o5_core_093 & popcount33_w6o5_core_092;
  assign popcount33_w6o5_core_097 = popcount33_w6o5_core_094 | popcount33_w6o5_core_096;
  assign popcount33_w6o5_core_099 = input_a[8] & input_a[1];
  assign popcount33_w6o5_core_100 = popcount33_w6o5_core_076 | popcount33_w6o5_core_097;
  assign popcount33_w6o5_core_103 = ~(input_a[29] ^ input_a[11]);
  assign popcount33_w6o5_core_104 = ~input_a[10];
  assign popcount33_w6o5_core_105 = popcount33_w6o5_core_059 ^ popcount33_w6o5_core_095;
  assign popcount33_w6o5_core_106 = popcount33_w6o5_core_059 & popcount33_w6o5_core_095;
  assign popcount33_w6o5_core_108 = input_a[20] & input_a[14];
  assign popcount33_w6o5_core_110 = popcount33_w6o5_core_066 ^ popcount33_w6o5_core_100;
  assign popcount33_w6o5_core_111 = popcount33_w6o5_core_066 & popcount33_w6o5_core_100;
  assign popcount33_w6o5_core_112 = popcount33_w6o5_core_110 ^ popcount33_w6o5_core_106;
  assign popcount33_w6o5_core_113 = popcount33_w6o5_core_110 & popcount33_w6o5_core_106;
  assign popcount33_w6o5_core_114 = popcount33_w6o5_core_111 | popcount33_w6o5_core_113;
  assign popcount33_w6o5_core_116 = ~(input_a[11] | input_a[11]);
  assign popcount33_w6o5_core_117 = popcount33_w6o5_core_065 | popcount33_w6o5_core_114;
  assign popcount33_w6o5_core_121 = input_a[25] & input_a[23];
  assign popcount33_w6o5_core_122 = input_a[4] ^ input_a[23];
  assign popcount33_w6o5_core_124 = input_a[13] | input_a[30];
  assign popcount33_w6o5_core_125 = ~(input_a[27] | input_a[32]);
  assign popcount33_w6o5_core_128 = ~(input_a[24] ^ input_a[18]);
  assign popcount33_w6o5_core_129 = ~(input_a[10] ^ input_a[4]);
  assign popcount33_w6o5_core_131 = ~(input_a[8] ^ input_a[31]);
  assign popcount33_w6o5_core_132 = ~(input_a[5] ^ input_a[11]);
  assign popcount33_w6o5_core_133 = ~(input_a[13] | input_a[25]);
  assign popcount33_w6o5_core_134 = input_a[24] ^ input_a[12];
  assign popcount33_w6o5_core_135 = ~(input_a[7] ^ input_a[16]);
  assign popcount33_w6o5_core_137 = ~input_a[30];
  assign popcount33_w6o5_core_138 = ~input_a[2];
  assign popcount33_w6o5_core_141 = ~(input_a[8] & input_a[14]);
  assign popcount33_w6o5_core_142_not = ~input_a[14];
  assign popcount33_w6o5_core_145 = input_a[30] | input_a[7];
  assign popcount33_w6o5_core_149 = ~(input_a[27] ^ input_a[17]);
  assign popcount33_w6o5_core_150 = input_a[31] & input_a[7];
  assign popcount33_w6o5_core_152 = ~input_a[6];
  assign popcount33_w6o5_core_153 = input_a[11] | input_a[4];
  assign popcount33_w6o5_core_154 = input_a[7] & input_a[3];
  assign popcount33_w6o5_core_156 = ~(input_a[28] ^ input_a[6]);
  assign popcount33_w6o5_core_157 = ~(input_a[20] | input_a[5]);
  assign popcount33_w6o5_core_158 = ~input_a[17];
  assign popcount33_w6o5_core_159 = input_a[22] ^ input_a[18];
  assign popcount33_w6o5_core_160 = ~input_a[16];
  assign popcount33_w6o5_core_161 = ~input_a[31];
  assign popcount33_w6o5_core_163 = input_a[16] ^ input_a[16];
  assign popcount33_w6o5_core_165 = ~(input_a[18] | input_a[13]);
  assign popcount33_w6o5_core_168 = input_a[20] ^ input_a[1];
  assign popcount33_w6o5_core_169 = input_a[7] ^ input_a[9];
  assign popcount33_w6o5_core_170 = input_a[11] & input_a[29];
  assign popcount33_w6o5_core_171 = ~(input_a[2] & input_a[32]);
  assign popcount33_w6o5_core_172 = input_a[20] ^ input_a[19];
  assign popcount33_w6o5_core_173 = ~(input_a[13] & input_a[30]);
  assign popcount33_w6o5_core_174 = ~(input_a[11] ^ input_a[10]);
  assign popcount33_w6o5_core_176 = ~(input_a[32] & input_a[21]);
  assign popcount33_w6o5_core_178 = ~input_a[20];
  assign popcount33_w6o5_core_179 = ~(input_a[0] | input_a[32]);
  assign popcount33_w6o5_core_181 = input_a[13] & input_a[17];
  assign popcount33_w6o5_core_183 = input_a[4] ^ input_a[6];
  assign popcount33_w6o5_core_184 = ~(input_a[28] & input_a[29]);
  assign popcount33_w6o5_core_185 = input_a[11] & input_a[9];
  assign popcount33_w6o5_core_188 = ~input_a[13];
  assign popcount33_w6o5_core_189 = input_a[15] ^ input_a[10];
  assign popcount33_w6o5_core_190 = ~input_a[6];
  assign popcount33_w6o5_core_191 = ~(input_a[8] & input_a[9]);
  assign popcount33_w6o5_core_192 = input_a[29] | input_a[19];
  assign popcount33_w6o5_core_193 = ~(input_a[12] | input_a[25]);
  assign popcount33_w6o5_core_195 = popcount33_w6o5_core_181 & input_a[21];
  assign popcount33_w6o5_core_196 = ~input_a[28];
  assign popcount33_w6o5_core_197 = ~(input_a[11] ^ input_a[2]);
  assign popcount33_w6o5_core_198 = input_a[1] | input_a[7];
  assign popcount33_w6o5_core_199 = ~(input_a[29] ^ input_a[14]);
  assign popcount33_w6o5_core_200 = input_a[12] & input_a[2];
  assign popcount33_w6o5_core_201 = input_a[20] ^ input_a[28];
  assign popcount33_w6o5_core_202 = input_a[2] ^ input_a[7];
  assign popcount33_w6o5_core_203 = ~(input_a[26] ^ input_a[2]);
  assign popcount33_w6o5_core_204_not = ~input_a[2];
  assign popcount33_w6o5_core_205 = ~input_a[15];
  assign popcount33_w6o5_core_206 = ~(input_a[26] | input_a[15]);
  assign popcount33_w6o5_core_207 = ~input_a[14];
  assign popcount33_w6o5_core_210 = input_a[23] ^ input_a[6];
  assign popcount33_w6o5_core_211 = input_a[12] ^ input_a[11];
  assign popcount33_w6o5_core_212 = ~input_a[25];
  assign popcount33_w6o5_core_214 = ~(input_a[4] ^ input_a[23]);
  assign popcount33_w6o5_core_215 = input_a[16] | input_a[6];
  assign popcount33_w6o5_core_216 = ~(input_a[25] | input_a[31]);
  assign popcount33_w6o5_core_217 = ~(input_a[12] ^ input_a[12]);
  assign popcount33_w6o5_core_220 = ~(input_a[19] | input_a[18]);
  assign popcount33_w6o5_core_224 = popcount33_w6o5_core_112 ^ popcount33_w6o5_core_105;
  assign popcount33_w6o5_core_225 = popcount33_w6o5_core_112 & popcount33_w6o5_core_105;
  assign popcount33_w6o5_core_229 = popcount33_w6o5_core_117 ^ popcount33_w6o5_core_225;
  assign popcount33_w6o5_core_230 = popcount33_w6o5_core_117 & popcount33_w6o5_core_225;
  assign popcount33_w6o5_core_232 = input_a[15] | popcount33_w6o5_core_195;
  assign popcount33_w6o5_core_233 = input_a[18] | input_a[7];
  assign popcount33_w6o5_core_234 = popcount33_w6o5_core_232 ^ popcount33_w6o5_core_230;
  assign popcount33_w6o5_core_235 = popcount33_w6o5_core_232 & popcount33_w6o5_core_230;
  assign popcount33_w6o5_core_236 = input_a[13] ^ input_a[14];
  assign popcount33_w6o5_core_238 = ~(input_a[19] & input_a[14]);

  assign popcount33_w6o5_out[0] = input_a[31];
  assign popcount33_w6o5_out[1] = popcount33_w6o5_core_205;
  assign popcount33_w6o5_out[2] = popcount33_w6o5_core_224;
  assign popcount33_w6o5_out[3] = popcount33_w6o5_core_229;
  assign popcount33_w6o5_out[4] = popcount33_w6o5_core_234;
  assign popcount33_w6o5_out[5] = popcount33_w6o5_core_235;
endmodule