// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.50915
// WCE=19.0
// EP=0.87489%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_ay4z(input [35:0] input_a, output [5:0] popcount36_ay4z_out);
  wire popcount36_ay4z_core_039;
  wire popcount36_ay4z_core_040;
  wire popcount36_ay4z_core_041;
  wire popcount36_ay4z_core_043;
  wire popcount36_ay4z_core_045;
  wire popcount36_ay4z_core_046;
  wire popcount36_ay4z_core_048;
  wire popcount36_ay4z_core_050;
  wire popcount36_ay4z_core_051;
  wire popcount36_ay4z_core_052;
  wire popcount36_ay4z_core_054;
  wire popcount36_ay4z_core_059;
  wire popcount36_ay4z_core_061;
  wire popcount36_ay4z_core_062;
  wire popcount36_ay4z_core_063;
  wire popcount36_ay4z_core_064;
  wire popcount36_ay4z_core_065;
  wire popcount36_ay4z_core_068;
  wire popcount36_ay4z_core_069;
  wire popcount36_ay4z_core_073;
  wire popcount36_ay4z_core_075;
  wire popcount36_ay4z_core_077;
  wire popcount36_ay4z_core_078;
  wire popcount36_ay4z_core_079;
  wire popcount36_ay4z_core_080;
  wire popcount36_ay4z_core_082;
  wire popcount36_ay4z_core_084;
  wire popcount36_ay4z_core_085;
  wire popcount36_ay4z_core_088;
  wire popcount36_ay4z_core_089;
  wire popcount36_ay4z_core_090;
  wire popcount36_ay4z_core_092;
  wire popcount36_ay4z_core_093;
  wire popcount36_ay4z_core_094;
  wire popcount36_ay4z_core_095;
  wire popcount36_ay4z_core_096;
  wire popcount36_ay4z_core_097;
  wire popcount36_ay4z_core_098;
  wire popcount36_ay4z_core_099;
  wire popcount36_ay4z_core_100_not;
  wire popcount36_ay4z_core_101;
  wire popcount36_ay4z_core_102;
  wire popcount36_ay4z_core_103;
  wire popcount36_ay4z_core_104;
  wire popcount36_ay4z_core_106;
  wire popcount36_ay4z_core_109;
  wire popcount36_ay4z_core_113;
  wire popcount36_ay4z_core_115;
  wire popcount36_ay4z_core_116;
  wire popcount36_ay4z_core_117;
  wire popcount36_ay4z_core_119;
  wire popcount36_ay4z_core_121;
  wire popcount36_ay4z_core_123;
  wire popcount36_ay4z_core_126;
  wire popcount36_ay4z_core_127;
  wire popcount36_ay4z_core_128;
  wire popcount36_ay4z_core_129;
  wire popcount36_ay4z_core_130;
  wire popcount36_ay4z_core_133;
  wire popcount36_ay4z_core_134;
  wire popcount36_ay4z_core_135;
  wire popcount36_ay4z_core_136;
  wire popcount36_ay4z_core_137;
  wire popcount36_ay4z_core_143;
  wire popcount36_ay4z_core_144;
  wire popcount36_ay4z_core_148;
  wire popcount36_ay4z_core_151;
  wire popcount36_ay4z_core_152;
  wire popcount36_ay4z_core_154;
  wire popcount36_ay4z_core_157;
  wire popcount36_ay4z_core_158;
  wire popcount36_ay4z_core_159;
  wire popcount36_ay4z_core_160;
  wire popcount36_ay4z_core_162;
  wire popcount36_ay4z_core_163;
  wire popcount36_ay4z_core_164;
  wire popcount36_ay4z_core_165;
  wire popcount36_ay4z_core_168;
  wire popcount36_ay4z_core_169;
  wire popcount36_ay4z_core_173;
  wire popcount36_ay4z_core_175;
  wire popcount36_ay4z_core_176;
  wire popcount36_ay4z_core_177;
  wire popcount36_ay4z_core_178;
  wire popcount36_ay4z_core_179;
  wire popcount36_ay4z_core_180;
  wire popcount36_ay4z_core_181;
  wire popcount36_ay4z_core_184;
  wire popcount36_ay4z_core_185;
  wire popcount36_ay4z_core_186;
  wire popcount36_ay4z_core_188;
  wire popcount36_ay4z_core_189;
  wire popcount36_ay4z_core_190;
  wire popcount36_ay4z_core_191;
  wire popcount36_ay4z_core_195;
  wire popcount36_ay4z_core_196;
  wire popcount36_ay4z_core_197;
  wire popcount36_ay4z_core_198;
  wire popcount36_ay4z_core_201;
  wire popcount36_ay4z_core_202;
  wire popcount36_ay4z_core_204_not;
  wire popcount36_ay4z_core_206;
  wire popcount36_ay4z_core_210;
  wire popcount36_ay4z_core_211;
  wire popcount36_ay4z_core_212;
  wire popcount36_ay4z_core_214;
  wire popcount36_ay4z_core_216;
  wire popcount36_ay4z_core_217;
  wire popcount36_ay4z_core_221;
  wire popcount36_ay4z_core_222;
  wire popcount36_ay4z_core_224;
  wire popcount36_ay4z_core_226;
  wire popcount36_ay4z_core_227;
  wire popcount36_ay4z_core_228;
  wire popcount36_ay4z_core_229;
  wire popcount36_ay4z_core_230;
  wire popcount36_ay4z_core_231;
  wire popcount36_ay4z_core_232;
  wire popcount36_ay4z_core_233;
  wire popcount36_ay4z_core_234;
  wire popcount36_ay4z_core_235;
  wire popcount36_ay4z_core_236;
  wire popcount36_ay4z_core_237;
  wire popcount36_ay4z_core_238;
  wire popcount36_ay4z_core_239;
  wire popcount36_ay4z_core_240;
  wire popcount36_ay4z_core_241;
  wire popcount36_ay4z_core_243;
  wire popcount36_ay4z_core_245;
  wire popcount36_ay4z_core_246;
  wire popcount36_ay4z_core_248;
  wire popcount36_ay4z_core_249;
  wire popcount36_ay4z_core_250;
  wire popcount36_ay4z_core_252;
  wire popcount36_ay4z_core_255;
  wire popcount36_ay4z_core_257;
  wire popcount36_ay4z_core_259;
  wire popcount36_ay4z_core_260;
  wire popcount36_ay4z_core_262;
  wire popcount36_ay4z_core_264;
  wire popcount36_ay4z_core_266;
  wire popcount36_ay4z_core_267;
  wire popcount36_ay4z_core_268;
  wire popcount36_ay4z_core_270;
  wire popcount36_ay4z_core_271;
  wire popcount36_ay4z_core_272;
  wire popcount36_ay4z_core_273;
  wire popcount36_ay4z_core_274;
  wire popcount36_ay4z_core_275;

  assign popcount36_ay4z_core_039 = ~(input_a[9] ^ input_a[3]);
  assign popcount36_ay4z_core_040 = ~(input_a[21] | input_a[19]);
  assign popcount36_ay4z_core_041 = ~(input_a[16] | input_a[8]);
  assign popcount36_ay4z_core_043 = input_a[20] | input_a[30];
  assign popcount36_ay4z_core_045 = ~(input_a[16] & input_a[12]);
  assign popcount36_ay4z_core_046 = ~(input_a[31] | input_a[19]);
  assign popcount36_ay4z_core_048 = ~(input_a[32] & input_a[24]);
  assign popcount36_ay4z_core_050 = ~(input_a[25] | input_a[3]);
  assign popcount36_ay4z_core_051 = ~(input_a[9] ^ input_a[3]);
  assign popcount36_ay4z_core_052 = ~(input_a[18] | input_a[30]);
  assign popcount36_ay4z_core_054 = input_a[12] | input_a[28];
  assign popcount36_ay4z_core_059 = ~(input_a[20] ^ input_a[17]);
  assign popcount36_ay4z_core_061 = ~(input_a[29] & input_a[16]);
  assign popcount36_ay4z_core_062 = input_a[33] | input_a[32];
  assign popcount36_ay4z_core_063 = ~(input_a[6] ^ input_a[30]);
  assign popcount36_ay4z_core_064 = ~(input_a[3] & input_a[25]);
  assign popcount36_ay4z_core_065 = ~(input_a[26] & input_a[14]);
  assign popcount36_ay4z_core_068 = input_a[18] & input_a[33];
  assign popcount36_ay4z_core_069 = input_a[7] | input_a[2];
  assign popcount36_ay4z_core_073 = input_a[26] ^ input_a[30];
  assign popcount36_ay4z_core_075 = ~(input_a[23] | input_a[27]);
  assign popcount36_ay4z_core_077 = ~input_a[29];
  assign popcount36_ay4z_core_078 = input_a[31] | input_a[5];
  assign popcount36_ay4z_core_079 = ~(input_a[6] & input_a[32]);
  assign popcount36_ay4z_core_080 = ~input_a[13];
  assign popcount36_ay4z_core_082 = ~(input_a[25] | input_a[18]);
  assign popcount36_ay4z_core_084 = ~(input_a[15] | input_a[0]);
  assign popcount36_ay4z_core_085 = ~(input_a[26] & input_a[26]);
  assign popcount36_ay4z_core_088 = ~(input_a[14] ^ input_a[35]);
  assign popcount36_ay4z_core_089 = input_a[9] ^ input_a[28];
  assign popcount36_ay4z_core_090 = input_a[30] & input_a[16];
  assign popcount36_ay4z_core_092 = input_a[34] | input_a[30];
  assign popcount36_ay4z_core_093 = ~(input_a[18] ^ input_a[21]);
  assign popcount36_ay4z_core_094 = ~(input_a[19] | input_a[19]);
  assign popcount36_ay4z_core_095 = input_a[23] & input_a[19];
  assign popcount36_ay4z_core_096 = ~(input_a[26] & input_a[8]);
  assign popcount36_ay4z_core_097 = ~(input_a[8] ^ input_a[9]);
  assign popcount36_ay4z_core_098 = ~(input_a[11] & input_a[12]);
  assign popcount36_ay4z_core_099 = input_a[29] ^ input_a[18];
  assign popcount36_ay4z_core_100_not = ~input_a[4];
  assign popcount36_ay4z_core_101 = input_a[12] | input_a[29];
  assign popcount36_ay4z_core_102 = input_a[19] & input_a[31];
  assign popcount36_ay4z_core_103 = ~(input_a[7] | input_a[26]);
  assign popcount36_ay4z_core_104 = ~input_a[17];
  assign popcount36_ay4z_core_106 = ~(input_a[12] | input_a[16]);
  assign popcount36_ay4z_core_109 = ~input_a[21];
  assign popcount36_ay4z_core_113 = ~(input_a[31] | input_a[17]);
  assign popcount36_ay4z_core_115 = input_a[23] & input_a[11];
  assign popcount36_ay4z_core_116 = input_a[34] ^ input_a[30];
  assign popcount36_ay4z_core_117 = input_a[5] | input_a[34];
  assign popcount36_ay4z_core_119 = input_a[4] | input_a[18];
  assign popcount36_ay4z_core_121 = input_a[7] ^ input_a[35];
  assign popcount36_ay4z_core_123 = ~input_a[32];
  assign popcount36_ay4z_core_126 = ~(input_a[5] | input_a[15]);
  assign popcount36_ay4z_core_127 = ~(input_a[25] & input_a[1]);
  assign popcount36_ay4z_core_128 = ~(input_a[8] & input_a[10]);
  assign popcount36_ay4z_core_129 = input_a[16] & input_a[13];
  assign popcount36_ay4z_core_130 = input_a[14] | input_a[2];
  assign popcount36_ay4z_core_133 = ~(input_a[6] & input_a[29]);
  assign popcount36_ay4z_core_134 = input_a[20] | input_a[29];
  assign popcount36_ay4z_core_135 = ~(input_a[26] ^ input_a[19]);
  assign popcount36_ay4z_core_136 = ~(input_a[15] & input_a[29]);
  assign popcount36_ay4z_core_137 = ~(input_a[20] & input_a[29]);
  assign popcount36_ay4z_core_143 = input_a[16] | input_a[32];
  assign popcount36_ay4z_core_144 = input_a[23] ^ input_a[22];
  assign popcount36_ay4z_core_148 = ~(input_a[28] ^ input_a[13]);
  assign popcount36_ay4z_core_151 = input_a[29] ^ input_a[24];
  assign popcount36_ay4z_core_152 = input_a[26] ^ input_a[17];
  assign popcount36_ay4z_core_154 = ~input_a[28];
  assign popcount36_ay4z_core_157 = input_a[22] & input_a[1];
  assign popcount36_ay4z_core_158 = ~(input_a[30] | input_a[22]);
  assign popcount36_ay4z_core_159 = ~(input_a[15] | input_a[8]);
  assign popcount36_ay4z_core_160 = ~input_a[4];
  assign popcount36_ay4z_core_162 = ~(input_a[0] & input_a[24]);
  assign popcount36_ay4z_core_163 = input_a[31] | input_a[35];
  assign popcount36_ay4z_core_164 = ~(input_a[3] ^ input_a[31]);
  assign popcount36_ay4z_core_165 = input_a[18] & input_a[33];
  assign popcount36_ay4z_core_168 = ~(input_a[11] & input_a[7]);
  assign popcount36_ay4z_core_169 = ~input_a[17];
  assign popcount36_ay4z_core_173 = input_a[34] & input_a[29];
  assign popcount36_ay4z_core_175 = input_a[30] | input_a[32];
  assign popcount36_ay4z_core_176 = ~(input_a[34] | input_a[29]);
  assign popcount36_ay4z_core_177 = input_a[21] | input_a[23];
  assign popcount36_ay4z_core_178 = ~input_a[32];
  assign popcount36_ay4z_core_179 = input_a[19] ^ input_a[24];
  assign popcount36_ay4z_core_180 = ~(input_a[17] | input_a[19]);
  assign popcount36_ay4z_core_181 = input_a[8] | input_a[25];
  assign popcount36_ay4z_core_184 = input_a[11] & input_a[3];
  assign popcount36_ay4z_core_185 = ~input_a[0];
  assign popcount36_ay4z_core_186 = ~(input_a[23] ^ input_a[28]);
  assign popcount36_ay4z_core_188 = ~(input_a[28] | input_a[14]);
  assign popcount36_ay4z_core_189 = input_a[10] | input_a[13];
  assign popcount36_ay4z_core_190 = ~(input_a[24] | input_a[31]);
  assign popcount36_ay4z_core_191 = ~(input_a[6] | input_a[14]);
  assign popcount36_ay4z_core_195 = ~input_a[21];
  assign popcount36_ay4z_core_196 = ~input_a[33];
  assign popcount36_ay4z_core_197 = input_a[9] & input_a[33];
  assign popcount36_ay4z_core_198 = input_a[5] & input_a[23];
  assign popcount36_ay4z_core_201 = input_a[13] ^ input_a[18];
  assign popcount36_ay4z_core_202 = input_a[1] | input_a[35];
  assign popcount36_ay4z_core_204_not = ~input_a[24];
  assign popcount36_ay4z_core_206 = input_a[35] | input_a[21];
  assign popcount36_ay4z_core_210 = input_a[6] & input_a[18];
  assign popcount36_ay4z_core_211 = input_a[26] | input_a[21];
  assign popcount36_ay4z_core_212 = ~(input_a[13] ^ input_a[32]);
  assign popcount36_ay4z_core_214 = ~(input_a[8] | input_a[29]);
  assign popcount36_ay4z_core_216 = ~input_a[8];
  assign popcount36_ay4z_core_217 = ~(input_a[2] | input_a[13]);
  assign popcount36_ay4z_core_221 = input_a[22] | input_a[12];
  assign popcount36_ay4z_core_222 = input_a[25] & input_a[21];
  assign popcount36_ay4z_core_224 = ~(input_a[10] & input_a[29]);
  assign popcount36_ay4z_core_226 = ~(input_a[27] ^ input_a[30]);
  assign popcount36_ay4z_core_227 = input_a[5] | input_a[6];
  assign popcount36_ay4z_core_228 = input_a[23] & input_a[7];
  assign popcount36_ay4z_core_229 = input_a[4] & input_a[34];
  assign popcount36_ay4z_core_230 = ~(input_a[33] | input_a[7]);
  assign popcount36_ay4z_core_231 = input_a[14] | input_a[23];
  assign popcount36_ay4z_core_232 = ~(input_a[8] ^ input_a[0]);
  assign popcount36_ay4z_core_233 = ~(input_a[7] & input_a[21]);
  assign popcount36_ay4z_core_234 = ~input_a[11];
  assign popcount36_ay4z_core_235 = ~(input_a[11] ^ input_a[10]);
  assign popcount36_ay4z_core_236 = ~(input_a[16] ^ input_a[14]);
  assign popcount36_ay4z_core_237 = input_a[21] | input_a[25];
  assign popcount36_ay4z_core_238 = ~(input_a[26] | input_a[21]);
  assign popcount36_ay4z_core_239 = input_a[0] & input_a[2];
  assign popcount36_ay4z_core_240 = ~(input_a[6] & input_a[20]);
  assign popcount36_ay4z_core_241 = ~(input_a[12] ^ input_a[24]);
  assign popcount36_ay4z_core_243 = input_a[9] | input_a[18];
  assign popcount36_ay4z_core_245 = input_a[29] & input_a[27];
  assign popcount36_ay4z_core_246 = input_a[17] | input_a[4];
  assign popcount36_ay4z_core_248 = ~input_a[18];
  assign popcount36_ay4z_core_249 = input_a[24] & input_a[1];
  assign popcount36_ay4z_core_250 = ~(input_a[22] ^ input_a[33]);
  assign popcount36_ay4z_core_252 = ~input_a[2];
  assign popcount36_ay4z_core_255 = ~input_a[27];
  assign popcount36_ay4z_core_257 = input_a[11] | input_a[32];
  assign popcount36_ay4z_core_259 = ~(input_a[35] & input_a[2]);
  assign popcount36_ay4z_core_260 = ~(input_a[31] | input_a[31]);
  assign popcount36_ay4z_core_262 = ~(input_a[11] | input_a[28]);
  assign popcount36_ay4z_core_264 = input_a[1] & input_a[20];
  assign popcount36_ay4z_core_266 = ~(input_a[1] ^ input_a[17]);
  assign popcount36_ay4z_core_267 = ~(input_a[31] ^ input_a[13]);
  assign popcount36_ay4z_core_268 = ~(input_a[17] | input_a[20]);
  assign popcount36_ay4z_core_270 = ~(input_a[11] & input_a[18]);
  assign popcount36_ay4z_core_271 = ~input_a[15];
  assign popcount36_ay4z_core_272 = ~(input_a[8] | input_a[27]);
  assign popcount36_ay4z_core_273 = ~(input_a[11] | input_a[7]);
  assign popcount36_ay4z_core_274 = ~(input_a[17] | input_a[1]);
  assign popcount36_ay4z_core_275 = input_a[11] & input_a[20];

  assign popcount36_ay4z_out[0] = input_a[5];
  assign popcount36_ay4z_out[1] = 1'b1;
  assign popcount36_ay4z_out[2] = 1'b0;
  assign popcount36_ay4z_out[3] = 1'b0;
  assign popcount36_ay4z_out[4] = 1'b1;
  assign popcount36_ay4z_out[5] = 1'b0;
endmodule