// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.49838
// WCE=13.0
// EP=0.792877%
// Printed PDK parameters:
//  Area=55410982.0
//  Delay=68461520.0
//  Power=3002500.0

module popcount30_wgv4(input [29:0] input_a, output [4:0] popcount30_wgv4_out);
  wire popcount30_wgv4_core_032;
  wire popcount30_wgv4_core_033;
  wire popcount30_wgv4_core_035;
  wire popcount30_wgv4_core_036;
  wire popcount30_wgv4_core_038;
  wire popcount30_wgv4_core_039;
  wire popcount30_wgv4_core_042;
  wire popcount30_wgv4_core_044;
  wire popcount30_wgv4_core_045;
  wire popcount30_wgv4_core_046;
  wire popcount30_wgv4_core_047;
  wire popcount30_wgv4_core_049;
  wire popcount30_wgv4_core_050;
  wire popcount30_wgv4_core_051;
  wire popcount30_wgv4_core_052;
  wire popcount30_wgv4_core_053;
  wire popcount30_wgv4_core_054;
  wire popcount30_wgv4_core_055;
  wire popcount30_wgv4_core_057;
  wire popcount30_wgv4_core_058;
  wire popcount30_wgv4_core_059;
  wire popcount30_wgv4_core_061;
  wire popcount30_wgv4_core_062;
  wire popcount30_wgv4_core_064;
  wire popcount30_wgv4_core_065;
  wire popcount30_wgv4_core_066_not;
  wire popcount30_wgv4_core_067;
  wire popcount30_wgv4_core_068;
  wire popcount30_wgv4_core_070;
  wire popcount30_wgv4_core_073;
  wire popcount30_wgv4_core_077;
  wire popcount30_wgv4_core_078;
  wire popcount30_wgv4_core_080;
  wire popcount30_wgv4_core_081;
  wire popcount30_wgv4_core_082;
  wire popcount30_wgv4_core_084;
  wire popcount30_wgv4_core_085;
  wire popcount30_wgv4_core_087;
  wire popcount30_wgv4_core_093;
  wire popcount30_wgv4_core_094;
  wire popcount30_wgv4_core_096;
  wire popcount30_wgv4_core_097;
  wire popcount30_wgv4_core_098;
  wire popcount30_wgv4_core_102;
  wire popcount30_wgv4_core_103;
  wire popcount30_wgv4_core_104;
  wire popcount30_wgv4_core_105;
  wire popcount30_wgv4_core_106;
  wire popcount30_wgv4_core_108;
  wire popcount30_wgv4_core_111;
  wire popcount30_wgv4_core_115;
  wire popcount30_wgv4_core_116;
  wire popcount30_wgv4_core_118;
  wire popcount30_wgv4_core_119;
  wire popcount30_wgv4_core_120;
  wire popcount30_wgv4_core_121;
  wire popcount30_wgv4_core_122;
  wire popcount30_wgv4_core_123;
  wire popcount30_wgv4_core_124;
  wire popcount30_wgv4_core_126;
  wire popcount30_wgv4_core_131;
  wire popcount30_wgv4_core_132;
  wire popcount30_wgv4_core_133;
  wire popcount30_wgv4_core_134;
  wire popcount30_wgv4_core_135;
  wire popcount30_wgv4_core_138;
  wire popcount30_wgv4_core_141;
  wire popcount30_wgv4_core_142;
  wire popcount30_wgv4_core_143;
  wire popcount30_wgv4_core_144;
  wire popcount30_wgv4_core_145;
  wire popcount30_wgv4_core_146;
  wire popcount30_wgv4_core_147;
  wire popcount30_wgv4_core_148;
  wire popcount30_wgv4_core_149;
  wire popcount30_wgv4_core_150;
  wire popcount30_wgv4_core_152;
  wire popcount30_wgv4_core_153;
  wire popcount30_wgv4_core_154;
  wire popcount30_wgv4_core_155;
  wire popcount30_wgv4_core_156;
  wire popcount30_wgv4_core_157;
  wire popcount30_wgv4_core_158;
  wire popcount30_wgv4_core_159;
  wire popcount30_wgv4_core_160;
  wire popcount30_wgv4_core_161;
  wire popcount30_wgv4_core_163;
  wire popcount30_wgv4_core_164;
  wire popcount30_wgv4_core_165;
  wire popcount30_wgv4_core_166;
  wire popcount30_wgv4_core_167;
  wire popcount30_wgv4_core_168;
  wire popcount30_wgv4_core_169;
  wire popcount30_wgv4_core_170;
  wire popcount30_wgv4_core_171;
  wire popcount30_wgv4_core_172;
  wire popcount30_wgv4_core_175;
  wire popcount30_wgv4_core_176;
  wire popcount30_wgv4_core_177;
  wire popcount30_wgv4_core_178;
  wire popcount30_wgv4_core_182;
  wire popcount30_wgv4_core_183;
  wire popcount30_wgv4_core_184;
  wire popcount30_wgv4_core_185;
  wire popcount30_wgv4_core_186;
  wire popcount30_wgv4_core_188;
  wire popcount30_wgv4_core_190;
  wire popcount30_wgv4_core_192;
  wire popcount30_wgv4_core_193;
  wire popcount30_wgv4_core_195;
  wire popcount30_wgv4_core_199;
  wire popcount30_wgv4_core_200;
  wire popcount30_wgv4_core_201;
  wire popcount30_wgv4_core_202;
  wire popcount30_wgv4_core_203;
  wire popcount30_wgv4_core_204;
  wire popcount30_wgv4_core_205;
  wire popcount30_wgv4_core_206;
  wire popcount30_wgv4_core_207;
  wire popcount30_wgv4_core_208;
  wire popcount30_wgv4_core_210;
  wire popcount30_wgv4_core_211;

  assign popcount30_wgv4_core_032 = input_a[16] | input_a[15];
  assign popcount30_wgv4_core_033 = input_a[14] & input_a[10];
  assign popcount30_wgv4_core_035 = input_a[11] & popcount30_wgv4_core_032;
  assign popcount30_wgv4_core_036 = popcount30_wgv4_core_033 | popcount30_wgv4_core_035;
  assign popcount30_wgv4_core_038 = input_a[3] ^ input_a[5];
  assign popcount30_wgv4_core_039 = input_a[3] & input_a[4];
  assign popcount30_wgv4_core_042 = ~(input_a[3] | input_a[23]);
  assign popcount30_wgv4_core_044 = input_a[4] ^ input_a[5];
  assign popcount30_wgv4_core_045 = popcount30_wgv4_core_039 & input_a[5];
  assign popcount30_wgv4_core_046 = popcount30_wgv4_core_044 | popcount30_wgv4_core_038;
  assign popcount30_wgv4_core_047 = ~(input_a[8] ^ input_a[5]);
  assign popcount30_wgv4_core_049 = input_a[14] & input_a[4];
  assign popcount30_wgv4_core_050 = input_a[0] & input_a[8];
  assign popcount30_wgv4_core_051 = popcount30_wgv4_core_036 ^ popcount30_wgv4_core_046;
  assign popcount30_wgv4_core_052 = popcount30_wgv4_core_036 & popcount30_wgv4_core_046;
  assign popcount30_wgv4_core_053 = popcount30_wgv4_core_051 ^ popcount30_wgv4_core_050;
  assign popcount30_wgv4_core_054 = popcount30_wgv4_core_051 & popcount30_wgv4_core_050;
  assign popcount30_wgv4_core_055 = popcount30_wgv4_core_052 | popcount30_wgv4_core_054;
  assign popcount30_wgv4_core_057 = ~(input_a[13] ^ input_a[29]);
  assign popcount30_wgv4_core_058 = popcount30_wgv4_core_045 | popcount30_wgv4_core_055;
  assign popcount30_wgv4_core_059 = input_a[28] | input_a[20];
  assign popcount30_wgv4_core_061 = ~(input_a[27] ^ input_a[29]);
  assign popcount30_wgv4_core_062 = input_a[12] & input_a[16];
  assign popcount30_wgv4_core_064 = input_a[2] & input_a[9];
  assign popcount30_wgv4_core_065 = ~(input_a[25] ^ input_a[2]);
  assign popcount30_wgv4_core_066_not = ~input_a[13];
  assign popcount30_wgv4_core_067 = popcount30_wgv4_core_062 | popcount30_wgv4_core_064;
  assign popcount30_wgv4_core_068 = input_a[0] | input_a[3];
  assign popcount30_wgv4_core_070 = input_a[20] & input_a[27];
  assign popcount30_wgv4_core_073 = ~(input_a[18] & input_a[1]);
  assign popcount30_wgv4_core_077 = ~(input_a[10] & input_a[10]);
  assign popcount30_wgv4_core_078 = ~input_a[2];
  assign popcount30_wgv4_core_080 = input_a[7] & input_a[6];
  assign popcount30_wgv4_core_081 = ~(input_a[3] | input_a[24]);
  assign popcount30_wgv4_core_082 = ~(input_a[13] | input_a[29]);
  assign popcount30_wgv4_core_084 = input_a[28] & input_a[15];
  assign popcount30_wgv4_core_085 = popcount30_wgv4_core_067 | popcount30_wgv4_core_080;
  assign popcount30_wgv4_core_087 = ~popcount30_wgv4_core_085;
  assign popcount30_wgv4_core_093 = input_a[22] ^ input_a[9];
  assign popcount30_wgv4_core_094 = ~(input_a[19] | input_a[11]);
  assign popcount30_wgv4_core_096 = ~(input_a[11] & input_a[17]);
  assign popcount30_wgv4_core_097 = popcount30_wgv4_core_053 ^ popcount30_wgv4_core_087;
  assign popcount30_wgv4_core_098 = popcount30_wgv4_core_053 & popcount30_wgv4_core_087;
  assign popcount30_wgv4_core_102 = popcount30_wgv4_core_058 ^ popcount30_wgv4_core_085;
  assign popcount30_wgv4_core_103 = popcount30_wgv4_core_058 & popcount30_wgv4_core_085;
  assign popcount30_wgv4_core_104 = popcount30_wgv4_core_102 ^ popcount30_wgv4_core_098;
  assign popcount30_wgv4_core_105 = popcount30_wgv4_core_102 & popcount30_wgv4_core_098;
  assign popcount30_wgv4_core_106 = popcount30_wgv4_core_103 | popcount30_wgv4_core_105;
  assign popcount30_wgv4_core_108 = input_a[27] ^ input_a[0];
  assign popcount30_wgv4_core_111 = input_a[19] & input_a[29];
  assign popcount30_wgv4_core_115 = ~(input_a[10] | input_a[17]);
  assign popcount30_wgv4_core_116 = input_a[17] | input_a[1];
  assign popcount30_wgv4_core_118 = input_a[18] ^ input_a[19];
  assign popcount30_wgv4_core_119 = input_a[18] & input_a[19];
  assign popcount30_wgv4_core_120 = input_a[20] ^ input_a[21];
  assign popcount30_wgv4_core_121 = input_a[20] & input_a[21];
  assign popcount30_wgv4_core_122 = popcount30_wgv4_core_118 ^ popcount30_wgv4_core_120;
  assign popcount30_wgv4_core_123 = popcount30_wgv4_core_118 & popcount30_wgv4_core_120;
  assign popcount30_wgv4_core_124 = popcount30_wgv4_core_119 ^ popcount30_wgv4_core_121;
  assign popcount30_wgv4_core_126 = popcount30_wgv4_core_124 | popcount30_wgv4_core_123;
  assign popcount30_wgv4_core_131 = popcount30_wgv4_core_116 ^ popcount30_wgv4_core_126;
  assign popcount30_wgv4_core_132 = popcount30_wgv4_core_116 & popcount30_wgv4_core_126;
  assign popcount30_wgv4_core_133 = popcount30_wgv4_core_131 ^ popcount30_wgv4_core_122;
  assign popcount30_wgv4_core_134 = popcount30_wgv4_core_131 & popcount30_wgv4_core_122;
  assign popcount30_wgv4_core_135 = popcount30_wgv4_core_132 | popcount30_wgv4_core_134;
  assign popcount30_wgv4_core_138 = popcount30_wgv4_core_119 | popcount30_wgv4_core_135;
  assign popcount30_wgv4_core_141 = input_a[22] ^ input_a[23];
  assign popcount30_wgv4_core_142 = input_a[22] & input_a[23];
  assign popcount30_wgv4_core_143 = input_a[24] ^ input_a[25];
  assign popcount30_wgv4_core_144 = input_a[24] & input_a[25];
  assign popcount30_wgv4_core_145 = popcount30_wgv4_core_141 ^ popcount30_wgv4_core_143;
  assign popcount30_wgv4_core_146 = popcount30_wgv4_core_141 & popcount30_wgv4_core_143;
  assign popcount30_wgv4_core_147 = popcount30_wgv4_core_142 ^ popcount30_wgv4_core_144;
  assign popcount30_wgv4_core_148 = input_a[23] & popcount30_wgv4_core_144;
  assign popcount30_wgv4_core_149 = popcount30_wgv4_core_147 | popcount30_wgv4_core_146;
  assign popcount30_wgv4_core_150 = input_a[12] & input_a[13];
  assign popcount30_wgv4_core_152 = input_a[26] ^ input_a[27];
  assign popcount30_wgv4_core_153 = input_a[26] & input_a[27];
  assign popcount30_wgv4_core_154 = input_a[28] ^ input_a[29];
  assign popcount30_wgv4_core_155 = input_a[28] & input_a[29];
  assign popcount30_wgv4_core_156 = popcount30_wgv4_core_152 ^ popcount30_wgv4_core_154;
  assign popcount30_wgv4_core_157 = popcount30_wgv4_core_152 & popcount30_wgv4_core_154;
  assign popcount30_wgv4_core_158 = popcount30_wgv4_core_153 ^ popcount30_wgv4_core_155;
  assign popcount30_wgv4_core_159 = popcount30_wgv4_core_153 & input_a[29];
  assign popcount30_wgv4_core_160 = popcount30_wgv4_core_158 | popcount30_wgv4_core_157;
  assign popcount30_wgv4_core_161 = input_a[25] | input_a[11];
  assign popcount30_wgv4_core_163 = ~input_a[23];
  assign popcount30_wgv4_core_164 = popcount30_wgv4_core_145 & popcount30_wgv4_core_156;
  assign popcount30_wgv4_core_165 = popcount30_wgv4_core_149 ^ popcount30_wgv4_core_160;
  assign popcount30_wgv4_core_166 = popcount30_wgv4_core_149 & popcount30_wgv4_core_160;
  assign popcount30_wgv4_core_167 = popcount30_wgv4_core_165 ^ popcount30_wgv4_core_164;
  assign popcount30_wgv4_core_168 = popcount30_wgv4_core_165 & popcount30_wgv4_core_164;
  assign popcount30_wgv4_core_169 = popcount30_wgv4_core_166 | popcount30_wgv4_core_168;
  assign popcount30_wgv4_core_170 = popcount30_wgv4_core_148 | popcount30_wgv4_core_159;
  assign popcount30_wgv4_core_171 = ~(input_a[19] ^ input_a[9]);
  assign popcount30_wgv4_core_172 = popcount30_wgv4_core_170 | popcount30_wgv4_core_169;
  assign popcount30_wgv4_core_175 = ~(input_a[14] ^ input_a[5]);
  assign popcount30_wgv4_core_176 = input_a[17] & input_a[4];
  assign popcount30_wgv4_core_177 = popcount30_wgv4_core_133 ^ popcount30_wgv4_core_167;
  assign popcount30_wgv4_core_178 = popcount30_wgv4_core_133 & popcount30_wgv4_core_167;
  assign popcount30_wgv4_core_182 = popcount30_wgv4_core_138 ^ popcount30_wgv4_core_172;
  assign popcount30_wgv4_core_183 = popcount30_wgv4_core_138 & popcount30_wgv4_core_172;
  assign popcount30_wgv4_core_184 = popcount30_wgv4_core_182 ^ popcount30_wgv4_core_178;
  assign popcount30_wgv4_core_185 = popcount30_wgv4_core_182 & popcount30_wgv4_core_178;
  assign popcount30_wgv4_core_186 = popcount30_wgv4_core_183 | popcount30_wgv4_core_185;
  assign popcount30_wgv4_core_188 = ~(input_a[29] ^ input_a[4]);
  assign popcount30_wgv4_core_190 = ~(input_a[6] & input_a[2]);
  assign popcount30_wgv4_core_192 = ~(input_a[13] | input_a[24]);
  assign popcount30_wgv4_core_193 = ~input_a[14];
  assign popcount30_wgv4_core_195 = popcount30_wgv4_core_097 & popcount30_wgv4_core_177;
  assign popcount30_wgv4_core_199 = popcount30_wgv4_core_104 ^ popcount30_wgv4_core_184;
  assign popcount30_wgv4_core_200 = popcount30_wgv4_core_104 & popcount30_wgv4_core_184;
  assign popcount30_wgv4_core_201 = popcount30_wgv4_core_199 ^ popcount30_wgv4_core_195;
  assign popcount30_wgv4_core_202 = popcount30_wgv4_core_199 & popcount30_wgv4_core_195;
  assign popcount30_wgv4_core_203 = popcount30_wgv4_core_200 | popcount30_wgv4_core_202;
  assign popcount30_wgv4_core_204 = popcount30_wgv4_core_106 ^ popcount30_wgv4_core_186;
  assign popcount30_wgv4_core_205 = popcount30_wgv4_core_106 & popcount30_wgv4_core_186;
  assign popcount30_wgv4_core_206 = popcount30_wgv4_core_204 ^ popcount30_wgv4_core_203;
  assign popcount30_wgv4_core_207 = popcount30_wgv4_core_204 & popcount30_wgv4_core_203;
  assign popcount30_wgv4_core_208 = popcount30_wgv4_core_205 | popcount30_wgv4_core_207;
  assign popcount30_wgv4_core_210 = input_a[1] ^ input_a[13];
  assign popcount30_wgv4_core_211 = ~(input_a[21] | input_a[28]);

  assign popcount30_wgv4_out[0] = popcount30_wgv4_core_206;
  assign popcount30_wgv4_out[1] = input_a[13];
  assign popcount30_wgv4_out[2] = popcount30_wgv4_core_201;
  assign popcount30_wgv4_out[3] = popcount30_wgv4_core_206;
  assign popcount30_wgv4_out[4] = popcount30_wgv4_core_208;
endmodule