// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.40858
// WCE=33.0
// EP=0.944491%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_ugbo(input [35:0] input_a, output [5:0] popcount36_ugbo_out);
  wire popcount36_ugbo_core_038;
  wire popcount36_ugbo_core_039;
  wire popcount36_ugbo_core_040;
  wire popcount36_ugbo_core_041;
  wire popcount36_ugbo_core_042;
  wire popcount36_ugbo_core_044;
  wire popcount36_ugbo_core_045;
  wire popcount36_ugbo_core_048;
  wire popcount36_ugbo_core_049;
  wire popcount36_ugbo_core_052;
  wire popcount36_ugbo_core_053;
  wire popcount36_ugbo_core_054;
  wire popcount36_ugbo_core_056;
  wire popcount36_ugbo_core_057;
  wire popcount36_ugbo_core_058;
  wire popcount36_ugbo_core_060;
  wire popcount36_ugbo_core_062;
  wire popcount36_ugbo_core_063;
  wire popcount36_ugbo_core_064;
  wire popcount36_ugbo_core_065;
  wire popcount36_ugbo_core_066;
  wire popcount36_ugbo_core_067;
  wire popcount36_ugbo_core_069;
  wire popcount36_ugbo_core_070;
  wire popcount36_ugbo_core_071;
  wire popcount36_ugbo_core_072;
  wire popcount36_ugbo_core_073;
  wire popcount36_ugbo_core_074;
  wire popcount36_ugbo_core_075;
  wire popcount36_ugbo_core_077;
  wire popcount36_ugbo_core_078;
  wire popcount36_ugbo_core_082;
  wire popcount36_ugbo_core_083;
  wire popcount36_ugbo_core_084;
  wire popcount36_ugbo_core_087;
  wire popcount36_ugbo_core_088;
  wire popcount36_ugbo_core_090;
  wire popcount36_ugbo_core_091;
  wire popcount36_ugbo_core_092;
  wire popcount36_ugbo_core_093;
  wire popcount36_ugbo_core_095;
  wire popcount36_ugbo_core_096;
  wire popcount36_ugbo_core_097;
  wire popcount36_ugbo_core_098;
  wire popcount36_ugbo_core_100;
  wire popcount36_ugbo_core_101;
  wire popcount36_ugbo_core_102;
  wire popcount36_ugbo_core_104;
  wire popcount36_ugbo_core_105;
  wire popcount36_ugbo_core_108;
  wire popcount36_ugbo_core_109;
  wire popcount36_ugbo_core_111;
  wire popcount36_ugbo_core_112;
  wire popcount36_ugbo_core_113;
  wire popcount36_ugbo_core_115;
  wire popcount36_ugbo_core_116;
  wire popcount36_ugbo_core_117;
  wire popcount36_ugbo_core_118;
  wire popcount36_ugbo_core_120;
  wire popcount36_ugbo_core_121;
  wire popcount36_ugbo_core_122;
  wire popcount36_ugbo_core_123;
  wire popcount36_ugbo_core_124;
  wire popcount36_ugbo_core_125;
  wire popcount36_ugbo_core_126;
  wire popcount36_ugbo_core_127;
  wire popcount36_ugbo_core_128;
  wire popcount36_ugbo_core_131;
  wire popcount36_ugbo_core_132;
  wire popcount36_ugbo_core_133;
  wire popcount36_ugbo_core_134;
  wire popcount36_ugbo_core_136;
  wire popcount36_ugbo_core_137;
  wire popcount36_ugbo_core_138;
  wire popcount36_ugbo_core_140;
  wire popcount36_ugbo_core_141;
  wire popcount36_ugbo_core_143;
  wire popcount36_ugbo_core_145;
  wire popcount36_ugbo_core_146;
  wire popcount36_ugbo_core_148;
  wire popcount36_ugbo_core_149;
  wire popcount36_ugbo_core_151;
  wire popcount36_ugbo_core_152;
  wire popcount36_ugbo_core_153;
  wire popcount36_ugbo_core_154_not;
  wire popcount36_ugbo_core_155;
  wire popcount36_ugbo_core_156;
  wire popcount36_ugbo_core_157;
  wire popcount36_ugbo_core_160;
  wire popcount36_ugbo_core_161;
  wire popcount36_ugbo_core_166;
  wire popcount36_ugbo_core_168;
  wire popcount36_ugbo_core_169;
  wire popcount36_ugbo_core_171;
  wire popcount36_ugbo_core_172;
  wire popcount36_ugbo_core_173;
  wire popcount36_ugbo_core_174;
  wire popcount36_ugbo_core_175;
  wire popcount36_ugbo_core_177;
  wire popcount36_ugbo_core_180;
  wire popcount36_ugbo_core_181;
  wire popcount36_ugbo_core_183;
  wire popcount36_ugbo_core_184;
  wire popcount36_ugbo_core_185;
  wire popcount36_ugbo_core_186;
  wire popcount36_ugbo_core_187_not;
  wire popcount36_ugbo_core_188;
  wire popcount36_ugbo_core_189;
  wire popcount36_ugbo_core_191;
  wire popcount36_ugbo_core_192;
  wire popcount36_ugbo_core_193;
  wire popcount36_ugbo_core_194;
  wire popcount36_ugbo_core_195;
  wire popcount36_ugbo_core_196;
  wire popcount36_ugbo_core_197;
  wire popcount36_ugbo_core_198;
  wire popcount36_ugbo_core_199;
  wire popcount36_ugbo_core_203;
  wire popcount36_ugbo_core_204;
  wire popcount36_ugbo_core_205;
  wire popcount36_ugbo_core_206_not;
  wire popcount36_ugbo_core_207;
  wire popcount36_ugbo_core_210;
  wire popcount36_ugbo_core_211;
  wire popcount36_ugbo_core_213_not;
  wire popcount36_ugbo_core_215;
  wire popcount36_ugbo_core_216;
  wire popcount36_ugbo_core_217;
  wire popcount36_ugbo_core_223;
  wire popcount36_ugbo_core_224;
  wire popcount36_ugbo_core_227;
  wire popcount36_ugbo_core_229;
  wire popcount36_ugbo_core_231;
  wire popcount36_ugbo_core_232;
  wire popcount36_ugbo_core_233;
  wire popcount36_ugbo_core_236;
  wire popcount36_ugbo_core_237;
  wire popcount36_ugbo_core_238;
  wire popcount36_ugbo_core_240_not;
  wire popcount36_ugbo_core_243;
  wire popcount36_ugbo_core_245;
  wire popcount36_ugbo_core_247;
  wire popcount36_ugbo_core_248;
  wire popcount36_ugbo_core_250;
  wire popcount36_ugbo_core_251_not;
  wire popcount36_ugbo_core_252;
  wire popcount36_ugbo_core_255;
  wire popcount36_ugbo_core_256;
  wire popcount36_ugbo_core_257;
  wire popcount36_ugbo_core_261;
  wire popcount36_ugbo_core_262;
  wire popcount36_ugbo_core_263;
  wire popcount36_ugbo_core_265;
  wire popcount36_ugbo_core_266;
  wire popcount36_ugbo_core_267;
  wire popcount36_ugbo_core_268;
  wire popcount36_ugbo_core_269;
  wire popcount36_ugbo_core_271;
  wire popcount36_ugbo_core_273;
  wire popcount36_ugbo_core_274;
  wire popcount36_ugbo_core_276_not;

  assign popcount36_ugbo_core_038 = ~input_a[22];
  assign popcount36_ugbo_core_039 = ~(input_a[6] ^ input_a[35]);
  assign popcount36_ugbo_core_040 = ~(input_a[3] ^ input_a[34]);
  assign popcount36_ugbo_core_041 = input_a[4] | input_a[22];
  assign popcount36_ugbo_core_042 = input_a[16] | input_a[5];
  assign popcount36_ugbo_core_044 = ~(input_a[15] ^ input_a[6]);
  assign popcount36_ugbo_core_045 = ~input_a[7];
  assign popcount36_ugbo_core_048 = ~(input_a[17] ^ input_a[12]);
  assign popcount36_ugbo_core_049 = input_a[22] ^ input_a[6];
  assign popcount36_ugbo_core_052 = ~(input_a[3] & input_a[8]);
  assign popcount36_ugbo_core_053 = ~(input_a[0] ^ input_a[24]);
  assign popcount36_ugbo_core_054 = input_a[18] | input_a[33];
  assign popcount36_ugbo_core_056 = ~input_a[26];
  assign popcount36_ugbo_core_057 = ~input_a[6];
  assign popcount36_ugbo_core_058 = input_a[30] ^ input_a[30];
  assign popcount36_ugbo_core_060 = ~input_a[9];
  assign popcount36_ugbo_core_062 = input_a[11] ^ input_a[32];
  assign popcount36_ugbo_core_063 = ~(input_a[35] ^ input_a[6]);
  assign popcount36_ugbo_core_064 = ~(input_a[18] | input_a[14]);
  assign popcount36_ugbo_core_065 = input_a[14] ^ input_a[35];
  assign popcount36_ugbo_core_066 = input_a[0] ^ input_a[23];
  assign popcount36_ugbo_core_067 = ~(input_a[14] ^ input_a[6]);
  assign popcount36_ugbo_core_069 = ~input_a[21];
  assign popcount36_ugbo_core_070 = ~(input_a[7] ^ input_a[0]);
  assign popcount36_ugbo_core_071 = input_a[25] ^ input_a[7];
  assign popcount36_ugbo_core_072 = ~(input_a[18] | input_a[9]);
  assign popcount36_ugbo_core_073 = ~(input_a[34] ^ input_a[7]);
  assign popcount36_ugbo_core_074 = input_a[10] ^ input_a[26];
  assign popcount36_ugbo_core_075 = input_a[7] ^ input_a[28];
  assign popcount36_ugbo_core_077 = ~(input_a[17] ^ input_a[20]);
  assign popcount36_ugbo_core_078 = ~input_a[21];
  assign popcount36_ugbo_core_082 = input_a[2] ^ input_a[4];
  assign popcount36_ugbo_core_083 = input_a[6] ^ input_a[30];
  assign popcount36_ugbo_core_084 = ~(input_a[34] & input_a[12]);
  assign popcount36_ugbo_core_087 = input_a[22] | input_a[3];
  assign popcount36_ugbo_core_088 = input_a[12] | input_a[32];
  assign popcount36_ugbo_core_090 = input_a[3] | input_a[17];
  assign popcount36_ugbo_core_091 = ~(input_a[11] ^ input_a[14]);
  assign popcount36_ugbo_core_092 = ~(input_a[33] ^ input_a[28]);
  assign popcount36_ugbo_core_093 = ~(input_a[23] & input_a[11]);
  assign popcount36_ugbo_core_095 = input_a[22] | input_a[2];
  assign popcount36_ugbo_core_096 = input_a[6] & input_a[27];
  assign popcount36_ugbo_core_097 = input_a[28] ^ input_a[35];
  assign popcount36_ugbo_core_098 = ~(input_a[35] & input_a[33]);
  assign popcount36_ugbo_core_100 = ~(input_a[18] ^ input_a[20]);
  assign popcount36_ugbo_core_101 = ~(input_a[5] & input_a[29]);
  assign popcount36_ugbo_core_102 = ~(input_a[26] & input_a[30]);
  assign popcount36_ugbo_core_104 = ~(input_a[34] ^ input_a[20]);
  assign popcount36_ugbo_core_105 = input_a[4] | input_a[27];
  assign popcount36_ugbo_core_108 = ~(input_a[11] ^ input_a[32]);
  assign popcount36_ugbo_core_109 = input_a[17] | input_a[26];
  assign popcount36_ugbo_core_111 = ~(input_a[1] & input_a[34]);
  assign popcount36_ugbo_core_112 = input_a[35] & input_a[25];
  assign popcount36_ugbo_core_113 = ~(input_a[26] ^ input_a[10]);
  assign popcount36_ugbo_core_115 = input_a[14] & input_a[3];
  assign popcount36_ugbo_core_116 = input_a[32] & input_a[12];
  assign popcount36_ugbo_core_117 = input_a[12] ^ input_a[9];
  assign popcount36_ugbo_core_118 = input_a[21] ^ input_a[20];
  assign popcount36_ugbo_core_120 = input_a[11] ^ input_a[22];
  assign popcount36_ugbo_core_121 = input_a[0] & input_a[27];
  assign popcount36_ugbo_core_122 = input_a[31] & input_a[12];
  assign popcount36_ugbo_core_123 = ~input_a[4];
  assign popcount36_ugbo_core_124 = ~(input_a[22] ^ input_a[27]);
  assign popcount36_ugbo_core_125 = ~(input_a[12] | input_a[21]);
  assign popcount36_ugbo_core_126 = ~(input_a[30] | input_a[16]);
  assign popcount36_ugbo_core_127 = input_a[19] | input_a[11];
  assign popcount36_ugbo_core_128 = ~input_a[12];
  assign popcount36_ugbo_core_131 = ~(input_a[23] | input_a[31]);
  assign popcount36_ugbo_core_132 = input_a[23] | input_a[1];
  assign popcount36_ugbo_core_133 = ~(input_a[23] & input_a[30]);
  assign popcount36_ugbo_core_134 = ~(input_a[20] ^ input_a[18]);
  assign popcount36_ugbo_core_136 = input_a[34] | input_a[18];
  assign popcount36_ugbo_core_137 = ~(input_a[24] | input_a[31]);
  assign popcount36_ugbo_core_138 = ~(input_a[14] & input_a[29]);
  assign popcount36_ugbo_core_140 = input_a[19] & input_a[15];
  assign popcount36_ugbo_core_141 = ~(input_a[17] & input_a[34]);
  assign popcount36_ugbo_core_143 = ~(input_a[26] & input_a[18]);
  assign popcount36_ugbo_core_145 = ~input_a[25];
  assign popcount36_ugbo_core_146 = ~(input_a[23] ^ input_a[9]);
  assign popcount36_ugbo_core_148 = input_a[3] & input_a[3];
  assign popcount36_ugbo_core_149 = input_a[11] | input_a[20];
  assign popcount36_ugbo_core_151 = ~(input_a[7] | input_a[18]);
  assign popcount36_ugbo_core_152 = input_a[7] ^ input_a[16];
  assign popcount36_ugbo_core_153 = input_a[12] & input_a[20];
  assign popcount36_ugbo_core_154_not = ~input_a[5];
  assign popcount36_ugbo_core_155 = input_a[27] | input_a[34];
  assign popcount36_ugbo_core_156 = ~(input_a[7] & input_a[32]);
  assign popcount36_ugbo_core_157 = ~(input_a[0] & input_a[31]);
  assign popcount36_ugbo_core_160 = input_a[24] | input_a[20];
  assign popcount36_ugbo_core_161 = ~input_a[31];
  assign popcount36_ugbo_core_166 = ~(input_a[25] & input_a[24]);
  assign popcount36_ugbo_core_168 = ~(input_a[18] | input_a[33]);
  assign popcount36_ugbo_core_169 = ~(input_a[3] & input_a[26]);
  assign popcount36_ugbo_core_171 = ~(input_a[2] & input_a[6]);
  assign popcount36_ugbo_core_172 = ~input_a[0];
  assign popcount36_ugbo_core_173 = ~(input_a[2] | input_a[13]);
  assign popcount36_ugbo_core_174 = ~input_a[22];
  assign popcount36_ugbo_core_175 = ~(input_a[23] & input_a[12]);
  assign popcount36_ugbo_core_177 = input_a[7] & input_a[1];
  assign popcount36_ugbo_core_180 = input_a[21] | input_a[29];
  assign popcount36_ugbo_core_181 = input_a[32] | input_a[33];
  assign popcount36_ugbo_core_183 = ~input_a[4];
  assign popcount36_ugbo_core_184 = input_a[9] ^ input_a[25];
  assign popcount36_ugbo_core_185 = ~(input_a[30] | input_a[30]);
  assign popcount36_ugbo_core_186 = input_a[28] | input_a[2];
  assign popcount36_ugbo_core_187_not = ~input_a[22];
  assign popcount36_ugbo_core_188 = ~input_a[18];
  assign popcount36_ugbo_core_189 = ~(input_a[17] | input_a[12]);
  assign popcount36_ugbo_core_191 = ~(input_a[11] | input_a[11]);
  assign popcount36_ugbo_core_192 = ~(input_a[12] ^ input_a[26]);
  assign popcount36_ugbo_core_193 = input_a[5] | input_a[10];
  assign popcount36_ugbo_core_194 = ~(input_a[28] ^ input_a[27]);
  assign popcount36_ugbo_core_195 = ~(input_a[12] | input_a[0]);
  assign popcount36_ugbo_core_196 = ~(input_a[9] | input_a[6]);
  assign popcount36_ugbo_core_197 = ~input_a[0];
  assign popcount36_ugbo_core_198 = ~(input_a[11] ^ input_a[21]);
  assign popcount36_ugbo_core_199 = ~(input_a[22] ^ input_a[17]);
  assign popcount36_ugbo_core_203 = input_a[30] | input_a[30];
  assign popcount36_ugbo_core_204 = ~input_a[28];
  assign popcount36_ugbo_core_205 = ~input_a[7];
  assign popcount36_ugbo_core_206_not = ~input_a[28];
  assign popcount36_ugbo_core_207 = ~(input_a[14] ^ input_a[35]);
  assign popcount36_ugbo_core_210 = ~(input_a[26] & input_a[28]);
  assign popcount36_ugbo_core_211 = ~(input_a[8] & input_a[33]);
  assign popcount36_ugbo_core_213_not = ~input_a[23];
  assign popcount36_ugbo_core_215 = ~(input_a[20] & input_a[25]);
  assign popcount36_ugbo_core_216 = input_a[27] | input_a[0];
  assign popcount36_ugbo_core_217 = ~(input_a[7] ^ input_a[7]);
  assign popcount36_ugbo_core_223 = ~(input_a[26] | input_a[17]);
  assign popcount36_ugbo_core_224 = ~(input_a[27] ^ input_a[30]);
  assign popcount36_ugbo_core_227 = ~(input_a[30] ^ input_a[0]);
  assign popcount36_ugbo_core_229 = ~(input_a[30] & input_a[6]);
  assign popcount36_ugbo_core_231 = input_a[30] | input_a[5];
  assign popcount36_ugbo_core_232 = input_a[15] | input_a[29];
  assign popcount36_ugbo_core_233 = ~(input_a[22] & input_a[11]);
  assign popcount36_ugbo_core_236 = ~input_a[14];
  assign popcount36_ugbo_core_237 = input_a[19] | input_a[26];
  assign popcount36_ugbo_core_238 = ~input_a[12];
  assign popcount36_ugbo_core_240_not = ~input_a[25];
  assign popcount36_ugbo_core_243 = ~(input_a[2] ^ input_a[7]);
  assign popcount36_ugbo_core_245 = ~input_a[35];
  assign popcount36_ugbo_core_247 = input_a[23] & input_a[32];
  assign popcount36_ugbo_core_248 = ~(input_a[19] & input_a[7]);
  assign popcount36_ugbo_core_250 = ~(input_a[24] | input_a[2]);
  assign popcount36_ugbo_core_251_not = ~input_a[20];
  assign popcount36_ugbo_core_252 = ~(input_a[8] ^ input_a[31]);
  assign popcount36_ugbo_core_255 = input_a[13] ^ input_a[12];
  assign popcount36_ugbo_core_256 = ~(input_a[33] | input_a[16]);
  assign popcount36_ugbo_core_257 = ~input_a[19];
  assign popcount36_ugbo_core_261 = ~input_a[12];
  assign popcount36_ugbo_core_262 = ~(input_a[8] | input_a[7]);
  assign popcount36_ugbo_core_263 = ~(input_a[17] ^ input_a[14]);
  assign popcount36_ugbo_core_265 = ~(input_a[35] ^ input_a[9]);
  assign popcount36_ugbo_core_266 = input_a[27] & input_a[8];
  assign popcount36_ugbo_core_267 = ~input_a[9];
  assign popcount36_ugbo_core_268 = input_a[13] & input_a[27];
  assign popcount36_ugbo_core_269 = ~(input_a[5] & input_a[28]);
  assign popcount36_ugbo_core_271 = ~(input_a[11] | input_a[0]);
  assign popcount36_ugbo_core_273 = input_a[4] ^ input_a[35];
  assign popcount36_ugbo_core_274 = ~(input_a[25] ^ input_a[29]);
  assign popcount36_ugbo_core_276_not = ~input_a[3];

  assign popcount36_ugbo_out[0] = input_a[18];
  assign popcount36_ugbo_out[1] = 1'b1;
  assign popcount36_ugbo_out[2] = input_a[22];
  assign popcount36_ugbo_out[3] = 1'b0;
  assign popcount36_ugbo_out[4] = input_a[0];
  assign popcount36_ugbo_out[5] = 1'b0;
endmodule