// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.50741
// WCE=20.0
// EP=0.874629%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_ee7v(input [38:0] input_a, output [5:0] popcount39_ee7v_out);
  wire popcount39_ee7v_core_041;
  wire popcount39_ee7v_core_043;
  wire popcount39_ee7v_core_045;
  wire popcount39_ee7v_core_046;
  wire popcount39_ee7v_core_048;
  wire popcount39_ee7v_core_049;
  wire popcount39_ee7v_core_050;
  wire popcount39_ee7v_core_051;
  wire popcount39_ee7v_core_052;
  wire popcount39_ee7v_core_058;
  wire popcount39_ee7v_core_061;
  wire popcount39_ee7v_core_062;
  wire popcount39_ee7v_core_063;
  wire popcount39_ee7v_core_066_not;
  wire popcount39_ee7v_core_067;
  wire popcount39_ee7v_core_068;
  wire popcount39_ee7v_core_069;
  wire popcount39_ee7v_core_070;
  wire popcount39_ee7v_core_071;
  wire popcount39_ee7v_core_072;
  wire popcount39_ee7v_core_074;
  wire popcount39_ee7v_core_075_not;
  wire popcount39_ee7v_core_076;
  wire popcount39_ee7v_core_077;
  wire popcount39_ee7v_core_078;
  wire popcount39_ee7v_core_085;
  wire popcount39_ee7v_core_086;
  wire popcount39_ee7v_core_088;
  wire popcount39_ee7v_core_091;
  wire popcount39_ee7v_core_092;
  wire popcount39_ee7v_core_093;
  wire popcount39_ee7v_core_095;
  wire popcount39_ee7v_core_096;
  wire popcount39_ee7v_core_097;
  wire popcount39_ee7v_core_100;
  wire popcount39_ee7v_core_103;
  wire popcount39_ee7v_core_105;
  wire popcount39_ee7v_core_106;
  wire popcount39_ee7v_core_107;
  wire popcount39_ee7v_core_108;
  wire popcount39_ee7v_core_109;
  wire popcount39_ee7v_core_110;
  wire popcount39_ee7v_core_111;
  wire popcount39_ee7v_core_112;
  wire popcount39_ee7v_core_114;
  wire popcount39_ee7v_core_116;
  wire popcount39_ee7v_core_117;
  wire popcount39_ee7v_core_118;
  wire popcount39_ee7v_core_123;
  wire popcount39_ee7v_core_124;
  wire popcount39_ee7v_core_125;
  wire popcount39_ee7v_core_129;
  wire popcount39_ee7v_core_130_not;
  wire popcount39_ee7v_core_132_not;
  wire popcount39_ee7v_core_139;
  wire popcount39_ee7v_core_140;
  wire popcount39_ee7v_core_142;
  wire popcount39_ee7v_core_144;
  wire popcount39_ee7v_core_145;
  wire popcount39_ee7v_core_146;
  wire popcount39_ee7v_core_147;
  wire popcount39_ee7v_core_148;
  wire popcount39_ee7v_core_149;
  wire popcount39_ee7v_core_150;
  wire popcount39_ee7v_core_153;
  wire popcount39_ee7v_core_155;
  wire popcount39_ee7v_core_156;
  wire popcount39_ee7v_core_158;
  wire popcount39_ee7v_core_160;
  wire popcount39_ee7v_core_161;
  wire popcount39_ee7v_core_162;
  wire popcount39_ee7v_core_163;
  wire popcount39_ee7v_core_164;
  wire popcount39_ee7v_core_165;
  wire popcount39_ee7v_core_167;
  wire popcount39_ee7v_core_168;
  wire popcount39_ee7v_core_169;
  wire popcount39_ee7v_core_170;
  wire popcount39_ee7v_core_171;
  wire popcount39_ee7v_core_173;
  wire popcount39_ee7v_core_175;
  wire popcount39_ee7v_core_176;
  wire popcount39_ee7v_core_177;
  wire popcount39_ee7v_core_178;
  wire popcount39_ee7v_core_179;
  wire popcount39_ee7v_core_182;
  wire popcount39_ee7v_core_184;
  wire popcount39_ee7v_core_187;
  wire popcount39_ee7v_core_190;
  wire popcount39_ee7v_core_192;
  wire popcount39_ee7v_core_193;
  wire popcount39_ee7v_core_194;
  wire popcount39_ee7v_core_195;
  wire popcount39_ee7v_core_196;
  wire popcount39_ee7v_core_197;
  wire popcount39_ee7v_core_198;
  wire popcount39_ee7v_core_199;
  wire popcount39_ee7v_core_200;
  wire popcount39_ee7v_core_201;
  wire popcount39_ee7v_core_202;
  wire popcount39_ee7v_core_204;
  wire popcount39_ee7v_core_205;
  wire popcount39_ee7v_core_206;
  wire popcount39_ee7v_core_207;
  wire popcount39_ee7v_core_211;
  wire popcount39_ee7v_core_212;
  wire popcount39_ee7v_core_215;
  wire popcount39_ee7v_core_217;
  wire popcount39_ee7v_core_218;
  wire popcount39_ee7v_core_220;
  wire popcount39_ee7v_core_223;
  wire popcount39_ee7v_core_225;
  wire popcount39_ee7v_core_226;
  wire popcount39_ee7v_core_227;
  wire popcount39_ee7v_core_231;
  wire popcount39_ee7v_core_232;
  wire popcount39_ee7v_core_233;
  wire popcount39_ee7v_core_235;
  wire popcount39_ee7v_core_236;
  wire popcount39_ee7v_core_239;
  wire popcount39_ee7v_core_242;
  wire popcount39_ee7v_core_243;
  wire popcount39_ee7v_core_246;
  wire popcount39_ee7v_core_247;
  wire popcount39_ee7v_core_249;
  wire popcount39_ee7v_core_250;
  wire popcount39_ee7v_core_256;
  wire popcount39_ee7v_core_257;
  wire popcount39_ee7v_core_258;
  wire popcount39_ee7v_core_259;
  wire popcount39_ee7v_core_260;
  wire popcount39_ee7v_core_261;
  wire popcount39_ee7v_core_262;
  wire popcount39_ee7v_core_263;
  wire popcount39_ee7v_core_264;
  wire popcount39_ee7v_core_265;
  wire popcount39_ee7v_core_266;
  wire popcount39_ee7v_core_267;
  wire popcount39_ee7v_core_270;
  wire popcount39_ee7v_core_271;
  wire popcount39_ee7v_core_272;
  wire popcount39_ee7v_core_273;
  wire popcount39_ee7v_core_274;
  wire popcount39_ee7v_core_275;
  wire popcount39_ee7v_core_276;
  wire popcount39_ee7v_core_277_not;
  wire popcount39_ee7v_core_278;
  wire popcount39_ee7v_core_282;
  wire popcount39_ee7v_core_283;
  wire popcount39_ee7v_core_285;
  wire popcount39_ee7v_core_286;
  wire popcount39_ee7v_core_287;
  wire popcount39_ee7v_core_288;
  wire popcount39_ee7v_core_289;
  wire popcount39_ee7v_core_291;
  wire popcount39_ee7v_core_292;
  wire popcount39_ee7v_core_294;
  wire popcount39_ee7v_core_295;
  wire popcount39_ee7v_core_296;
  wire popcount39_ee7v_core_297;
  wire popcount39_ee7v_core_298;
  wire popcount39_ee7v_core_299;
  wire popcount39_ee7v_core_300;
  wire popcount39_ee7v_core_303;
  wire popcount39_ee7v_core_304;
  wire popcount39_ee7v_core_305;

  assign popcount39_ee7v_core_041 = ~(input_a[34] & input_a[31]);
  assign popcount39_ee7v_core_043 = ~(input_a[11] ^ input_a[9]);
  assign popcount39_ee7v_core_045 = ~(input_a[34] ^ input_a[14]);
  assign popcount39_ee7v_core_046 = ~(input_a[7] & input_a[14]);
  assign popcount39_ee7v_core_048 = input_a[30] | input_a[36];
  assign popcount39_ee7v_core_049 = input_a[38] & input_a[16];
  assign popcount39_ee7v_core_050 = input_a[1] & input_a[34];
  assign popcount39_ee7v_core_051 = input_a[15] | input_a[33];
  assign popcount39_ee7v_core_052 = ~(input_a[28] | input_a[30]);
  assign popcount39_ee7v_core_058 = ~(input_a[10] & input_a[27]);
  assign popcount39_ee7v_core_061 = ~input_a[23];
  assign popcount39_ee7v_core_062 = ~(input_a[9] | input_a[31]);
  assign popcount39_ee7v_core_063 = ~input_a[12];
  assign popcount39_ee7v_core_066_not = ~input_a[6];
  assign popcount39_ee7v_core_067 = ~(input_a[15] & input_a[23]);
  assign popcount39_ee7v_core_068 = ~(input_a[18] | input_a[27]);
  assign popcount39_ee7v_core_069 = input_a[18] & input_a[2];
  assign popcount39_ee7v_core_070 = ~input_a[28];
  assign popcount39_ee7v_core_071 = input_a[17] & input_a[36];
  assign popcount39_ee7v_core_072 = input_a[32] | input_a[32];
  assign popcount39_ee7v_core_074 = ~(input_a[26] ^ input_a[3]);
  assign popcount39_ee7v_core_075_not = ~input_a[30];
  assign popcount39_ee7v_core_076 = input_a[5] | input_a[31];
  assign popcount39_ee7v_core_077 = input_a[0] ^ input_a[24];
  assign popcount39_ee7v_core_078 = input_a[34] & input_a[1];
  assign popcount39_ee7v_core_085 = ~(input_a[28] & input_a[7]);
  assign popcount39_ee7v_core_086 = input_a[34] & input_a[31];
  assign popcount39_ee7v_core_088 = ~(input_a[31] ^ input_a[15]);
  assign popcount39_ee7v_core_091 = input_a[33] | input_a[31];
  assign popcount39_ee7v_core_092 = ~input_a[37];
  assign popcount39_ee7v_core_093 = ~(input_a[22] & input_a[17]);
  assign popcount39_ee7v_core_095 = ~(input_a[0] & input_a[8]);
  assign popcount39_ee7v_core_096 = input_a[19] & input_a[13];
  assign popcount39_ee7v_core_097 = input_a[27] ^ input_a[5];
  assign popcount39_ee7v_core_100 = ~(input_a[18] ^ input_a[16]);
  assign popcount39_ee7v_core_103 = ~(input_a[11] | input_a[0]);
  assign popcount39_ee7v_core_105 = input_a[32] ^ input_a[2];
  assign popcount39_ee7v_core_106 = ~(input_a[31] & input_a[30]);
  assign popcount39_ee7v_core_107 = input_a[28] | input_a[3];
  assign popcount39_ee7v_core_108 = ~(input_a[4] & input_a[38]);
  assign popcount39_ee7v_core_109 = input_a[23] & input_a[8];
  assign popcount39_ee7v_core_110 = input_a[26] & input_a[27];
  assign popcount39_ee7v_core_111 = ~(input_a[20] | input_a[34]);
  assign popcount39_ee7v_core_112 = ~(input_a[10] ^ input_a[22]);
  assign popcount39_ee7v_core_114 = ~(input_a[0] & input_a[25]);
  assign popcount39_ee7v_core_116 = input_a[25] & input_a[11];
  assign popcount39_ee7v_core_117 = input_a[24] ^ input_a[1];
  assign popcount39_ee7v_core_118 = ~(input_a[4] ^ input_a[3]);
  assign popcount39_ee7v_core_123 = input_a[17] | input_a[9];
  assign popcount39_ee7v_core_124 = ~(input_a[16] | input_a[36]);
  assign popcount39_ee7v_core_125 = input_a[11] & input_a[3];
  assign popcount39_ee7v_core_129 = input_a[36] & input_a[14];
  assign popcount39_ee7v_core_130_not = ~input_a[35];
  assign popcount39_ee7v_core_132_not = ~input_a[21];
  assign popcount39_ee7v_core_139 = ~(input_a[1] & input_a[22]);
  assign popcount39_ee7v_core_140 = ~(input_a[17] & input_a[11]);
  assign popcount39_ee7v_core_142 = ~(input_a[20] & input_a[27]);
  assign popcount39_ee7v_core_144 = input_a[19] | input_a[1];
  assign popcount39_ee7v_core_145 = ~(input_a[33] ^ input_a[7]);
  assign popcount39_ee7v_core_146 = input_a[13] & input_a[24];
  assign popcount39_ee7v_core_147 = input_a[10] & input_a[4];
  assign popcount39_ee7v_core_148 = ~(input_a[3] & input_a[21]);
  assign popcount39_ee7v_core_149 = ~(input_a[13] | input_a[32]);
  assign popcount39_ee7v_core_150 = input_a[18] ^ input_a[9];
  assign popcount39_ee7v_core_153 = input_a[22] | input_a[21];
  assign popcount39_ee7v_core_155 = input_a[22] | input_a[36];
  assign popcount39_ee7v_core_156 = input_a[25] & input_a[22];
  assign popcount39_ee7v_core_158 = ~input_a[3];
  assign popcount39_ee7v_core_160 = ~input_a[37];
  assign popcount39_ee7v_core_161 = input_a[23] | input_a[32];
  assign popcount39_ee7v_core_162 = ~(input_a[34] | input_a[30]);
  assign popcount39_ee7v_core_163 = input_a[29] | input_a[10];
  assign popcount39_ee7v_core_164 = ~(input_a[5] & input_a[17]);
  assign popcount39_ee7v_core_165 = ~(input_a[23] ^ input_a[26]);
  assign popcount39_ee7v_core_167 = ~input_a[29];
  assign popcount39_ee7v_core_168 = ~(input_a[0] & input_a[31]);
  assign popcount39_ee7v_core_169 = ~(input_a[19] | input_a[17]);
  assign popcount39_ee7v_core_170 = input_a[11] & input_a[34];
  assign popcount39_ee7v_core_171 = ~(input_a[29] & input_a[36]);
  assign popcount39_ee7v_core_173 = input_a[20] | input_a[8];
  assign popcount39_ee7v_core_175 = ~input_a[7];
  assign popcount39_ee7v_core_176 = ~(input_a[34] | input_a[21]);
  assign popcount39_ee7v_core_177 = ~(input_a[25] ^ input_a[11]);
  assign popcount39_ee7v_core_178 = ~(input_a[0] & input_a[30]);
  assign popcount39_ee7v_core_179 = ~(input_a[4] ^ input_a[10]);
  assign popcount39_ee7v_core_182 = ~(input_a[15] | input_a[11]);
  assign popcount39_ee7v_core_184 = ~(input_a[10] | input_a[8]);
  assign popcount39_ee7v_core_187 = ~input_a[16];
  assign popcount39_ee7v_core_190 = input_a[19] | input_a[38];
  assign popcount39_ee7v_core_192 = ~(input_a[5] & input_a[15]);
  assign popcount39_ee7v_core_193 = ~(input_a[29] ^ input_a[3]);
  assign popcount39_ee7v_core_194 = ~(input_a[28] ^ input_a[25]);
  assign popcount39_ee7v_core_195 = ~(input_a[29] | input_a[23]);
  assign popcount39_ee7v_core_196 = input_a[13] | input_a[0];
  assign popcount39_ee7v_core_197 = ~(input_a[38] | input_a[29]);
  assign popcount39_ee7v_core_198 = input_a[27] & input_a[1];
  assign popcount39_ee7v_core_199 = ~input_a[1];
  assign popcount39_ee7v_core_200 = ~(input_a[25] | input_a[13]);
  assign popcount39_ee7v_core_201 = ~input_a[20];
  assign popcount39_ee7v_core_202 = input_a[24] ^ input_a[3];
  assign popcount39_ee7v_core_204 = ~(input_a[14] | input_a[4]);
  assign popcount39_ee7v_core_205 = ~(input_a[32] | input_a[16]);
  assign popcount39_ee7v_core_206 = input_a[34] ^ input_a[7];
  assign popcount39_ee7v_core_207 = ~(input_a[1] | input_a[26]);
  assign popcount39_ee7v_core_211 = ~(input_a[23] ^ input_a[14]);
  assign popcount39_ee7v_core_212 = ~(input_a[4] & input_a[16]);
  assign popcount39_ee7v_core_215 = input_a[4] & input_a[10];
  assign popcount39_ee7v_core_217 = ~(input_a[7] & input_a[10]);
  assign popcount39_ee7v_core_218 = input_a[28] ^ input_a[38];
  assign popcount39_ee7v_core_220 = input_a[13] & input_a[37];
  assign popcount39_ee7v_core_223 = input_a[17] ^ input_a[15];
  assign popcount39_ee7v_core_225 = ~(input_a[6] | input_a[20]);
  assign popcount39_ee7v_core_226 = ~(input_a[31] ^ input_a[12]);
  assign popcount39_ee7v_core_227 = input_a[11] & input_a[21];
  assign popcount39_ee7v_core_231 = ~(input_a[28] ^ input_a[14]);
  assign popcount39_ee7v_core_232 = ~(input_a[6] | input_a[26]);
  assign popcount39_ee7v_core_233 = ~(input_a[24] & input_a[18]);
  assign popcount39_ee7v_core_235 = input_a[11] | input_a[26];
  assign popcount39_ee7v_core_236 = input_a[23] | input_a[4];
  assign popcount39_ee7v_core_239 = ~input_a[16];
  assign popcount39_ee7v_core_242 = ~(input_a[25] ^ input_a[9]);
  assign popcount39_ee7v_core_243 = ~input_a[23];
  assign popcount39_ee7v_core_246 = ~input_a[30];
  assign popcount39_ee7v_core_247 = input_a[16] & input_a[13];
  assign popcount39_ee7v_core_249 = ~(input_a[32] | input_a[3]);
  assign popcount39_ee7v_core_250 = ~input_a[18];
  assign popcount39_ee7v_core_256 = input_a[21] | input_a[13];
  assign popcount39_ee7v_core_257 = ~(input_a[7] ^ input_a[35]);
  assign popcount39_ee7v_core_258 = ~(input_a[13] ^ input_a[23]);
  assign popcount39_ee7v_core_259 = input_a[13] ^ input_a[34];
  assign popcount39_ee7v_core_260 = input_a[12] & input_a[18];
  assign popcount39_ee7v_core_261 = input_a[21] & input_a[7];
  assign popcount39_ee7v_core_262 = ~(input_a[25] & input_a[11]);
  assign popcount39_ee7v_core_263 = ~input_a[17];
  assign popcount39_ee7v_core_264 = input_a[13] & input_a[9];
  assign popcount39_ee7v_core_265 = ~(input_a[5] | input_a[21]);
  assign popcount39_ee7v_core_266 = ~(input_a[1] | input_a[27]);
  assign popcount39_ee7v_core_267 = ~(input_a[9] ^ input_a[16]);
  assign popcount39_ee7v_core_270 = input_a[38] ^ input_a[6];
  assign popcount39_ee7v_core_271 = input_a[26] | input_a[22];
  assign popcount39_ee7v_core_272 = input_a[2] & input_a[35];
  assign popcount39_ee7v_core_273 = input_a[38] ^ input_a[31];
  assign popcount39_ee7v_core_274 = ~(input_a[13] ^ input_a[25]);
  assign popcount39_ee7v_core_275 = ~(input_a[12] | input_a[1]);
  assign popcount39_ee7v_core_276 = ~(input_a[9] | input_a[27]);
  assign popcount39_ee7v_core_277_not = ~input_a[9];
  assign popcount39_ee7v_core_278 = ~(input_a[13] | input_a[18]);
  assign popcount39_ee7v_core_282 = ~(input_a[18] ^ input_a[34]);
  assign popcount39_ee7v_core_283 = ~(input_a[17] ^ input_a[20]);
  assign popcount39_ee7v_core_285 = ~(input_a[21] & input_a[25]);
  assign popcount39_ee7v_core_286 = ~(input_a[37] ^ input_a[31]);
  assign popcount39_ee7v_core_287 = input_a[9] & input_a[19];
  assign popcount39_ee7v_core_288 = ~(input_a[4] ^ input_a[23]);
  assign popcount39_ee7v_core_289 = input_a[2] & input_a[21];
  assign popcount39_ee7v_core_291 = input_a[8] & input_a[2];
  assign popcount39_ee7v_core_292 = input_a[16] ^ input_a[15];
  assign popcount39_ee7v_core_294 = input_a[17] & input_a[37];
  assign popcount39_ee7v_core_295 = ~(input_a[18] ^ input_a[34]);
  assign popcount39_ee7v_core_296 = input_a[25] | input_a[13];
  assign popcount39_ee7v_core_297 = input_a[34] | input_a[29];
  assign popcount39_ee7v_core_298 = input_a[27] ^ input_a[26];
  assign popcount39_ee7v_core_299 = ~(input_a[29] ^ input_a[8]);
  assign popcount39_ee7v_core_300 = ~(input_a[36] ^ input_a[24]);
  assign popcount39_ee7v_core_303 = ~(input_a[31] | input_a[24]);
  assign popcount39_ee7v_core_304 = ~(input_a[21] ^ input_a[6]);
  assign popcount39_ee7v_core_305 = ~(input_a[26] ^ input_a[2]);

  assign popcount39_ee7v_out[0] = 1'b0;
  assign popcount39_ee7v_out[1] = 1'b0;
  assign popcount39_ee7v_out[2] = 1'b1;
  assign popcount39_ee7v_out[3] = 1'b0;
  assign popcount39_ee7v_out[4] = 1'b1;
  assign popcount39_ee7v_out[5] = 1'b0;
endmodule