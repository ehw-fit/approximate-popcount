// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.53964
// WCE=28.0
// EP=0.986587%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_030e(input [37:0] input_a, output [5:0] popcount38_030e_out);
  wire popcount38_030e_core_042;
  wire popcount38_030e_core_043;
  wire popcount38_030e_core_044;
  wire popcount38_030e_core_047;
  wire popcount38_030e_core_048;
  wire popcount38_030e_core_049;
  wire popcount38_030e_core_050;
  wire popcount38_030e_core_051;
  wire popcount38_030e_core_052;
  wire popcount38_030e_core_053;
  wire popcount38_030e_core_057;
  wire popcount38_030e_core_058;
  wire popcount38_030e_core_060;
  wire popcount38_030e_core_063_not;
  wire popcount38_030e_core_065;
  wire popcount38_030e_core_066;
  wire popcount38_030e_core_068;
  wire popcount38_030e_core_069;
  wire popcount38_030e_core_070;
  wire popcount38_030e_core_073;
  wire popcount38_030e_core_075;
  wire popcount38_030e_core_077;
  wire popcount38_030e_core_079;
  wire popcount38_030e_core_081;
  wire popcount38_030e_core_084;
  wire popcount38_030e_core_085;
  wire popcount38_030e_core_087;
  wire popcount38_030e_core_088;
  wire popcount38_030e_core_089;
  wire popcount38_030e_core_091;
  wire popcount38_030e_core_093;
  wire popcount38_030e_core_094;
  wire popcount38_030e_core_095;
  wire popcount38_030e_core_096;
  wire popcount38_030e_core_097;
  wire popcount38_030e_core_098;
  wire popcount38_030e_core_101;
  wire popcount38_030e_core_102;
  wire popcount38_030e_core_104;
  wire popcount38_030e_core_106;
  wire popcount38_030e_core_110;
  wire popcount38_030e_core_111;
  wire popcount38_030e_core_112;
  wire popcount38_030e_core_113;
  wire popcount38_030e_core_114;
  wire popcount38_030e_core_117;
  wire popcount38_030e_core_118;
  wire popcount38_030e_core_119;
  wire popcount38_030e_core_120;
  wire popcount38_030e_core_121;
  wire popcount38_030e_core_124;
  wire popcount38_030e_core_125;
  wire popcount38_030e_core_127;
  wire popcount38_030e_core_129;
  wire popcount38_030e_core_130;
  wire popcount38_030e_core_132;
  wire popcount38_030e_core_134;
  wire popcount38_030e_core_135;
  wire popcount38_030e_core_136;
  wire popcount38_030e_core_137;
  wire popcount38_030e_core_139;
  wire popcount38_030e_core_140;
  wire popcount38_030e_core_141;
  wire popcount38_030e_core_143;
  wire popcount38_030e_core_144;
  wire popcount38_030e_core_146;
  wire popcount38_030e_core_147;
  wire popcount38_030e_core_149;
  wire popcount38_030e_core_151;
  wire popcount38_030e_core_152;
  wire popcount38_030e_core_153;
  wire popcount38_030e_core_154;
  wire popcount38_030e_core_155;
  wire popcount38_030e_core_156;
  wire popcount38_030e_core_157;
  wire popcount38_030e_core_159_not;
  wire popcount38_030e_core_161;
  wire popcount38_030e_core_163;
  wire popcount38_030e_core_166;
  wire popcount38_030e_core_167;
  wire popcount38_030e_core_169;
  wire popcount38_030e_core_172;
  wire popcount38_030e_core_173;
  wire popcount38_030e_core_174;
  wire popcount38_030e_core_176;
  wire popcount38_030e_core_177;
  wire popcount38_030e_core_178;
  wire popcount38_030e_core_179;
  wire popcount38_030e_core_181;
  wire popcount38_030e_core_183;
  wire popcount38_030e_core_184;
  wire popcount38_030e_core_186;
  wire popcount38_030e_core_187;
  wire popcount38_030e_core_188;
  wire popcount38_030e_core_190;
  wire popcount38_030e_core_195;
  wire popcount38_030e_core_196;
  wire popcount38_030e_core_197;
  wire popcount38_030e_core_199;
  wire popcount38_030e_core_201;
  wire popcount38_030e_core_202;
  wire popcount38_030e_core_204;
  wire popcount38_030e_core_205;
  wire popcount38_030e_core_207;
  wire popcount38_030e_core_208;
  wire popcount38_030e_core_209;
  wire popcount38_030e_core_211;
  wire popcount38_030e_core_212;
  wire popcount38_030e_core_213;
  wire popcount38_030e_core_216;
  wire popcount38_030e_core_217;
  wire popcount38_030e_core_218;
  wire popcount38_030e_core_219;
  wire popcount38_030e_core_222;
  wire popcount38_030e_core_223;
  wire popcount38_030e_core_225;
  wire popcount38_030e_core_226;
  wire popcount38_030e_core_227;
  wire popcount38_030e_core_228;
  wire popcount38_030e_core_230;
  wire popcount38_030e_core_231_not;
  wire popcount38_030e_core_233;
  wire popcount38_030e_core_235;
  wire popcount38_030e_core_236;
  wire popcount38_030e_core_239;
  wire popcount38_030e_core_240;
  wire popcount38_030e_core_242;
  wire popcount38_030e_core_247;
  wire popcount38_030e_core_248;
  wire popcount38_030e_core_250;
  wire popcount38_030e_core_252;
  wire popcount38_030e_core_253;
  wire popcount38_030e_core_256;
  wire popcount38_030e_core_259;
  wire popcount38_030e_core_260;
  wire popcount38_030e_core_261;
  wire popcount38_030e_core_263;
  wire popcount38_030e_core_267;
  wire popcount38_030e_core_268;
  wire popcount38_030e_core_269;
  wire popcount38_030e_core_270;
  wire popcount38_030e_core_271;
  wire popcount38_030e_core_272;
  wire popcount38_030e_core_274;
  wire popcount38_030e_core_275;
  wire popcount38_030e_core_276;
  wire popcount38_030e_core_278;
  wire popcount38_030e_core_279;
  wire popcount38_030e_core_280;
  wire popcount38_030e_core_282;
  wire popcount38_030e_core_283;
  wire popcount38_030e_core_285;
  wire popcount38_030e_core_286;
  wire popcount38_030e_core_288;
  wire popcount38_030e_core_290;
  wire popcount38_030e_core_291;
  wire popcount38_030e_core_292;
  wire popcount38_030e_core_294;
  wire popcount38_030e_core_296;

  assign popcount38_030e_core_042 = input_a[28] ^ input_a[32];
  assign popcount38_030e_core_043 = input_a[30] ^ input_a[8];
  assign popcount38_030e_core_044 = ~(input_a[37] ^ input_a[24]);
  assign popcount38_030e_core_047 = input_a[15] | input_a[32];
  assign popcount38_030e_core_048 = input_a[8] & input_a[34];
  assign popcount38_030e_core_049 = ~(input_a[32] ^ input_a[1]);
  assign popcount38_030e_core_050 = input_a[26] ^ input_a[6];
  assign popcount38_030e_core_051 = ~(input_a[1] | input_a[4]);
  assign popcount38_030e_core_052 = input_a[36] & input_a[24];
  assign popcount38_030e_core_053 = ~(input_a[4] | input_a[7]);
  assign popcount38_030e_core_057 = ~(input_a[12] ^ input_a[17]);
  assign popcount38_030e_core_058 = input_a[28] | input_a[29];
  assign popcount38_030e_core_060 = ~(input_a[26] ^ input_a[16]);
  assign popcount38_030e_core_063_not = ~input_a[32];
  assign popcount38_030e_core_065 = input_a[25] | input_a[4];
  assign popcount38_030e_core_066 = ~(input_a[37] & input_a[1]);
  assign popcount38_030e_core_068 = input_a[1] ^ input_a[23];
  assign popcount38_030e_core_069 = ~(input_a[2] | input_a[12]);
  assign popcount38_030e_core_070 = ~input_a[5];
  assign popcount38_030e_core_073 = ~input_a[6];
  assign popcount38_030e_core_075 = ~(input_a[25] & input_a[35]);
  assign popcount38_030e_core_077 = ~input_a[6];
  assign popcount38_030e_core_079 = ~(input_a[6] | input_a[4]);
  assign popcount38_030e_core_081 = ~(input_a[10] | input_a[23]);
  assign popcount38_030e_core_084 = input_a[8] ^ input_a[8];
  assign popcount38_030e_core_085 = ~(input_a[17] & input_a[18]);
  assign popcount38_030e_core_087 = ~input_a[26];
  assign popcount38_030e_core_088 = input_a[22] & input_a[20];
  assign popcount38_030e_core_089 = ~input_a[2];
  assign popcount38_030e_core_091 = input_a[12] | input_a[7];
  assign popcount38_030e_core_093 = input_a[14] & input_a[20];
  assign popcount38_030e_core_094 = ~(input_a[4] ^ input_a[10]);
  assign popcount38_030e_core_095 = input_a[7] ^ input_a[1];
  assign popcount38_030e_core_096 = ~(input_a[22] & input_a[1]);
  assign popcount38_030e_core_097 = input_a[13] | input_a[1];
  assign popcount38_030e_core_098 = ~(input_a[30] ^ input_a[19]);
  assign popcount38_030e_core_101 = ~input_a[27];
  assign popcount38_030e_core_102 = ~(input_a[23] | input_a[11]);
  assign popcount38_030e_core_104 = ~(input_a[17] ^ input_a[35]);
  assign popcount38_030e_core_106 = ~(input_a[4] | input_a[33]);
  assign popcount38_030e_core_110 = ~(input_a[6] ^ input_a[4]);
  assign popcount38_030e_core_111 = ~(input_a[1] & input_a[20]);
  assign popcount38_030e_core_112 = input_a[20] & input_a[29];
  assign popcount38_030e_core_113 = ~input_a[8];
  assign popcount38_030e_core_114 = ~(input_a[21] | input_a[9]);
  assign popcount38_030e_core_117 = input_a[5] | input_a[14];
  assign popcount38_030e_core_118 = input_a[25] | input_a[33];
  assign popcount38_030e_core_119 = ~(input_a[31] | input_a[36]);
  assign popcount38_030e_core_120 = input_a[29] & input_a[27];
  assign popcount38_030e_core_121 = input_a[10] ^ input_a[9];
  assign popcount38_030e_core_124 = ~input_a[8];
  assign popcount38_030e_core_125 = input_a[32] ^ input_a[32];
  assign popcount38_030e_core_127 = input_a[21] ^ input_a[34];
  assign popcount38_030e_core_129 = input_a[37] | input_a[13];
  assign popcount38_030e_core_130 = ~(input_a[0] | input_a[36]);
  assign popcount38_030e_core_132 = ~(input_a[3] | input_a[10]);
  assign popcount38_030e_core_134 = input_a[17] & input_a[11];
  assign popcount38_030e_core_135 = input_a[21] & input_a[34];
  assign popcount38_030e_core_136 = input_a[1] | input_a[33];
  assign popcount38_030e_core_137 = ~(input_a[14] ^ input_a[16]);
  assign popcount38_030e_core_139 = ~input_a[13];
  assign popcount38_030e_core_140 = ~(input_a[12] ^ input_a[31]);
  assign popcount38_030e_core_141 = input_a[27] ^ input_a[3];
  assign popcount38_030e_core_143 = ~(input_a[11] ^ input_a[37]);
  assign popcount38_030e_core_144 = input_a[20] ^ input_a[4];
  assign popcount38_030e_core_146 = input_a[25] | input_a[14];
  assign popcount38_030e_core_147 = ~input_a[11];
  assign popcount38_030e_core_149 = input_a[32] & input_a[9];
  assign popcount38_030e_core_151 = ~(input_a[5] & input_a[30]);
  assign popcount38_030e_core_152 = ~(input_a[17] & input_a[30]);
  assign popcount38_030e_core_153 = ~input_a[8];
  assign popcount38_030e_core_154 = ~(input_a[5] ^ input_a[27]);
  assign popcount38_030e_core_155 = input_a[31] | input_a[23];
  assign popcount38_030e_core_156 = input_a[20] | input_a[16];
  assign popcount38_030e_core_157 = input_a[15] ^ input_a[24];
  assign popcount38_030e_core_159_not = ~input_a[4];
  assign popcount38_030e_core_161 = ~(input_a[33] | input_a[16]);
  assign popcount38_030e_core_163 = ~(input_a[27] ^ input_a[23]);
  assign popcount38_030e_core_166 = ~(input_a[9] | input_a[19]);
  assign popcount38_030e_core_167 = ~(input_a[15] & input_a[28]);
  assign popcount38_030e_core_169 = ~input_a[1];
  assign popcount38_030e_core_172 = ~(input_a[11] | input_a[17]);
  assign popcount38_030e_core_173 = ~input_a[10];
  assign popcount38_030e_core_174 = ~(input_a[35] | input_a[17]);
  assign popcount38_030e_core_176 = input_a[4] ^ input_a[32];
  assign popcount38_030e_core_177 = ~(input_a[37] | input_a[32]);
  assign popcount38_030e_core_178 = input_a[17] | input_a[15];
  assign popcount38_030e_core_179 = ~(input_a[37] | input_a[28]);
  assign popcount38_030e_core_181 = input_a[22] & input_a[5];
  assign popcount38_030e_core_183 = ~(input_a[21] & input_a[24]);
  assign popcount38_030e_core_184 = input_a[34] & input_a[11];
  assign popcount38_030e_core_186 = ~(input_a[31] & input_a[9]);
  assign popcount38_030e_core_187 = input_a[0] ^ input_a[17];
  assign popcount38_030e_core_188 = ~(input_a[16] & input_a[25]);
  assign popcount38_030e_core_190 = ~(input_a[25] ^ input_a[23]);
  assign popcount38_030e_core_195 = input_a[16] & input_a[37];
  assign popcount38_030e_core_196 = ~(input_a[13] ^ input_a[1]);
  assign popcount38_030e_core_197 = ~(input_a[15] | input_a[19]);
  assign popcount38_030e_core_199 = ~(input_a[24] ^ input_a[5]);
  assign popcount38_030e_core_201 = ~input_a[12];
  assign popcount38_030e_core_202 = input_a[29] | input_a[16];
  assign popcount38_030e_core_204 = ~(input_a[11] | input_a[36]);
  assign popcount38_030e_core_205 = input_a[26] | input_a[33];
  assign popcount38_030e_core_207 = input_a[2] | input_a[6];
  assign popcount38_030e_core_208 = ~(input_a[30] & input_a[21]);
  assign popcount38_030e_core_209 = input_a[7] & input_a[36];
  assign popcount38_030e_core_211 = ~(input_a[33] | input_a[31]);
  assign popcount38_030e_core_212 = input_a[32] ^ input_a[4];
  assign popcount38_030e_core_213 = ~input_a[37];
  assign popcount38_030e_core_216 = input_a[24] ^ input_a[8];
  assign popcount38_030e_core_217 = ~(input_a[17] ^ input_a[12]);
  assign popcount38_030e_core_218 = input_a[16] | input_a[2];
  assign popcount38_030e_core_219 = input_a[35] | input_a[14];
  assign popcount38_030e_core_222 = ~(input_a[22] ^ input_a[5]);
  assign popcount38_030e_core_223 = ~input_a[19];
  assign popcount38_030e_core_225 = ~input_a[29];
  assign popcount38_030e_core_226 = ~(input_a[20] ^ input_a[9]);
  assign popcount38_030e_core_227 = ~(input_a[22] & input_a[29]);
  assign popcount38_030e_core_228 = input_a[37] | input_a[25];
  assign popcount38_030e_core_230 = input_a[13] & input_a[31];
  assign popcount38_030e_core_231_not = ~input_a[2];
  assign popcount38_030e_core_233 = ~(input_a[7] & input_a[11]);
  assign popcount38_030e_core_235 = input_a[31] | input_a[28];
  assign popcount38_030e_core_236 = input_a[8] | input_a[20];
  assign popcount38_030e_core_239 = input_a[36] & input_a[26];
  assign popcount38_030e_core_240 = input_a[18] | input_a[37];
  assign popcount38_030e_core_242 = ~(input_a[36] | input_a[18]);
  assign popcount38_030e_core_247 = input_a[11] & input_a[13];
  assign popcount38_030e_core_248 = ~(input_a[8] & input_a[30]);
  assign popcount38_030e_core_250 = ~(input_a[31] & input_a[4]);
  assign popcount38_030e_core_252 = input_a[14] | input_a[14];
  assign popcount38_030e_core_253 = ~(input_a[22] | input_a[19]);
  assign popcount38_030e_core_256 = ~(input_a[4] ^ input_a[34]);
  assign popcount38_030e_core_259 = ~(input_a[3] & input_a[20]);
  assign popcount38_030e_core_260 = input_a[12] ^ input_a[8];
  assign popcount38_030e_core_261 = ~input_a[7];
  assign popcount38_030e_core_263 = ~(input_a[14] & input_a[30]);
  assign popcount38_030e_core_267 = ~(input_a[29] ^ input_a[5]);
  assign popcount38_030e_core_268 = input_a[31] ^ input_a[19];
  assign popcount38_030e_core_269 = ~(input_a[21] ^ input_a[15]);
  assign popcount38_030e_core_270 = input_a[23] | input_a[32];
  assign popcount38_030e_core_271 = input_a[23] ^ input_a[6];
  assign popcount38_030e_core_272 = ~(input_a[12] & input_a[28]);
  assign popcount38_030e_core_274 = input_a[2] | input_a[4];
  assign popcount38_030e_core_275 = ~(input_a[12] ^ input_a[29]);
  assign popcount38_030e_core_276 = ~input_a[29];
  assign popcount38_030e_core_278 = ~(input_a[12] & input_a[26]);
  assign popcount38_030e_core_279 = ~(input_a[1] | input_a[33]);
  assign popcount38_030e_core_280 = input_a[19] ^ input_a[37];
  assign popcount38_030e_core_282 = ~(input_a[18] ^ input_a[8]);
  assign popcount38_030e_core_283 = input_a[37] & input_a[24];
  assign popcount38_030e_core_285 = input_a[12] & input_a[34];
  assign popcount38_030e_core_286 = input_a[18] | input_a[12];
  assign popcount38_030e_core_288 = input_a[8] ^ input_a[33];
  assign popcount38_030e_core_290 = ~(input_a[5] | input_a[4]);
  assign popcount38_030e_core_291 = ~(input_a[2] ^ input_a[36]);
  assign popcount38_030e_core_292 = input_a[23] | input_a[7];
  assign popcount38_030e_core_294 = input_a[22] | input_a[7];
  assign popcount38_030e_core_296 = input_a[29] | input_a[2];

  assign popcount38_030e_out[0] = input_a[23];
  assign popcount38_030e_out[1] = input_a[25];
  assign popcount38_030e_out[2] = 1'b1;
  assign popcount38_030e_out[3] = 1'b1;
  assign popcount38_030e_out[4] = 1'b0;
  assign popcount38_030e_out[5] = 1'b0;
endmodule