// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=19.5143
// WCE=59.0
// EP=0.994645%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount40_ghhv(input [39:0] input_a, output [5:0] popcount40_ghhv_out);
  wire popcount40_ghhv_core_042;
  wire popcount40_ghhv_core_043_not;
  wire popcount40_ghhv_core_047;
  wire popcount40_ghhv_core_048;
  wire popcount40_ghhv_core_049;
  wire popcount40_ghhv_core_051;
  wire popcount40_ghhv_core_055;
  wire popcount40_ghhv_core_056;
  wire popcount40_ghhv_core_057;
  wire popcount40_ghhv_core_058;
  wire popcount40_ghhv_core_059;
  wire popcount40_ghhv_core_061;
  wire popcount40_ghhv_core_063;
  wire popcount40_ghhv_core_064;
  wire popcount40_ghhv_core_065;
  wire popcount40_ghhv_core_067;
  wire popcount40_ghhv_core_069;
  wire popcount40_ghhv_core_070;
  wire popcount40_ghhv_core_072;
  wire popcount40_ghhv_core_073;
  wire popcount40_ghhv_core_075;
  wire popcount40_ghhv_core_076;
  wire popcount40_ghhv_core_077;
  wire popcount40_ghhv_core_079;
  wire popcount40_ghhv_core_080;
  wire popcount40_ghhv_core_084;
  wire popcount40_ghhv_core_085;
  wire popcount40_ghhv_core_086;
  wire popcount40_ghhv_core_088_not;
  wire popcount40_ghhv_core_089;
  wire popcount40_ghhv_core_090;
  wire popcount40_ghhv_core_092;
  wire popcount40_ghhv_core_093;
  wire popcount40_ghhv_core_094;
  wire popcount40_ghhv_core_098;
  wire popcount40_ghhv_core_099;
  wire popcount40_ghhv_core_100;
  wire popcount40_ghhv_core_102;
  wire popcount40_ghhv_core_104;
  wire popcount40_ghhv_core_107;
  wire popcount40_ghhv_core_108;
  wire popcount40_ghhv_core_109;
  wire popcount40_ghhv_core_112;
  wire popcount40_ghhv_core_115;
  wire popcount40_ghhv_core_119;
  wire popcount40_ghhv_core_120;
  wire popcount40_ghhv_core_123;
  wire popcount40_ghhv_core_124;
  wire popcount40_ghhv_core_125;
  wire popcount40_ghhv_core_127;
  wire popcount40_ghhv_core_128;
  wire popcount40_ghhv_core_130;
  wire popcount40_ghhv_core_131;
  wire popcount40_ghhv_core_133;
  wire popcount40_ghhv_core_134;
  wire popcount40_ghhv_core_135;
  wire popcount40_ghhv_core_138;
  wire popcount40_ghhv_core_139;
  wire popcount40_ghhv_core_140;
  wire popcount40_ghhv_core_143;
  wire popcount40_ghhv_core_145;
  wire popcount40_ghhv_core_146;
  wire popcount40_ghhv_core_147;
  wire popcount40_ghhv_core_148;
  wire popcount40_ghhv_core_150;
  wire popcount40_ghhv_core_151;
  wire popcount40_ghhv_core_152;
  wire popcount40_ghhv_core_157;
  wire popcount40_ghhv_core_158;
  wire popcount40_ghhv_core_159;
  wire popcount40_ghhv_core_160;
  wire popcount40_ghhv_core_161;
  wire popcount40_ghhv_core_162;
  wire popcount40_ghhv_core_163;
  wire popcount40_ghhv_core_164;
  wire popcount40_ghhv_core_165;
  wire popcount40_ghhv_core_166;
  wire popcount40_ghhv_core_167;
  wire popcount40_ghhv_core_169;
  wire popcount40_ghhv_core_170;
  wire popcount40_ghhv_core_171;
  wire popcount40_ghhv_core_172;
  wire popcount40_ghhv_core_173;
  wire popcount40_ghhv_core_175;
  wire popcount40_ghhv_core_177;
  wire popcount40_ghhv_core_178;
  wire popcount40_ghhv_core_180;
  wire popcount40_ghhv_core_182_not;
  wire popcount40_ghhv_core_183;
  wire popcount40_ghhv_core_184;
  wire popcount40_ghhv_core_185;
  wire popcount40_ghhv_core_186;
  wire popcount40_ghhv_core_187;
  wire popcount40_ghhv_core_188;
  wire popcount40_ghhv_core_189;
  wire popcount40_ghhv_core_190;
  wire popcount40_ghhv_core_191;
  wire popcount40_ghhv_core_192;
  wire popcount40_ghhv_core_193;
  wire popcount40_ghhv_core_194_not;
  wire popcount40_ghhv_core_198;
  wire popcount40_ghhv_core_202;
  wire popcount40_ghhv_core_203;
  wire popcount40_ghhv_core_204;
  wire popcount40_ghhv_core_206;
  wire popcount40_ghhv_core_208;
  wire popcount40_ghhv_core_209;
  wire popcount40_ghhv_core_210;
  wire popcount40_ghhv_core_211;
  wire popcount40_ghhv_core_212;
  wire popcount40_ghhv_core_213;
  wire popcount40_ghhv_core_215;
  wire popcount40_ghhv_core_216;
  wire popcount40_ghhv_core_218;
  wire popcount40_ghhv_core_219;
  wire popcount40_ghhv_core_220_not;
  wire popcount40_ghhv_core_222;
  wire popcount40_ghhv_core_224;
  wire popcount40_ghhv_core_225;
  wire popcount40_ghhv_core_226;
  wire popcount40_ghhv_core_228;
  wire popcount40_ghhv_core_229;
  wire popcount40_ghhv_core_230;
  wire popcount40_ghhv_core_231;
  wire popcount40_ghhv_core_232;
  wire popcount40_ghhv_core_234;
  wire popcount40_ghhv_core_235;
  wire popcount40_ghhv_core_236;
  wire popcount40_ghhv_core_237;
  wire popcount40_ghhv_core_239;
  wire popcount40_ghhv_core_244;
  wire popcount40_ghhv_core_246;
  wire popcount40_ghhv_core_247;
  wire popcount40_ghhv_core_248;
  wire popcount40_ghhv_core_249;
  wire popcount40_ghhv_core_250;
  wire popcount40_ghhv_core_251;
  wire popcount40_ghhv_core_252;
  wire popcount40_ghhv_core_253;
  wire popcount40_ghhv_core_255;
  wire popcount40_ghhv_core_256;
  wire popcount40_ghhv_core_257;
  wire popcount40_ghhv_core_258;
  wire popcount40_ghhv_core_260;
  wire popcount40_ghhv_core_261;
  wire popcount40_ghhv_core_262;
  wire popcount40_ghhv_core_263;
  wire popcount40_ghhv_core_269;
  wire popcount40_ghhv_core_271;
  wire popcount40_ghhv_core_272;
  wire popcount40_ghhv_core_273;
  wire popcount40_ghhv_core_275;
  wire popcount40_ghhv_core_276;
  wire popcount40_ghhv_core_277;
  wire popcount40_ghhv_core_280;
  wire popcount40_ghhv_core_283;
  wire popcount40_ghhv_core_284;
  wire popcount40_ghhv_core_285;
  wire popcount40_ghhv_core_287;
  wire popcount40_ghhv_core_288;
  wire popcount40_ghhv_core_291;
  wire popcount40_ghhv_core_294;
  wire popcount40_ghhv_core_296;
  wire popcount40_ghhv_core_297;
  wire popcount40_ghhv_core_299;
  wire popcount40_ghhv_core_300;
  wire popcount40_ghhv_core_306;
  wire popcount40_ghhv_core_307;
  wire popcount40_ghhv_core_310;
  wire popcount40_ghhv_core_311;
  wire popcount40_ghhv_core_313;
  wire popcount40_ghhv_core_315;
  wire popcount40_ghhv_core_316;

  assign popcount40_ghhv_core_042 = input_a[37] ^ input_a[27];
  assign popcount40_ghhv_core_043_not = ~input_a[14];
  assign popcount40_ghhv_core_047 = input_a[25] ^ input_a[16];
  assign popcount40_ghhv_core_048 = input_a[17] | input_a[7];
  assign popcount40_ghhv_core_049 = ~(input_a[31] | input_a[15]);
  assign popcount40_ghhv_core_051 = ~(input_a[8] & input_a[15]);
  assign popcount40_ghhv_core_055 = input_a[14] ^ input_a[0];
  assign popcount40_ghhv_core_056 = input_a[17] | input_a[24];
  assign popcount40_ghhv_core_057 = input_a[28] | input_a[12];
  assign popcount40_ghhv_core_058 = input_a[29] | input_a[13];
  assign popcount40_ghhv_core_059 = ~(input_a[15] & input_a[35]);
  assign popcount40_ghhv_core_061 = input_a[13] & input_a[7];
  assign popcount40_ghhv_core_063 = input_a[12] ^ input_a[20];
  assign popcount40_ghhv_core_064 = ~(input_a[25] ^ input_a[31]);
  assign popcount40_ghhv_core_065 = input_a[35] & input_a[1];
  assign popcount40_ghhv_core_067 = input_a[15] | input_a[25];
  assign popcount40_ghhv_core_069 = ~(input_a[2] & input_a[2]);
  assign popcount40_ghhv_core_070 = input_a[38] | input_a[28];
  assign popcount40_ghhv_core_072 = ~input_a[19];
  assign popcount40_ghhv_core_073 = ~(input_a[10] & input_a[26]);
  assign popcount40_ghhv_core_075 = input_a[39] ^ input_a[36];
  assign popcount40_ghhv_core_076 = input_a[39] ^ input_a[8];
  assign popcount40_ghhv_core_077 = input_a[26] ^ input_a[31];
  assign popcount40_ghhv_core_079 = ~(input_a[2] & input_a[12]);
  assign popcount40_ghhv_core_080 = input_a[0] | input_a[25];
  assign popcount40_ghhv_core_084 = ~input_a[11];
  assign popcount40_ghhv_core_085 = ~(input_a[32] ^ input_a[15]);
  assign popcount40_ghhv_core_086 = ~(input_a[4] | input_a[25]);
  assign popcount40_ghhv_core_088_not = ~input_a[12];
  assign popcount40_ghhv_core_089 = ~(input_a[10] & input_a[31]);
  assign popcount40_ghhv_core_090 = input_a[16] & input_a[34];
  assign popcount40_ghhv_core_092 = ~(input_a[3] & input_a[20]);
  assign popcount40_ghhv_core_093 = input_a[34] ^ input_a[7];
  assign popcount40_ghhv_core_094 = ~(input_a[19] ^ input_a[21]);
  assign popcount40_ghhv_core_098 = ~(input_a[25] | input_a[1]);
  assign popcount40_ghhv_core_099 = ~(input_a[18] & input_a[35]);
  assign popcount40_ghhv_core_100 = ~(input_a[26] ^ input_a[18]);
  assign popcount40_ghhv_core_102 = input_a[32] & input_a[6];
  assign popcount40_ghhv_core_104 = ~(input_a[1] ^ input_a[31]);
  assign popcount40_ghhv_core_107 = input_a[36] ^ input_a[15];
  assign popcount40_ghhv_core_108 = ~(input_a[14] | input_a[5]);
  assign popcount40_ghhv_core_109 = ~input_a[34];
  assign popcount40_ghhv_core_112 = input_a[8] & input_a[13];
  assign popcount40_ghhv_core_115 = ~(input_a[4] ^ input_a[12]);
  assign popcount40_ghhv_core_119 = ~(input_a[39] ^ input_a[26]);
  assign popcount40_ghhv_core_120 = input_a[37] ^ input_a[33];
  assign popcount40_ghhv_core_123 = ~input_a[39];
  assign popcount40_ghhv_core_124 = input_a[14] ^ input_a[36];
  assign popcount40_ghhv_core_125 = input_a[2] | input_a[37];
  assign popcount40_ghhv_core_127 = input_a[1] | input_a[8];
  assign popcount40_ghhv_core_128 = ~(input_a[37] | input_a[39]);
  assign popcount40_ghhv_core_130 = input_a[0] & input_a[13];
  assign popcount40_ghhv_core_131 = input_a[3] ^ input_a[18];
  assign popcount40_ghhv_core_133 = input_a[10] & input_a[3];
  assign popcount40_ghhv_core_134 = input_a[25] | input_a[24];
  assign popcount40_ghhv_core_135 = input_a[9] ^ input_a[17];
  assign popcount40_ghhv_core_138 = ~input_a[32];
  assign popcount40_ghhv_core_139 = ~(input_a[16] & input_a[9]);
  assign popcount40_ghhv_core_140 = input_a[12] | input_a[12];
  assign popcount40_ghhv_core_143 = input_a[33] ^ input_a[21];
  assign popcount40_ghhv_core_145 = ~input_a[36];
  assign popcount40_ghhv_core_146 = ~input_a[7];
  assign popcount40_ghhv_core_147 = input_a[29] | input_a[11];
  assign popcount40_ghhv_core_148 = input_a[15] ^ input_a[29];
  assign popcount40_ghhv_core_150 = ~(input_a[31] | input_a[18]);
  assign popcount40_ghhv_core_151 = ~input_a[24];
  assign popcount40_ghhv_core_152 = ~(input_a[21] ^ input_a[31]);
  assign popcount40_ghhv_core_157 = input_a[27] | input_a[34];
  assign popcount40_ghhv_core_158 = input_a[7] ^ input_a[6];
  assign popcount40_ghhv_core_159 = input_a[19] & input_a[19];
  assign popcount40_ghhv_core_160 = ~(input_a[38] | input_a[27]);
  assign popcount40_ghhv_core_161 = input_a[1] ^ input_a[20];
  assign popcount40_ghhv_core_162 = ~(input_a[37] ^ input_a[27]);
  assign popcount40_ghhv_core_163 = ~(input_a[22] & input_a[35]);
  assign popcount40_ghhv_core_164 = input_a[12] ^ input_a[28];
  assign popcount40_ghhv_core_165 = input_a[18] ^ input_a[18];
  assign popcount40_ghhv_core_166 = input_a[15] ^ input_a[2];
  assign popcount40_ghhv_core_167 = input_a[1] ^ input_a[28];
  assign popcount40_ghhv_core_169 = ~(input_a[14] ^ input_a[36]);
  assign popcount40_ghhv_core_170 = input_a[29] & input_a[20];
  assign popcount40_ghhv_core_171 = input_a[14] | input_a[25];
  assign popcount40_ghhv_core_172 = ~(input_a[35] ^ input_a[9]);
  assign popcount40_ghhv_core_173 = ~input_a[2];
  assign popcount40_ghhv_core_175 = input_a[32] ^ input_a[38];
  assign popcount40_ghhv_core_177 = ~(input_a[3] & input_a[2]);
  assign popcount40_ghhv_core_178 = ~input_a[18];
  assign popcount40_ghhv_core_180 = input_a[17] & input_a[19];
  assign popcount40_ghhv_core_182_not = ~input_a[14];
  assign popcount40_ghhv_core_183 = input_a[34] ^ input_a[2];
  assign popcount40_ghhv_core_184 = ~(input_a[17] ^ input_a[11]);
  assign popcount40_ghhv_core_185 = input_a[4] & input_a[13];
  assign popcount40_ghhv_core_186 = ~(input_a[35] & input_a[22]);
  assign popcount40_ghhv_core_187 = ~(input_a[11] ^ input_a[5]);
  assign popcount40_ghhv_core_188 = ~(input_a[27] | input_a[18]);
  assign popcount40_ghhv_core_189 = ~(input_a[4] | input_a[33]);
  assign popcount40_ghhv_core_190 = input_a[13] & input_a[22];
  assign popcount40_ghhv_core_191 = input_a[19] & input_a[35];
  assign popcount40_ghhv_core_192 = input_a[22] | input_a[27];
  assign popcount40_ghhv_core_193 = ~(input_a[15] ^ input_a[32]);
  assign popcount40_ghhv_core_194_not = ~input_a[39];
  assign popcount40_ghhv_core_198 = input_a[28] ^ input_a[29];
  assign popcount40_ghhv_core_202 = ~(input_a[22] | input_a[13]);
  assign popcount40_ghhv_core_203 = input_a[19] ^ input_a[3];
  assign popcount40_ghhv_core_204 = input_a[20] | input_a[8];
  assign popcount40_ghhv_core_206 = ~(input_a[0] ^ input_a[13]);
  assign popcount40_ghhv_core_208 = ~input_a[39];
  assign popcount40_ghhv_core_209 = ~input_a[2];
  assign popcount40_ghhv_core_210 = input_a[17] & input_a[36];
  assign popcount40_ghhv_core_211 = input_a[24] | input_a[38];
  assign popcount40_ghhv_core_212 = input_a[10] | input_a[14];
  assign popcount40_ghhv_core_213 = input_a[37] & input_a[27];
  assign popcount40_ghhv_core_215 = input_a[8] ^ input_a[33];
  assign popcount40_ghhv_core_216 = input_a[23] | input_a[10];
  assign popcount40_ghhv_core_218 = input_a[16] ^ input_a[30];
  assign popcount40_ghhv_core_219 = ~input_a[21];
  assign popcount40_ghhv_core_220_not = ~input_a[4];
  assign popcount40_ghhv_core_222 = ~(input_a[29] ^ input_a[32]);
  assign popcount40_ghhv_core_224 = input_a[36] ^ input_a[7];
  assign popcount40_ghhv_core_225 = ~(input_a[9] & input_a[16]);
  assign popcount40_ghhv_core_226 = ~(input_a[28] ^ input_a[17]);
  assign popcount40_ghhv_core_228 = ~(input_a[14] & input_a[21]);
  assign popcount40_ghhv_core_229 = input_a[14] ^ input_a[26];
  assign popcount40_ghhv_core_230 = ~(input_a[26] ^ input_a[2]);
  assign popcount40_ghhv_core_231 = ~(input_a[29] ^ input_a[24]);
  assign popcount40_ghhv_core_232 = input_a[36] & input_a[24];
  assign popcount40_ghhv_core_234 = ~(input_a[18] & input_a[9]);
  assign popcount40_ghhv_core_235 = input_a[7] ^ input_a[14];
  assign popcount40_ghhv_core_236 = input_a[24] | input_a[39];
  assign popcount40_ghhv_core_237 = input_a[10] & input_a[16];
  assign popcount40_ghhv_core_239 = ~(input_a[12] | input_a[37]);
  assign popcount40_ghhv_core_244 = input_a[35] | input_a[23];
  assign popcount40_ghhv_core_246 = ~(input_a[3] & input_a[32]);
  assign popcount40_ghhv_core_247 = input_a[3] ^ input_a[29];
  assign popcount40_ghhv_core_248 = ~(input_a[36] | input_a[32]);
  assign popcount40_ghhv_core_249 = ~(input_a[37] | input_a[24]);
  assign popcount40_ghhv_core_250 = ~input_a[18];
  assign popcount40_ghhv_core_251 = ~(input_a[22] | input_a[33]);
  assign popcount40_ghhv_core_252 = ~input_a[2];
  assign popcount40_ghhv_core_253 = input_a[22] ^ input_a[7];
  assign popcount40_ghhv_core_255 = input_a[7] & input_a[6];
  assign popcount40_ghhv_core_256 = input_a[22] & input_a[17];
  assign popcount40_ghhv_core_257 = ~(input_a[33] ^ input_a[12]);
  assign popcount40_ghhv_core_258 = ~(input_a[37] & input_a[36]);
  assign popcount40_ghhv_core_260 = ~(input_a[14] ^ input_a[21]);
  assign popcount40_ghhv_core_261 = ~(input_a[21] ^ input_a[0]);
  assign popcount40_ghhv_core_262 = ~input_a[24];
  assign popcount40_ghhv_core_263 = ~(input_a[32] & input_a[21]);
  assign popcount40_ghhv_core_269 = ~(input_a[2] & input_a[32]);
  assign popcount40_ghhv_core_271 = input_a[2] ^ input_a[22];
  assign popcount40_ghhv_core_272 = ~(input_a[20] & input_a[30]);
  assign popcount40_ghhv_core_273 = ~(input_a[36] | input_a[31]);
  assign popcount40_ghhv_core_275 = ~input_a[35];
  assign popcount40_ghhv_core_276 = ~(input_a[23] ^ input_a[0]);
  assign popcount40_ghhv_core_277 = ~input_a[39];
  assign popcount40_ghhv_core_280 = ~input_a[9];
  assign popcount40_ghhv_core_283 = ~(input_a[26] | input_a[38]);
  assign popcount40_ghhv_core_284 = input_a[30] ^ input_a[23];
  assign popcount40_ghhv_core_285 = input_a[17] & input_a[37];
  assign popcount40_ghhv_core_287 = input_a[32] | input_a[21];
  assign popcount40_ghhv_core_288 = ~(input_a[0] & input_a[4]);
  assign popcount40_ghhv_core_291 = input_a[2] | input_a[3];
  assign popcount40_ghhv_core_294 = input_a[34] | input_a[34];
  assign popcount40_ghhv_core_296 = ~(input_a[25] ^ input_a[10]);
  assign popcount40_ghhv_core_297 = ~input_a[4];
  assign popcount40_ghhv_core_299 = ~input_a[19];
  assign popcount40_ghhv_core_300 = input_a[39] | input_a[14];
  assign popcount40_ghhv_core_306 = ~(input_a[32] ^ input_a[11]);
  assign popcount40_ghhv_core_307 = ~(input_a[16] ^ input_a[33]);
  assign popcount40_ghhv_core_310 = input_a[21] ^ input_a[18];
  assign popcount40_ghhv_core_311 = input_a[22] & input_a[10];
  assign popcount40_ghhv_core_313 = ~(input_a[24] & input_a[37]);
  assign popcount40_ghhv_core_315 = ~(input_a[39] ^ input_a[6]);
  assign popcount40_ghhv_core_316 = input_a[14] | input_a[13];

  assign popcount40_ghhv_out[0] = 1'b0;
  assign popcount40_ghhv_out[1] = 1'b1;
  assign popcount40_ghhv_out[2] = input_a[7];
  assign popcount40_ghhv_out[3] = 1'b1;
  assign popcount40_ghhv_out[4] = input_a[12];
  assign popcount40_ghhv_out[5] = input_a[33];
endmodule