// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.79938
// WCE=19.0
// EP=0.825257%
// Printed PDK parameters:
//  Area=45886051.0
//  Delay=58474496.0
//  Power=2302800.0

module popcount36_bd2s(input [35:0] input_a, output [5:0] popcount36_bd2s_out);
  wire popcount36_bd2s_core_038;
  wire popcount36_bd2s_core_039;
  wire popcount36_bd2s_core_040;
  wire popcount36_bd2s_core_041;
  wire popcount36_bd2s_core_043;
  wire popcount36_bd2s_core_045;
  wire popcount36_bd2s_core_046;
  wire popcount36_bd2s_core_050;
  wire popcount36_bd2s_core_051;
  wire popcount36_bd2s_core_055;
  wire popcount36_bd2s_core_057;
  wire popcount36_bd2s_core_058;
  wire popcount36_bd2s_core_059;
  wire popcount36_bd2s_core_061;
  wire popcount36_bd2s_core_062;
  wire popcount36_bd2s_core_063;
  wire popcount36_bd2s_core_067;
  wire popcount36_bd2s_core_068;
  wire popcount36_bd2s_core_069;
  wire popcount36_bd2s_core_071;
  wire popcount36_bd2s_core_073;
  wire popcount36_bd2s_core_074;
  wire popcount36_bd2s_core_075;
  wire popcount36_bd2s_core_077;
  wire popcount36_bd2s_core_081;
  wire popcount36_bd2s_core_082;
  wire popcount36_bd2s_core_083;
  wire popcount36_bd2s_core_084_not;
  wire popcount36_bd2s_core_086;
  wire popcount36_bd2s_core_088;
  wire popcount36_bd2s_core_089;
  wire popcount36_bd2s_core_091;
  wire popcount36_bd2s_core_092;
  wire popcount36_bd2s_core_093;
  wire popcount36_bd2s_core_094;
  wire popcount36_bd2s_core_095;
  wire popcount36_bd2s_core_096;
  wire popcount36_bd2s_core_097;
  wire popcount36_bd2s_core_099;
  wire popcount36_bd2s_core_101;
  wire popcount36_bd2s_core_102;
  wire popcount36_bd2s_core_103;
  wire popcount36_bd2s_core_105;
  wire popcount36_bd2s_core_109;
  wire popcount36_bd2s_core_110;
  wire popcount36_bd2s_core_111;
  wire popcount36_bd2s_core_115;
  wire popcount36_bd2s_core_116;
  wire popcount36_bd2s_core_117;
  wire popcount36_bd2s_core_118;
  wire popcount36_bd2s_core_119;
  wire popcount36_bd2s_core_121;
  wire popcount36_bd2s_core_123;
  wire popcount36_bd2s_core_125;
  wire popcount36_bd2s_core_127;
  wire popcount36_bd2s_core_128;
  wire popcount36_bd2s_core_129;
  wire popcount36_bd2s_core_132;
  wire popcount36_bd2s_core_135;
  wire popcount36_bd2s_core_136;
  wire popcount36_bd2s_core_137;
  wire popcount36_bd2s_core_138;
  wire popcount36_bd2s_core_140;
  wire popcount36_bd2s_core_144;
  wire popcount36_bd2s_core_145;
  wire popcount36_bd2s_core_146;
  wire popcount36_bd2s_core_147;
  wire popcount36_bd2s_core_148;
  wire popcount36_bd2s_core_150;
  wire popcount36_bd2s_core_151;
  wire popcount36_bd2s_core_152;
  wire popcount36_bd2s_core_156;
  wire popcount36_bd2s_core_158;
  wire popcount36_bd2s_core_160;
  wire popcount36_bd2s_core_161;
  wire popcount36_bd2s_core_163;
  wire popcount36_bd2s_core_164;
  wire popcount36_bd2s_core_165;
  wire popcount36_bd2s_core_166;
  wire popcount36_bd2s_core_167;
  wire popcount36_bd2s_core_168;
  wire popcount36_bd2s_core_169;
  wire popcount36_bd2s_core_172;
  wire popcount36_bd2s_core_173;
  wire popcount36_bd2s_core_174;
  wire popcount36_bd2s_core_175;
  wire popcount36_bd2s_core_179;
  wire popcount36_bd2s_core_180;
  wire popcount36_bd2s_core_181;
  wire popcount36_bd2s_core_182;
  wire popcount36_bd2s_core_183;
  wire popcount36_bd2s_core_185;
  wire popcount36_bd2s_core_186;
  wire popcount36_bd2s_core_187;
  wire popcount36_bd2s_core_188;
  wire popcount36_bd2s_core_190;
  wire popcount36_bd2s_core_192;
  wire popcount36_bd2s_core_193;
  wire popcount36_bd2s_core_194;
  wire popcount36_bd2s_core_197;
  wire popcount36_bd2s_core_198;
  wire popcount36_bd2s_core_199;
  wire popcount36_bd2s_core_200;
  wire popcount36_bd2s_core_201;
  wire popcount36_bd2s_core_202;
  wire popcount36_bd2s_core_203;
  wire popcount36_bd2s_core_207;
  wire popcount36_bd2s_core_208;
  wire popcount36_bd2s_core_209;
  wire popcount36_bd2s_core_210;
  wire popcount36_bd2s_core_211;
  wire popcount36_bd2s_core_214;
  wire popcount36_bd2s_core_215;
  wire popcount36_bd2s_core_216;
  wire popcount36_bd2s_core_217;
  wire popcount36_bd2s_core_223;
  wire popcount36_bd2s_core_226;
  wire popcount36_bd2s_core_227;
  wire popcount36_bd2s_core_228;
  wire popcount36_bd2s_core_229;
  wire popcount36_bd2s_core_230;
  wire popcount36_bd2s_core_231;
  wire popcount36_bd2s_core_233;
  wire popcount36_bd2s_core_235;
  wire popcount36_bd2s_core_236;
  wire popcount36_bd2s_core_237;
  wire popcount36_bd2s_core_238;
  wire popcount36_bd2s_core_239;
  wire popcount36_bd2s_core_242;
  wire popcount36_bd2s_core_246;
  wire popcount36_bd2s_core_248;
  wire popcount36_bd2s_core_249;
  wire popcount36_bd2s_core_252;
  wire popcount36_bd2s_core_253;
  wire popcount36_bd2s_core_254;
  wire popcount36_bd2s_core_255;
  wire popcount36_bd2s_core_256;
  wire popcount36_bd2s_core_257;
  wire popcount36_bd2s_core_258;
  wire popcount36_bd2s_core_259;
  wire popcount36_bd2s_core_260;
  wire popcount36_bd2s_core_261;
  wire popcount36_bd2s_core_262;
  wire popcount36_bd2s_core_263;
  wire popcount36_bd2s_core_264;
  wire popcount36_bd2s_core_265;
  wire popcount36_bd2s_core_266;
  wire popcount36_bd2s_core_268;
  wire popcount36_bd2s_core_269;
  wire popcount36_bd2s_core_273;

  assign popcount36_bd2s_core_038 = ~input_a[4];
  assign popcount36_bd2s_core_039 = input_a[0] & input_a[28];
  assign popcount36_bd2s_core_040 = ~(input_a[4] & input_a[18]);
  assign popcount36_bd2s_core_041 = ~(input_a[24] ^ input_a[35]);
  assign popcount36_bd2s_core_043 = input_a[10] & input_a[2];
  assign popcount36_bd2s_core_045 = input_a[1] & input_a[3];
  assign popcount36_bd2s_core_046 = popcount36_bd2s_core_039 | popcount36_bd2s_core_043;
  assign popcount36_bd2s_core_050 = input_a[4] & input_a[5];
  assign popcount36_bd2s_core_051 = input_a[9] ^ input_a[30];
  assign popcount36_bd2s_core_055 = ~input_a[25];
  assign popcount36_bd2s_core_057 = ~input_a[8];
  assign popcount36_bd2s_core_058 = input_a[27] & input_a[6];
  assign popcount36_bd2s_core_059 = input_a[1] | input_a[3];
  assign popcount36_bd2s_core_061 = popcount36_bd2s_core_059 | input_a[6];
  assign popcount36_bd2s_core_062 = popcount36_bd2s_core_059 & popcount36_bd2s_core_058;
  assign popcount36_bd2s_core_063 = popcount36_bd2s_core_050 | popcount36_bd2s_core_062;
  assign popcount36_bd2s_core_067 = input_a[12] ^ input_a[26];
  assign popcount36_bd2s_core_068 = ~input_a[30];
  assign popcount36_bd2s_core_069 = popcount36_bd2s_core_046 & popcount36_bd2s_core_061;
  assign popcount36_bd2s_core_071 = input_a[17] | input_a[32];
  assign popcount36_bd2s_core_073 = popcount36_bd2s_core_045 | popcount36_bd2s_core_063;
  assign popcount36_bd2s_core_074 = ~(input_a[30] ^ input_a[8]);
  assign popcount36_bd2s_core_075 = popcount36_bd2s_core_073 | popcount36_bd2s_core_069;
  assign popcount36_bd2s_core_077 = ~(input_a[19] & input_a[15]);
  assign popcount36_bd2s_core_081 = input_a[9] & input_a[7];
  assign popcount36_bd2s_core_082 = ~(input_a[11] & input_a[12]);
  assign popcount36_bd2s_core_083 = input_a[11] & input_a[12];
  assign popcount36_bd2s_core_084_not = ~popcount36_bd2s_core_082;
  assign popcount36_bd2s_core_086 = popcount36_bd2s_core_081 ^ popcount36_bd2s_core_083;
  assign popcount36_bd2s_core_088 = popcount36_bd2s_core_086 ^ popcount36_bd2s_core_082;
  assign popcount36_bd2s_core_089 = ~(input_a[30] & input_a[12]);
  assign popcount36_bd2s_core_091 = ~input_a[6];
  assign popcount36_bd2s_core_092 = input_a[13] & input_a[14];
  assign popcount36_bd2s_core_093 = ~input_a[9];
  assign popcount36_bd2s_core_094 = input_a[16] & input_a[17];
  assign popcount36_bd2s_core_095 = ~(input_a[13] | input_a[7]);
  assign popcount36_bd2s_core_096 = input_a[15] & input_a[29];
  assign popcount36_bd2s_core_097 = popcount36_bd2s_core_094 | popcount36_bd2s_core_096;
  assign popcount36_bd2s_core_099 = ~(input_a[29] | input_a[30]);
  assign popcount36_bd2s_core_101 = popcount36_bd2s_core_092 ^ popcount36_bd2s_core_097;
  assign popcount36_bd2s_core_102 = input_a[13] & popcount36_bd2s_core_097;
  assign popcount36_bd2s_core_103 = ~popcount36_bd2s_core_101;
  assign popcount36_bd2s_core_105 = popcount36_bd2s_core_102 | popcount36_bd2s_core_101;
  assign popcount36_bd2s_core_109 = input_a[34] ^ input_a[18];
  assign popcount36_bd2s_core_110 = popcount36_bd2s_core_088 ^ popcount36_bd2s_core_103;
  assign popcount36_bd2s_core_111 = popcount36_bd2s_core_088 & popcount36_bd2s_core_103;
  assign popcount36_bd2s_core_115 = popcount36_bd2s_core_081 ^ popcount36_bd2s_core_105;
  assign popcount36_bd2s_core_116 = popcount36_bd2s_core_081 & popcount36_bd2s_core_105;
  assign popcount36_bd2s_core_117 = popcount36_bd2s_core_115 ^ popcount36_bd2s_core_111;
  assign popcount36_bd2s_core_118 = popcount36_bd2s_core_115 & popcount36_bd2s_core_111;
  assign popcount36_bd2s_core_119 = popcount36_bd2s_core_116 | popcount36_bd2s_core_118;
  assign popcount36_bd2s_core_121 = input_a[35] | input_a[8];
  assign popcount36_bd2s_core_123 = input_a[6] | input_a[23];
  assign popcount36_bd2s_core_125 = input_a[21] ^ input_a[4];
  assign popcount36_bd2s_core_127 = input_a[17] ^ input_a[8];
  assign popcount36_bd2s_core_128 = input_a[0] ^ input_a[35];
  assign popcount36_bd2s_core_129 = popcount36_bd2s_core_075 ^ popcount36_bd2s_core_117;
  assign popcount36_bd2s_core_132 = input_a[31] & input_a[16];
  assign popcount36_bd2s_core_135 = ~input_a[3];
  assign popcount36_bd2s_core_136 = popcount36_bd2s_core_119 | popcount36_bd2s_core_075;
  assign popcount36_bd2s_core_137 = ~(input_a[15] | input_a[25]);
  assign popcount36_bd2s_core_138 = input_a[20] & input_a[6];
  assign popcount36_bd2s_core_140 = ~input_a[13];
  assign popcount36_bd2s_core_144 = input_a[18] ^ input_a[19];
  assign popcount36_bd2s_core_145 = input_a[18] & input_a[19];
  assign popcount36_bd2s_core_146 = input_a[8] & input_a[29];
  assign popcount36_bd2s_core_147 = input_a[20] & input_a[24];
  assign popcount36_bd2s_core_148 = input_a[11] | input_a[35];
  assign popcount36_bd2s_core_150 = input_a[19] ^ popcount36_bd2s_core_147;
  assign popcount36_bd2s_core_151 = popcount36_bd2s_core_145 & popcount36_bd2s_core_147;
  assign popcount36_bd2s_core_152 = popcount36_bd2s_core_150 | popcount36_bd2s_core_144;
  assign popcount36_bd2s_core_156 = input_a[22] & input_a[23];
  assign popcount36_bd2s_core_158 = input_a[25] & input_a[26];
  assign popcount36_bd2s_core_160 = input_a[21] & input_a[30];
  assign popcount36_bd2s_core_161 = popcount36_bd2s_core_158 | popcount36_bd2s_core_160;
  assign popcount36_bd2s_core_163 = ~input_a[21];
  assign popcount36_bd2s_core_164 = input_a[19] ^ input_a[4];
  assign popcount36_bd2s_core_165 = popcount36_bd2s_core_156 ^ popcount36_bd2s_core_161;
  assign popcount36_bd2s_core_166 = popcount36_bd2s_core_156 & popcount36_bd2s_core_161;
  assign popcount36_bd2s_core_167 = popcount36_bd2s_core_165 ^ input_a[8];
  assign popcount36_bd2s_core_168 = popcount36_bd2s_core_165 & input_a[8];
  assign popcount36_bd2s_core_169 = popcount36_bd2s_core_166 | popcount36_bd2s_core_168;
  assign popcount36_bd2s_core_172 = ~(input_a[27] & input_a[33]);
  assign popcount36_bd2s_core_173 = ~(input_a[1] & input_a[18]);
  assign popcount36_bd2s_core_174 = popcount36_bd2s_core_152 ^ popcount36_bd2s_core_167;
  assign popcount36_bd2s_core_175 = popcount36_bd2s_core_152 & popcount36_bd2s_core_167;
  assign popcount36_bd2s_core_179 = popcount36_bd2s_core_151 ^ popcount36_bd2s_core_169;
  assign popcount36_bd2s_core_180 = popcount36_bd2s_core_151 & popcount36_bd2s_core_169;
  assign popcount36_bd2s_core_181 = popcount36_bd2s_core_179 ^ popcount36_bd2s_core_175;
  assign popcount36_bd2s_core_182 = popcount36_bd2s_core_179 & popcount36_bd2s_core_175;
  assign popcount36_bd2s_core_183 = popcount36_bd2s_core_180 | popcount36_bd2s_core_182;
  assign popcount36_bd2s_core_185 = ~input_a[21];
  assign popcount36_bd2s_core_186 = input_a[24] | input_a[2];
  assign popcount36_bd2s_core_187 = input_a[30] ^ input_a[33];
  assign popcount36_bd2s_core_188 = ~(input_a[20] | input_a[10]);
  assign popcount36_bd2s_core_190 = input_a[17] & input_a[23];
  assign popcount36_bd2s_core_192 = ~(input_a[10] & input_a[30]);
  assign popcount36_bd2s_core_193 = ~(input_a[14] | input_a[10]);
  assign popcount36_bd2s_core_194 = input_a[10] | popcount36_bd2s_core_186;
  assign popcount36_bd2s_core_197 = input_a[31] ^ input_a[32];
  assign popcount36_bd2s_core_198 = input_a[31] & input_a[32];
  assign popcount36_bd2s_core_199 = input_a[34] | input_a[35];
  assign popcount36_bd2s_core_200 = input_a[34] & input_a[35];
  assign popcount36_bd2s_core_201 = ~(input_a[3] ^ input_a[23]);
  assign popcount36_bd2s_core_202 = input_a[33] & popcount36_bd2s_core_199;
  assign popcount36_bd2s_core_203 = popcount36_bd2s_core_200 | popcount36_bd2s_core_202;
  assign popcount36_bd2s_core_207 = popcount36_bd2s_core_198 ^ popcount36_bd2s_core_203;
  assign popcount36_bd2s_core_208 = input_a[31] & popcount36_bd2s_core_203;
  assign popcount36_bd2s_core_209 = popcount36_bd2s_core_207 ^ popcount36_bd2s_core_197;
  assign popcount36_bd2s_core_210 = popcount36_bd2s_core_207 & popcount36_bd2s_core_197;
  assign popcount36_bd2s_core_211 = popcount36_bd2s_core_208 | popcount36_bd2s_core_210;
  assign popcount36_bd2s_core_214 = ~input_a[32];
  assign popcount36_bd2s_core_215 = ~input_a[12];
  assign popcount36_bd2s_core_216 = popcount36_bd2s_core_194 ^ popcount36_bd2s_core_209;
  assign popcount36_bd2s_core_217 = popcount36_bd2s_core_194 & popcount36_bd2s_core_209;
  assign popcount36_bd2s_core_223 = popcount36_bd2s_core_211 | popcount36_bd2s_core_217;
  assign popcount36_bd2s_core_226 = input_a[12] | input_a[24];
  assign popcount36_bd2s_core_227 = ~(input_a[10] | input_a[22]);
  assign popcount36_bd2s_core_228 = ~(input_a[27] & input_a[14]);
  assign popcount36_bd2s_core_229 = ~input_a[0];
  assign popcount36_bd2s_core_230 = popcount36_bd2s_core_174 ^ popcount36_bd2s_core_216;
  assign popcount36_bd2s_core_231 = popcount36_bd2s_core_174 & popcount36_bd2s_core_216;
  assign popcount36_bd2s_core_233 = ~(input_a[20] ^ input_a[19]);
  assign popcount36_bd2s_core_235 = ~(popcount36_bd2s_core_181 & popcount36_bd2s_core_223);
  assign popcount36_bd2s_core_236 = popcount36_bd2s_core_181 & popcount36_bd2s_core_223;
  assign popcount36_bd2s_core_237 = popcount36_bd2s_core_235 ^ popcount36_bd2s_core_231;
  assign popcount36_bd2s_core_238 = popcount36_bd2s_core_235 & popcount36_bd2s_core_231;
  assign popcount36_bd2s_core_239 = popcount36_bd2s_core_236 | popcount36_bd2s_core_238;
  assign popcount36_bd2s_core_242 = popcount36_bd2s_core_183 ^ popcount36_bd2s_core_239;
  assign popcount36_bd2s_core_246 = ~input_a[0];
  assign popcount36_bd2s_core_248 = ~input_a[13];
  assign popcount36_bd2s_core_249 = ~(input_a[1] ^ input_a[20]);
  assign popcount36_bd2s_core_252 = popcount36_bd2s_core_110 ^ popcount36_bd2s_core_230;
  assign popcount36_bd2s_core_253 = popcount36_bd2s_core_110 & popcount36_bd2s_core_230;
  assign popcount36_bd2s_core_254 = popcount36_bd2s_core_252 ^ popcount36_bd2s_core_084_not;
  assign popcount36_bd2s_core_255 = popcount36_bd2s_core_252 & popcount36_bd2s_core_084_not;
  assign popcount36_bd2s_core_256 = popcount36_bd2s_core_253 | popcount36_bd2s_core_255;
  assign popcount36_bd2s_core_257 = popcount36_bd2s_core_129 ^ popcount36_bd2s_core_237;
  assign popcount36_bd2s_core_258 = popcount36_bd2s_core_129 & popcount36_bd2s_core_237;
  assign popcount36_bd2s_core_259 = popcount36_bd2s_core_257 ^ popcount36_bd2s_core_256;
  assign popcount36_bd2s_core_260 = popcount36_bd2s_core_257 & popcount36_bd2s_core_256;
  assign popcount36_bd2s_core_261 = popcount36_bd2s_core_258 | popcount36_bd2s_core_260;
  assign popcount36_bd2s_core_262 = popcount36_bd2s_core_136 ^ popcount36_bd2s_core_242;
  assign popcount36_bd2s_core_263 = popcount36_bd2s_core_136 & popcount36_bd2s_core_242;
  assign popcount36_bd2s_core_264 = popcount36_bd2s_core_262 ^ popcount36_bd2s_core_261;
  assign popcount36_bd2s_core_265 = popcount36_bd2s_core_262 & popcount36_bd2s_core_261;
  assign popcount36_bd2s_core_266 = popcount36_bd2s_core_263 | popcount36_bd2s_core_265;
  assign popcount36_bd2s_core_268 = ~(input_a[3] | input_a[27]);
  assign popcount36_bd2s_core_269 = popcount36_bd2s_core_183 | popcount36_bd2s_core_266;
  assign popcount36_bd2s_core_273 = input_a[9] ^ input_a[31];

  assign popcount36_bd2s_out[0] = popcount36_bd2s_core_262;
  assign popcount36_bd2s_out[1] = popcount36_bd2s_core_254;
  assign popcount36_bd2s_out[2] = popcount36_bd2s_core_259;
  assign popcount36_bd2s_out[3] = popcount36_bd2s_core_264;
  assign popcount36_bd2s_out[4] = popcount36_bd2s_core_269;
  assign popcount36_bd2s_out[5] = 1'b0;
endmodule