// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.93416
// WCE=12.0
// EP=0.83882%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_9965(input [23:0] input_a, output [4:0] popcount24_9965_out);
  wire popcount24_9965_core_027;
  wire popcount24_9965_core_028;
  wire popcount24_9965_core_029_not;
  wire popcount24_9965_core_030;
  wire popcount24_9965_core_031;
  wire popcount24_9965_core_033;
  wire popcount24_9965_core_038;
  wire popcount24_9965_core_039;
  wire popcount24_9965_core_041;
  wire popcount24_9965_core_042;
  wire popcount24_9965_core_043;
  wire popcount24_9965_core_045;
  wire popcount24_9965_core_047;
  wire popcount24_9965_core_050;
  wire popcount24_9965_core_051;
  wire popcount24_9965_core_053;
  wire popcount24_9965_core_054;
  wire popcount24_9965_core_055;
  wire popcount24_9965_core_056;
  wire popcount24_9965_core_061;
  wire popcount24_9965_core_064;
  wire popcount24_9965_core_067;
  wire popcount24_9965_core_070;
  wire popcount24_9965_core_071;
  wire popcount24_9965_core_072;
  wire popcount24_9965_core_073;
  wire popcount24_9965_core_075;
  wire popcount24_9965_core_079;
  wire popcount24_9965_core_082;
  wire popcount24_9965_core_083;
  wire popcount24_9965_core_086;
  wire popcount24_9965_core_089;
  wire popcount24_9965_core_090;
  wire popcount24_9965_core_091;
  wire popcount24_9965_core_093_not;
  wire popcount24_9965_core_096;
  wire popcount24_9965_core_098;
  wire popcount24_9965_core_100_not;
  wire popcount24_9965_core_101;
  wire popcount24_9965_core_102;
  wire popcount24_9965_core_103;
  wire popcount24_9965_core_104;
  wire popcount24_9965_core_105;
  wire popcount24_9965_core_106;
  wire popcount24_9965_core_108;
  wire popcount24_9965_core_109;
  wire popcount24_9965_core_110;
  wire popcount24_9965_core_112;
  wire popcount24_9965_core_113;
  wire popcount24_9965_core_114;
  wire popcount24_9965_core_117;
  wire popcount24_9965_core_118_not;
  wire popcount24_9965_core_119;
  wire popcount24_9965_core_121;
  wire popcount24_9965_core_123;
  wire popcount24_9965_core_125;
  wire popcount24_9965_core_126;
  wire popcount24_9965_core_127;
  wire popcount24_9965_core_128;
  wire popcount24_9965_core_129;
  wire popcount24_9965_core_130;
  wire popcount24_9965_core_131;
  wire popcount24_9965_core_133;
  wire popcount24_9965_core_134;
  wire popcount24_9965_core_137;
  wire popcount24_9965_core_141;
  wire popcount24_9965_core_143;
  wire popcount24_9965_core_146;
  wire popcount24_9965_core_147;
  wire popcount24_9965_core_151;
  wire popcount24_9965_core_153;
  wire popcount24_9965_core_156;
  wire popcount24_9965_core_157;
  wire popcount24_9965_core_158;
  wire popcount24_9965_core_159;
  wire popcount24_9965_core_160;
  wire popcount24_9965_core_161;
  wire popcount24_9965_core_162;
  wire popcount24_9965_core_163;
  wire popcount24_9965_core_165;
  wire popcount24_9965_core_166;
  wire popcount24_9965_core_167;
  wire popcount24_9965_core_168;
  wire popcount24_9965_core_169;
  wire popcount24_9965_core_170;
  wire popcount24_9965_core_171;
  wire popcount24_9965_core_172;
  wire popcount24_9965_core_176;
  wire popcount24_9965_core_177;

  assign popcount24_9965_core_027 = ~input_a[4];
  assign popcount24_9965_core_028 = ~(input_a[23] ^ input_a[2]);
  assign popcount24_9965_core_029_not = ~input_a[3];
  assign popcount24_9965_core_030 = ~(input_a[18] ^ input_a[21]);
  assign popcount24_9965_core_031 = ~input_a[14];
  assign popcount24_9965_core_033 = ~(input_a[0] | input_a[13]);
  assign popcount24_9965_core_038 = input_a[11] ^ input_a[13];
  assign popcount24_9965_core_039 = ~input_a[0];
  assign popcount24_9965_core_041 = ~(input_a[7] & input_a[6]);
  assign popcount24_9965_core_042 = ~(input_a[8] | input_a[9]);
  assign popcount24_9965_core_043 = input_a[2] | input_a[10];
  assign popcount24_9965_core_045 = input_a[5] ^ input_a[21];
  assign popcount24_9965_core_047 = ~input_a[21];
  assign popcount24_9965_core_050 = input_a[22] & input_a[16];
  assign popcount24_9965_core_051 = input_a[5] ^ input_a[1];
  assign popcount24_9965_core_053 = input_a[13] ^ input_a[13];
  assign popcount24_9965_core_054 = input_a[23] | input_a[15];
  assign popcount24_9965_core_055 = input_a[23] & input_a[5];
  assign popcount24_9965_core_056 = ~(input_a[4] & input_a[13]);
  assign popcount24_9965_core_061 = ~(input_a[13] & input_a[2]);
  assign popcount24_9965_core_064 = input_a[15] ^ input_a[18];
  assign popcount24_9965_core_067 = ~input_a[2];
  assign popcount24_9965_core_070 = ~(input_a[12] & input_a[5]);
  assign popcount24_9965_core_071 = input_a[18] | input_a[5];
  assign popcount24_9965_core_072 = input_a[7] | input_a[0];
  assign popcount24_9965_core_073 = ~input_a[22];
  assign popcount24_9965_core_075 = ~input_a[10];
  assign popcount24_9965_core_079 = ~(input_a[20] ^ input_a[9]);
  assign popcount24_9965_core_082 = input_a[21] | input_a[16];
  assign popcount24_9965_core_083 = input_a[23] & input_a[11];
  assign popcount24_9965_core_086 = ~(input_a[16] | input_a[13]);
  assign popcount24_9965_core_089 = input_a[11] | input_a[14];
  assign popcount24_9965_core_090 = input_a[12] ^ input_a[8];
  assign popcount24_9965_core_091 = input_a[17] & input_a[4];
  assign popcount24_9965_core_093_not = ~input_a[20];
  assign popcount24_9965_core_096 = ~(input_a[6] | input_a[18]);
  assign popcount24_9965_core_098 = input_a[7] | input_a[16];
  assign popcount24_9965_core_100_not = ~input_a[13];
  assign popcount24_9965_core_101 = input_a[9] | input_a[5];
  assign popcount24_9965_core_102 = ~(input_a[11] ^ input_a[8]);
  assign popcount24_9965_core_103 = ~(input_a[0] & input_a[13]);
  assign popcount24_9965_core_104 = ~input_a[21];
  assign popcount24_9965_core_105 = input_a[16] & input_a[10];
  assign popcount24_9965_core_106 = ~(input_a[12] | input_a[5]);
  assign popcount24_9965_core_108 = ~(input_a[11] & input_a[3]);
  assign popcount24_9965_core_109 = ~(input_a[16] & input_a[9]);
  assign popcount24_9965_core_110 = ~input_a[22];
  assign popcount24_9965_core_112 = ~(input_a[9] & input_a[15]);
  assign popcount24_9965_core_113 = ~(input_a[16] & input_a[2]);
  assign popcount24_9965_core_114 = ~(input_a[18] ^ input_a[0]);
  assign popcount24_9965_core_117 = ~(input_a[13] | input_a[22]);
  assign popcount24_9965_core_118_not = ~input_a[0];
  assign popcount24_9965_core_119 = input_a[16] & input_a[23];
  assign popcount24_9965_core_121 = input_a[13] & input_a[18];
  assign popcount24_9965_core_123 = ~(input_a[4] ^ input_a[9]);
  assign popcount24_9965_core_125 = input_a[19] & input_a[3];
  assign popcount24_9965_core_126 = ~(input_a[8] & input_a[21]);
  assign popcount24_9965_core_127 = ~(input_a[8] | input_a[10]);
  assign popcount24_9965_core_128 = input_a[12] | input_a[9];
  assign popcount24_9965_core_129 = ~(input_a[11] | input_a[18]);
  assign popcount24_9965_core_130 = ~(input_a[0] ^ input_a[1]);
  assign popcount24_9965_core_131 = ~(input_a[16] & input_a[20]);
  assign popcount24_9965_core_133 = ~(input_a[9] | input_a[0]);
  assign popcount24_9965_core_134 = ~(input_a[3] ^ input_a[16]);
  assign popcount24_9965_core_137 = ~(input_a[9] | input_a[8]);
  assign popcount24_9965_core_141 = input_a[13] ^ input_a[21];
  assign popcount24_9965_core_143 = ~input_a[9];
  assign popcount24_9965_core_146 = input_a[8] & input_a[7];
  assign popcount24_9965_core_147 = ~(input_a[8] & input_a[9]);
  assign popcount24_9965_core_151 = ~(input_a[5] | input_a[1]);
  assign popcount24_9965_core_153 = ~(input_a[15] & input_a[22]);
  assign popcount24_9965_core_156 = ~input_a[4];
  assign popcount24_9965_core_157 = ~(input_a[2] | input_a[13]);
  assign popcount24_9965_core_158 = input_a[6] & input_a[18];
  assign popcount24_9965_core_159 = input_a[1] & input_a[20];
  assign popcount24_9965_core_160 = ~(input_a[22] ^ input_a[10]);
  assign popcount24_9965_core_161 = ~input_a[14];
  assign popcount24_9965_core_162 = input_a[5] ^ input_a[15];
  assign popcount24_9965_core_163 = ~(input_a[22] | input_a[18]);
  assign popcount24_9965_core_165 = ~(input_a[11] ^ input_a[12]);
  assign popcount24_9965_core_166 = input_a[10] | input_a[19];
  assign popcount24_9965_core_167 = ~(input_a[12] & input_a[11]);
  assign popcount24_9965_core_168 = input_a[21] ^ input_a[17];
  assign popcount24_9965_core_169 = ~(input_a[6] | input_a[17]);
  assign popcount24_9965_core_170 = input_a[22] ^ input_a[17];
  assign popcount24_9965_core_171 = ~(input_a[4] ^ input_a[16]);
  assign popcount24_9965_core_172 = input_a[14] | input_a[2];
  assign popcount24_9965_core_176 = input_a[21] & input_a[6];
  assign popcount24_9965_core_177 = ~(input_a[6] & input_a[11]);

  assign popcount24_9965_out[0] = 1'b0;
  assign popcount24_9965_out[1] = 1'b0;
  assign popcount24_9965_out[2] = 1'b1;
  assign popcount24_9965_out[3] = 1'b1;
  assign popcount24_9965_out[4] = 1'b0;
endmodule