// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.44575
// WCE=22.0
// EP=0.934939%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_hc56(input [28:0] input_a, output [4:0] popcount29_hc56_out);
  wire popcount29_hc56_core_032;
  wire popcount29_hc56_core_034;
  wire popcount29_hc56_core_036;
  wire popcount29_hc56_core_038;
  wire popcount29_hc56_core_039_not;
  wire popcount29_hc56_core_042;
  wire popcount29_hc56_core_044;
  wire popcount29_hc56_core_045;
  wire popcount29_hc56_core_046;
  wire popcount29_hc56_core_048;
  wire popcount29_hc56_core_049;
  wire popcount29_hc56_core_051;
  wire popcount29_hc56_core_052;
  wire popcount29_hc56_core_054;
  wire popcount29_hc56_core_055;
  wire popcount29_hc56_core_056;
  wire popcount29_hc56_core_057;
  wire popcount29_hc56_core_058;
  wire popcount29_hc56_core_059;
  wire popcount29_hc56_core_063;
  wire popcount29_hc56_core_067;
  wire popcount29_hc56_core_068;
  wire popcount29_hc56_core_069;
  wire popcount29_hc56_core_070;
  wire popcount29_hc56_core_072;
  wire popcount29_hc56_core_073;
  wire popcount29_hc56_core_074;
  wire popcount29_hc56_core_076;
  wire popcount29_hc56_core_078;
  wire popcount29_hc56_core_080;
  wire popcount29_hc56_core_082;
  wire popcount29_hc56_core_086;
  wire popcount29_hc56_core_087;
  wire popcount29_hc56_core_088;
  wire popcount29_hc56_core_089;
  wire popcount29_hc56_core_090;
  wire popcount29_hc56_core_091;
  wire popcount29_hc56_core_092;
  wire popcount29_hc56_core_094;
  wire popcount29_hc56_core_095;
  wire popcount29_hc56_core_096;
  wire popcount29_hc56_core_097;
  wire popcount29_hc56_core_099;
  wire popcount29_hc56_core_100;
  wire popcount29_hc56_core_102;
  wire popcount29_hc56_core_103;
  wire popcount29_hc56_core_104;
  wire popcount29_hc56_core_107;
  wire popcount29_hc56_core_108;
  wire popcount29_hc56_core_109;
  wire popcount29_hc56_core_111;
  wire popcount29_hc56_core_112;
  wire popcount29_hc56_core_113;
  wire popcount29_hc56_core_114;
  wire popcount29_hc56_core_115;
  wire popcount29_hc56_core_117;
  wire popcount29_hc56_core_118;
  wire popcount29_hc56_core_119;
  wire popcount29_hc56_core_121;
  wire popcount29_hc56_core_122;
  wire popcount29_hc56_core_123;
  wire popcount29_hc56_core_124;
  wire popcount29_hc56_core_125;
  wire popcount29_hc56_core_126;
  wire popcount29_hc56_core_127;
  wire popcount29_hc56_core_128;
  wire popcount29_hc56_core_130;
  wire popcount29_hc56_core_131;
  wire popcount29_hc56_core_132;
  wire popcount29_hc56_core_133;
  wire popcount29_hc56_core_134;
  wire popcount29_hc56_core_135;
  wire popcount29_hc56_core_138;
  wire popcount29_hc56_core_139;
  wire popcount29_hc56_core_140;
  wire popcount29_hc56_core_144;
  wire popcount29_hc56_core_146;
  wire popcount29_hc56_core_147;
  wire popcount29_hc56_core_148;
  wire popcount29_hc56_core_149;
  wire popcount29_hc56_core_150;
  wire popcount29_hc56_core_151;
  wire popcount29_hc56_core_152;
  wire popcount29_hc56_core_154;
  wire popcount29_hc56_core_156;
  wire popcount29_hc56_core_157;
  wire popcount29_hc56_core_158;
  wire popcount29_hc56_core_159;
  wire popcount29_hc56_core_161;
  wire popcount29_hc56_core_162;
  wire popcount29_hc56_core_163_not;
  wire popcount29_hc56_core_165;
  wire popcount29_hc56_core_166;
  wire popcount29_hc56_core_168;
  wire popcount29_hc56_core_169;
  wire popcount29_hc56_core_172;
  wire popcount29_hc56_core_173;
  wire popcount29_hc56_core_174;
  wire popcount29_hc56_core_175;
  wire popcount29_hc56_core_176;
  wire popcount29_hc56_core_178_not;
  wire popcount29_hc56_core_179;
  wire popcount29_hc56_core_180;
  wire popcount29_hc56_core_183;
  wire popcount29_hc56_core_186;
  wire popcount29_hc56_core_187_not;
  wire popcount29_hc56_core_188;
  wire popcount29_hc56_core_191;
  wire popcount29_hc56_core_192;
  wire popcount29_hc56_core_194;
  wire popcount29_hc56_core_195;
  wire popcount29_hc56_core_196;
  wire popcount29_hc56_core_197;
  wire popcount29_hc56_core_198;
  wire popcount29_hc56_core_199;
  wire popcount29_hc56_core_201;
  wire popcount29_hc56_core_203;
  wire popcount29_hc56_core_204;
  wire popcount29_hc56_core_205;
  wire popcount29_hc56_core_206;
  wire popcount29_hc56_core_207;

  assign popcount29_hc56_core_032 = ~(input_a[21] | input_a[10]);
  assign popcount29_hc56_core_034 = ~(input_a[8] & input_a[0]);
  assign popcount29_hc56_core_036 = input_a[9] ^ input_a[18];
  assign popcount29_hc56_core_038 = ~(input_a[1] | input_a[9]);
  assign popcount29_hc56_core_039_not = ~input_a[8];
  assign popcount29_hc56_core_042 = ~input_a[20];
  assign popcount29_hc56_core_044 = input_a[16] & input_a[10];
  assign popcount29_hc56_core_045 = ~input_a[10];
  assign popcount29_hc56_core_046 = ~(input_a[28] | input_a[17]);
  assign popcount29_hc56_core_048 = ~(input_a[6] | input_a[13]);
  assign popcount29_hc56_core_049 = ~(input_a[6] & input_a[13]);
  assign popcount29_hc56_core_051 = ~(input_a[0] | input_a[26]);
  assign popcount29_hc56_core_052 = ~input_a[4];
  assign popcount29_hc56_core_054 = input_a[14] | input_a[0];
  assign popcount29_hc56_core_055 = input_a[26] ^ input_a[8];
  assign popcount29_hc56_core_056 = ~(input_a[1] & input_a[2]);
  assign popcount29_hc56_core_057 = input_a[28] & input_a[17];
  assign popcount29_hc56_core_058 = input_a[20] & input_a[0];
  assign popcount29_hc56_core_059 = input_a[25] & input_a[5];
  assign popcount29_hc56_core_063 = ~(input_a[19] & input_a[8]);
  assign popcount29_hc56_core_067 = input_a[24] & input_a[12];
  assign popcount29_hc56_core_068 = input_a[11] ^ input_a[7];
  assign popcount29_hc56_core_069 = input_a[19] & input_a[7];
  assign popcount29_hc56_core_070 = ~(input_a[15] & input_a[24]);
  assign popcount29_hc56_core_072 = ~(input_a[3] | input_a[18]);
  assign popcount29_hc56_core_073 = input_a[10] ^ input_a[27];
  assign popcount29_hc56_core_074 = ~input_a[28];
  assign popcount29_hc56_core_076 = input_a[4] ^ input_a[18];
  assign popcount29_hc56_core_078 = input_a[3] | input_a[7];
  assign popcount29_hc56_core_080 = ~(input_a[23] ^ input_a[2]);
  assign popcount29_hc56_core_082 = ~(input_a[24] | input_a[19]);
  assign popcount29_hc56_core_086 = input_a[24] & input_a[12];
  assign popcount29_hc56_core_087 = ~(input_a[18] ^ input_a[12]);
  assign popcount29_hc56_core_088 = ~(input_a[13] | input_a[25]);
  assign popcount29_hc56_core_089 = ~input_a[13];
  assign popcount29_hc56_core_090 = ~(input_a[23] | input_a[17]);
  assign popcount29_hc56_core_091 = ~(input_a[28] | input_a[25]);
  assign popcount29_hc56_core_092 = ~(input_a[19] & input_a[3]);
  assign popcount29_hc56_core_094 = input_a[25] ^ input_a[7];
  assign popcount29_hc56_core_095 = ~(input_a[28] & input_a[9]);
  assign popcount29_hc56_core_096 = ~input_a[27];
  assign popcount29_hc56_core_097 = ~(input_a[19] ^ input_a[19]);
  assign popcount29_hc56_core_099 = input_a[1] & input_a[20];
  assign popcount29_hc56_core_100 = ~(input_a[25] | input_a[0]);
  assign popcount29_hc56_core_102 = input_a[9] | input_a[4];
  assign popcount29_hc56_core_103 = ~(input_a[8] & input_a[23]);
  assign popcount29_hc56_core_104 = ~(input_a[1] | input_a[1]);
  assign popcount29_hc56_core_107 = input_a[6] ^ input_a[23];
  assign popcount29_hc56_core_108 = ~(input_a[10] | input_a[22]);
  assign popcount29_hc56_core_109 = ~(input_a[8] ^ input_a[25]);
  assign popcount29_hc56_core_111 = input_a[15] & input_a[24];
  assign popcount29_hc56_core_112 = input_a[3] ^ input_a[11];
  assign popcount29_hc56_core_113 = input_a[0] & input_a[11];
  assign popcount29_hc56_core_114 = ~(input_a[8] ^ input_a[14]);
  assign popcount29_hc56_core_115 = input_a[27] & input_a[1];
  assign popcount29_hc56_core_117 = ~(input_a[24] | input_a[0]);
  assign popcount29_hc56_core_118 = ~(input_a[5] ^ input_a[27]);
  assign popcount29_hc56_core_119 = ~input_a[23];
  assign popcount29_hc56_core_121 = input_a[12] ^ input_a[12];
  assign popcount29_hc56_core_122 = ~input_a[21];
  assign popcount29_hc56_core_123 = ~(input_a[0] | input_a[0]);
  assign popcount29_hc56_core_124 = ~(input_a[18] | input_a[27]);
  assign popcount29_hc56_core_125 = input_a[11] | input_a[26];
  assign popcount29_hc56_core_126 = ~(input_a[11] | input_a[24]);
  assign popcount29_hc56_core_127 = input_a[11] | input_a[24];
  assign popcount29_hc56_core_128 = input_a[5] ^ input_a[14];
  assign popcount29_hc56_core_130 = ~input_a[27];
  assign popcount29_hc56_core_131 = input_a[25] ^ input_a[12];
  assign popcount29_hc56_core_132 = ~(input_a[24] ^ input_a[10]);
  assign popcount29_hc56_core_133 = input_a[2] | input_a[3];
  assign popcount29_hc56_core_134 = ~input_a[28];
  assign popcount29_hc56_core_135 = input_a[6] & input_a[17];
  assign popcount29_hc56_core_138 = input_a[16] | input_a[19];
  assign popcount29_hc56_core_139 = ~(input_a[17] | input_a[5]);
  assign popcount29_hc56_core_140 = input_a[20] ^ input_a[26];
  assign popcount29_hc56_core_144 = ~(input_a[24] | input_a[8]);
  assign popcount29_hc56_core_146 = input_a[26] & input_a[22];
  assign popcount29_hc56_core_147 = ~(input_a[8] & input_a[9]);
  assign popcount29_hc56_core_148 = ~(input_a[24] ^ input_a[13]);
  assign popcount29_hc56_core_149 = ~(input_a[13] ^ input_a[19]);
  assign popcount29_hc56_core_150 = input_a[15] ^ input_a[4];
  assign popcount29_hc56_core_151 = ~(input_a[13] & input_a[4]);
  assign popcount29_hc56_core_152 = ~(input_a[8] & input_a[8]);
  assign popcount29_hc56_core_154 = ~input_a[0];
  assign popcount29_hc56_core_156 = input_a[25] ^ input_a[16];
  assign popcount29_hc56_core_157 = ~input_a[15];
  assign popcount29_hc56_core_158 = input_a[14] ^ input_a[12];
  assign popcount29_hc56_core_159 = ~input_a[21];
  assign popcount29_hc56_core_161 = input_a[9] & input_a[9];
  assign popcount29_hc56_core_162 = input_a[5] | input_a[1];
  assign popcount29_hc56_core_163_not = ~input_a[12];
  assign popcount29_hc56_core_165 = input_a[7] ^ input_a[4];
  assign popcount29_hc56_core_166 = ~input_a[16];
  assign popcount29_hc56_core_168 = input_a[17] ^ input_a[20];
  assign popcount29_hc56_core_169 = ~input_a[28];
  assign popcount29_hc56_core_172 = input_a[23] | input_a[9];
  assign popcount29_hc56_core_173 = ~(input_a[11] | input_a[17]);
  assign popcount29_hc56_core_174 = ~input_a[25];
  assign popcount29_hc56_core_175 = input_a[21] ^ input_a[21];
  assign popcount29_hc56_core_176 = ~input_a[21];
  assign popcount29_hc56_core_178_not = ~input_a[26];
  assign popcount29_hc56_core_179 = ~input_a[21];
  assign popcount29_hc56_core_180 = ~(input_a[3] & input_a[21]);
  assign popcount29_hc56_core_183 = ~(input_a[24] ^ input_a[11]);
  assign popcount29_hc56_core_186 = ~input_a[18];
  assign popcount29_hc56_core_187_not = ~input_a[23];
  assign popcount29_hc56_core_188 = ~(input_a[20] ^ input_a[0]);
  assign popcount29_hc56_core_191 = input_a[27] | input_a[27];
  assign popcount29_hc56_core_192 = ~(input_a[8] ^ input_a[27]);
  assign popcount29_hc56_core_194 = input_a[24] ^ input_a[18];
  assign popcount29_hc56_core_195 = input_a[26] & input_a[12];
  assign popcount29_hc56_core_196 = ~(input_a[9] ^ input_a[27]);
  assign popcount29_hc56_core_197 = ~(input_a[27] | input_a[25]);
  assign popcount29_hc56_core_198 = input_a[22] & input_a[26];
  assign popcount29_hc56_core_199 = ~(input_a[13] & input_a[14]);
  assign popcount29_hc56_core_201 = input_a[18] ^ input_a[2];
  assign popcount29_hc56_core_203 = ~input_a[14];
  assign popcount29_hc56_core_204 = ~(input_a[28] ^ input_a[8]);
  assign popcount29_hc56_core_205 = input_a[1] ^ input_a[23];
  assign popcount29_hc56_core_206 = input_a[26] | input_a[2];
  assign popcount29_hc56_core_207 = input_a[15] & input_a[11];

  assign popcount29_hc56_out[0] = input_a[27];
  assign popcount29_hc56_out[1] = input_a[8];
  assign popcount29_hc56_out[2] = 1'b1;
  assign popcount29_hc56_out[3] = input_a[28];
  assign popcount29_hc56_out[4] = 1'b0;
endmodule