// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.13779
// WCE=12.0
// EP=0.991153%
// Printed PDK parameters:
//  Area=25202425.0
//  Delay=45485016.0
//  Power=1153800.0

module popcount24_mubj(input [23:0] input_a, output [4:0] popcount24_mubj_out);
  wire popcount24_mubj_core_027;
  wire popcount24_mubj_core_028;
  wire popcount24_mubj_core_029;
  wire popcount24_mubj_core_032;
  wire popcount24_mubj_core_033;
  wire popcount24_mubj_core_036;
  wire popcount24_mubj_core_038;
  wire popcount24_mubj_core_040;
  wire popcount24_mubj_core_041;
  wire popcount24_mubj_core_043;
  wire popcount24_mubj_core_046;
  wire popcount24_mubj_core_048;
  wire popcount24_mubj_core_049;
  wire popcount24_mubj_core_051;
  wire popcount24_mubj_core_052;
  wire popcount24_mubj_core_056;
  wire popcount24_mubj_core_059;
  wire popcount24_mubj_core_061;
  wire popcount24_mubj_core_062;
  wire popcount24_mubj_core_063;
  wire popcount24_mubj_core_064;
  wire popcount24_mubj_core_065;
  wire popcount24_mubj_core_066;
  wire popcount24_mubj_core_068;
  wire popcount24_mubj_core_069;
  wire popcount24_mubj_core_070;
  wire popcount24_mubj_core_074;
  wire popcount24_mubj_core_075;
  wire popcount24_mubj_core_076;
  wire popcount24_mubj_core_078;
  wire popcount24_mubj_core_080;
  wire popcount24_mubj_core_081;
  wire popcount24_mubj_core_082;
  wire popcount24_mubj_core_083;
  wire popcount24_mubj_core_084;
  wire popcount24_mubj_core_085;
  wire popcount24_mubj_core_091;
  wire popcount24_mubj_core_093;
  wire popcount24_mubj_core_094;
  wire popcount24_mubj_core_096;
  wire popcount24_mubj_core_098;
  wire popcount24_mubj_core_099;
  wire popcount24_mubj_core_100;
  wire popcount24_mubj_core_101;
  wire popcount24_mubj_core_103;
  wire popcount24_mubj_core_104;
  wire popcount24_mubj_core_105_not;
  wire popcount24_mubj_core_106;
  wire popcount24_mubj_core_107;
  wire popcount24_mubj_core_108;
  wire popcount24_mubj_core_109;
  wire popcount24_mubj_core_110;
  wire popcount24_mubj_core_112;
  wire popcount24_mubj_core_114;
  wire popcount24_mubj_core_115;
  wire popcount24_mubj_core_116;
  wire popcount24_mubj_core_117;
  wire popcount24_mubj_core_118;
  wire popcount24_mubj_core_119;
  wire popcount24_mubj_core_121;
  wire popcount24_mubj_core_122;
  wire popcount24_mubj_core_123;
  wire popcount24_mubj_core_124;
  wire popcount24_mubj_core_125;
  wire popcount24_mubj_core_126;
  wire popcount24_mubj_core_127;
  wire popcount24_mubj_core_129;
  wire popcount24_mubj_core_130;
  wire popcount24_mubj_core_131;
  wire popcount24_mubj_core_132;
  wire popcount24_mubj_core_133;
  wire popcount24_mubj_core_137;
  wire popcount24_mubj_core_138;
  wire popcount24_mubj_core_139;
  wire popcount24_mubj_core_140;
  wire popcount24_mubj_core_141;
  wire popcount24_mubj_core_142;
  wire popcount24_mubj_core_144;
  wire popcount24_mubj_core_145;
  wire popcount24_mubj_core_146;
  wire popcount24_mubj_core_147;
  wire popcount24_mubj_core_148;
  wire popcount24_mubj_core_149;
  wire popcount24_mubj_core_150;
  wire popcount24_mubj_core_152;
  wire popcount24_mubj_core_154;
  wire popcount24_mubj_core_155;
  wire popcount24_mubj_core_156;
  wire popcount24_mubj_core_158;
  wire popcount24_mubj_core_159;
  wire popcount24_mubj_core_160;
  wire popcount24_mubj_core_161;
  wire popcount24_mubj_core_163;
  wire popcount24_mubj_core_164;
  wire popcount24_mubj_core_165;
  wire popcount24_mubj_core_166;
  wire popcount24_mubj_core_167;
  wire popcount24_mubj_core_168;
  wire popcount24_mubj_core_169;
  wire popcount24_mubj_core_170;
  wire popcount24_mubj_core_171;
  wire popcount24_mubj_core_172;
  wire popcount24_mubj_core_173;
  wire popcount24_mubj_core_174;
  wire popcount24_mubj_core_175;
  wire popcount24_mubj_core_177;

  assign popcount24_mubj_core_027 = input_a[14] & input_a[2];
  assign popcount24_mubj_core_028 = input_a[19] ^ input_a[11];
  assign popcount24_mubj_core_029 = input_a[2] | input_a[18];
  assign popcount24_mubj_core_032 = input_a[10] & input_a[10];
  assign popcount24_mubj_core_033 = input_a[21] | input_a[10];
  assign popcount24_mubj_core_036 = input_a[4] | input_a[1];
  assign popcount24_mubj_core_038 = input_a[18] | input_a[16];
  assign popcount24_mubj_core_040 = popcount24_mubj_core_027 ^ popcount24_mubj_core_036;
  assign popcount24_mubj_core_041 = popcount24_mubj_core_027 & popcount24_mubj_core_036;
  assign popcount24_mubj_core_043 = input_a[6] | input_a[22];
  assign popcount24_mubj_core_046 = input_a[5] ^ input_a[20];
  assign popcount24_mubj_core_048 = input_a[3] & input_a[5];
  assign popcount24_mubj_core_049 = input_a[2] & input_a[3];
  assign popcount24_mubj_core_051 = ~(input_a[17] | input_a[11]);
  assign popcount24_mubj_core_052 = input_a[6] & input_a[10];
  assign popcount24_mubj_core_056 = input_a[17] | input_a[5];
  assign popcount24_mubj_core_059 = input_a[3] | input_a[9];
  assign popcount24_mubj_core_061 = ~input_a[7];
  assign popcount24_mubj_core_062 = input_a[10] & input_a[19];
  assign popcount24_mubj_core_063 = input_a[17] ^ input_a[22];
  assign popcount24_mubj_core_064 = ~(input_a[19] ^ input_a[15]);
  assign popcount24_mubj_core_065 = ~input_a[18];
  assign popcount24_mubj_core_066 = input_a[9] | input_a[11];
  assign popcount24_mubj_core_068 = input_a[13] & input_a[9];
  assign popcount24_mubj_core_069 = input_a[23] | input_a[10];
  assign popcount24_mubj_core_070 = input_a[12] & input_a[22];
  assign popcount24_mubj_core_074 = input_a[23] | input_a[6];
  assign popcount24_mubj_core_075 = input_a[17] & input_a[0];
  assign popcount24_mubj_core_076 = popcount24_mubj_core_040 ^ popcount24_mubj_core_066;
  assign popcount24_mubj_core_078 = ~popcount24_mubj_core_076;
  assign popcount24_mubj_core_080 = popcount24_mubj_core_040 | popcount24_mubj_core_076;
  assign popcount24_mubj_core_081 = popcount24_mubj_core_041 ^ popcount24_mubj_core_069;
  assign popcount24_mubj_core_082 = popcount24_mubj_core_041 & popcount24_mubj_core_069;
  assign popcount24_mubj_core_083 = popcount24_mubj_core_081 ^ popcount24_mubj_core_080;
  assign popcount24_mubj_core_084 = popcount24_mubj_core_081 & popcount24_mubj_core_080;
  assign popcount24_mubj_core_085 = popcount24_mubj_core_082 | popcount24_mubj_core_084;
  assign popcount24_mubj_core_091 = ~(input_a[4] & input_a[5]);
  assign popcount24_mubj_core_093 = input_a[16] | input_a[10];
  assign popcount24_mubj_core_094 = input_a[17] & input_a[5];
  assign popcount24_mubj_core_096 = input_a[12] ^ input_a[23];
  assign popcount24_mubj_core_098 = input_a[16] & input_a[17];
  assign popcount24_mubj_core_099 = ~input_a[15];
  assign popcount24_mubj_core_100 = ~(input_a[0] & input_a[19]);
  assign popcount24_mubj_core_101 = popcount24_mubj_core_098 ^ input_a[15];
  assign popcount24_mubj_core_103 = input_a[12] ^ popcount24_mubj_core_099;
  assign popcount24_mubj_core_104 = input_a[12] & popcount24_mubj_core_099;
  assign popcount24_mubj_core_105_not = ~popcount24_mubj_core_101;
  assign popcount24_mubj_core_106 = input_a[17] & input_a[16];
  assign popcount24_mubj_core_107 = popcount24_mubj_core_105_not ^ popcount24_mubj_core_104;
  assign popcount24_mubj_core_108 = ~(input_a[8] | input_a[9]);
  assign popcount24_mubj_core_109 = popcount24_mubj_core_106 | input_a[12];
  assign popcount24_mubj_core_110 = input_a[13] | input_a[23];
  assign popcount24_mubj_core_112 = input_a[15] | popcount24_mubj_core_109;
  assign popcount24_mubj_core_114 = input_a[9] & input_a[11];
  assign popcount24_mubj_core_115 = input_a[4] | input_a[5];
  assign popcount24_mubj_core_116 = input_a[19] & input_a[20];
  assign popcount24_mubj_core_117 = ~(input_a[23] | input_a[1]);
  assign popcount24_mubj_core_118 = input_a[18] & input_a[7];
  assign popcount24_mubj_core_119 = popcount24_mubj_core_116 | popcount24_mubj_core_118;
  assign popcount24_mubj_core_121 = input_a[22] | input_a[21];
  assign popcount24_mubj_core_122 = input_a[0] & input_a[22];
  assign popcount24_mubj_core_123 = input_a[0] | input_a[23];
  assign popcount24_mubj_core_124 = input_a[21] & input_a[5];
  assign popcount24_mubj_core_125 = popcount24_mubj_core_122 | popcount24_mubj_core_124;
  assign popcount24_mubj_core_126 = ~(input_a[9] & input_a[9]);
  assign popcount24_mubj_core_127 = input_a[16] | input_a[16];
  assign popcount24_mubj_core_129 = popcount24_mubj_core_119 ^ popcount24_mubj_core_125;
  assign popcount24_mubj_core_130 = popcount24_mubj_core_119 & popcount24_mubj_core_125;
  assign popcount24_mubj_core_131 = popcount24_mubj_core_129 ^ input_a[8];
  assign popcount24_mubj_core_132 = popcount24_mubj_core_129 & input_a[8];
  assign popcount24_mubj_core_133 = popcount24_mubj_core_130 | popcount24_mubj_core_132;
  assign popcount24_mubj_core_137 = input_a[13] ^ input_a[1];
  assign popcount24_mubj_core_138 = ~(input_a[6] & input_a[11]);
  assign popcount24_mubj_core_139 = ~(input_a[18] ^ input_a[16]);
  assign popcount24_mubj_core_140 = popcount24_mubj_core_103 & input_a[3];
  assign popcount24_mubj_core_141 = input_a[16] & input_a[12];
  assign popcount24_mubj_core_142 = popcount24_mubj_core_107 & popcount24_mubj_core_131;
  assign popcount24_mubj_core_144 = input_a[13] & popcount24_mubj_core_140;
  assign popcount24_mubj_core_145 = popcount24_mubj_core_142 | popcount24_mubj_core_144;
  assign popcount24_mubj_core_146 = popcount24_mubj_core_112 ^ popcount24_mubj_core_133;
  assign popcount24_mubj_core_147 = popcount24_mubj_core_112 & popcount24_mubj_core_133;
  assign popcount24_mubj_core_148 = popcount24_mubj_core_146 ^ popcount24_mubj_core_145;
  assign popcount24_mubj_core_149 = popcount24_mubj_core_146 & popcount24_mubj_core_145;
  assign popcount24_mubj_core_150 = popcount24_mubj_core_147 | popcount24_mubj_core_149;
  assign popcount24_mubj_core_152 = ~(input_a[5] & input_a[1]);
  assign popcount24_mubj_core_154 = input_a[11] ^ input_a[5];
  assign popcount24_mubj_core_155 = ~(input_a[21] & input_a[21]);
  assign popcount24_mubj_core_156 = ~(input_a[23] & input_a[2]);
  assign popcount24_mubj_core_158 = popcount24_mubj_core_078 ^ input_a[6];
  assign popcount24_mubj_core_159 = popcount24_mubj_core_078 & input_a[6];
  assign popcount24_mubj_core_160 = input_a[20] & input_a[19];
  assign popcount24_mubj_core_161 = input_a[7] ^ input_a[16];
  assign popcount24_mubj_core_163 = popcount24_mubj_core_083 ^ popcount24_mubj_core_148;
  assign popcount24_mubj_core_164 = popcount24_mubj_core_083 & popcount24_mubj_core_148;
  assign popcount24_mubj_core_165 = popcount24_mubj_core_163 ^ popcount24_mubj_core_159;
  assign popcount24_mubj_core_166 = popcount24_mubj_core_163 & popcount24_mubj_core_159;
  assign popcount24_mubj_core_167 = popcount24_mubj_core_164 | popcount24_mubj_core_166;
  assign popcount24_mubj_core_168 = popcount24_mubj_core_085 | popcount24_mubj_core_150;
  assign popcount24_mubj_core_169 = popcount24_mubj_core_085 & popcount24_mubj_core_150;
  assign popcount24_mubj_core_170 = input_a[20] & input_a[16];
  assign popcount24_mubj_core_171 = popcount24_mubj_core_168 & popcount24_mubj_core_167;
  assign popcount24_mubj_core_172 = popcount24_mubj_core_169 | popcount24_mubj_core_171;
  assign popcount24_mubj_core_173 = ~(input_a[2] & input_a[10]);
  assign popcount24_mubj_core_174 = ~input_a[18];
  assign popcount24_mubj_core_175 = ~(input_a[21] & input_a[6]);
  assign popcount24_mubj_core_177 = ~(input_a[6] | input_a[23]);

  assign popcount24_mubj_out[0] = popcount24_mubj_core_164;
  assign popcount24_mubj_out[1] = popcount24_mubj_core_158;
  assign popcount24_mubj_out[2] = popcount24_mubj_core_165;
  assign popcount24_mubj_out[3] = 1'b0;
  assign popcount24_mubj_out[4] = popcount24_mubj_core_172;
endmodule