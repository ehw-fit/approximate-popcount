// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.55435
// WCE=20.0
// EP=0.98678%
// Printed PDK parameters:
//  Area=46253898.0
//  Delay=84290448.0
//  Power=1981600.0

module popcount39_ub2f(input [38:0] input_a, output [5:0] popcount39_ub2f_out);
  wire popcount39_ub2f_core_041;
  wire popcount39_ub2f_core_042;
  wire popcount39_ub2f_core_043;
  wire popcount39_ub2f_core_044;
  wire popcount39_ub2f_core_045;
  wire popcount39_ub2f_core_046;
  wire popcount39_ub2f_core_047;
  wire popcount39_ub2f_core_048;
  wire popcount39_ub2f_core_049;
  wire popcount39_ub2f_core_050;
  wire popcount39_ub2f_core_052;
  wire popcount39_ub2f_core_053;
  wire popcount39_ub2f_core_054;
  wire popcount39_ub2f_core_055;
  wire popcount39_ub2f_core_056;
  wire popcount39_ub2f_core_057;
  wire popcount39_ub2f_core_061;
  wire popcount39_ub2f_core_062;
  wire popcount39_ub2f_core_063;
  wire popcount39_ub2f_core_070;
  wire popcount39_ub2f_core_072;
  wire popcount39_ub2f_core_074;
  wire popcount39_ub2f_core_075;
  wire popcount39_ub2f_core_076;
  wire popcount39_ub2f_core_077;
  wire popcount39_ub2f_core_078;
  wire popcount39_ub2f_core_079;
  wire popcount39_ub2f_core_082;
  wire popcount39_ub2f_core_083;
  wire popcount39_ub2f_core_084;
  wire popcount39_ub2f_core_085;
  wire popcount39_ub2f_core_086;
  wire popcount39_ub2f_core_087;
  wire popcount39_ub2f_core_088;
  wire popcount39_ub2f_core_089;
  wire popcount39_ub2f_core_091;
  wire popcount39_ub2f_core_092;
  wire popcount39_ub2f_core_093;
  wire popcount39_ub2f_core_094;
  wire popcount39_ub2f_core_095;
  wire popcount39_ub2f_core_096;
  wire popcount39_ub2f_core_097;
  wire popcount39_ub2f_core_099;
  wire popcount39_ub2f_core_101;
  wire popcount39_ub2f_core_103;
  wire popcount39_ub2f_core_104;
  wire popcount39_ub2f_core_105;
  wire popcount39_ub2f_core_106;
  wire popcount39_ub2f_core_108;
  wire popcount39_ub2f_core_109;
  wire popcount39_ub2f_core_110;
  wire popcount39_ub2f_core_111;
  wire popcount39_ub2f_core_113;
  wire popcount39_ub2f_core_116;
  wire popcount39_ub2f_core_118;
  wire popcount39_ub2f_core_119;
  wire popcount39_ub2f_core_120;
  wire popcount39_ub2f_core_121;
  wire popcount39_ub2f_core_122;
  wire popcount39_ub2f_core_123;
  wire popcount39_ub2f_core_124;
  wire popcount39_ub2f_core_125;
  wire popcount39_ub2f_core_126;
  wire popcount39_ub2f_core_127;
  wire popcount39_ub2f_core_128;
  wire popcount39_ub2f_core_130;
  wire popcount39_ub2f_core_133;
  wire popcount39_ub2f_core_134;
  wire popcount39_ub2f_core_135;
  wire popcount39_ub2f_core_136;
  wire popcount39_ub2f_core_138;
  wire popcount39_ub2f_core_139;
  wire popcount39_ub2f_core_141;
  wire popcount39_ub2f_core_142;
  wire popcount39_ub2f_core_143;
  wire popcount39_ub2f_core_144;
  wire popcount39_ub2f_core_145;
  wire popcount39_ub2f_core_146;
  wire popcount39_ub2f_core_147;
  wire popcount39_ub2f_core_148;
  wire popcount39_ub2f_core_149;
  wire popcount39_ub2f_core_150;
  wire popcount39_ub2f_core_151;
  wire popcount39_ub2f_core_153;
  wire popcount39_ub2f_core_154;
  wire popcount39_ub2f_core_156;
  wire popcount39_ub2f_core_157;
  wire popcount39_ub2f_core_158;
  wire popcount39_ub2f_core_159;
  wire popcount39_ub2f_core_160;
  wire popcount39_ub2f_core_161;
  wire popcount39_ub2f_core_162;
  wire popcount39_ub2f_core_163;
  wire popcount39_ub2f_core_166;
  wire popcount39_ub2f_core_168;
  wire popcount39_ub2f_core_169;
  wire popcount39_ub2f_core_170;
  wire popcount39_ub2f_core_171;
  wire popcount39_ub2f_core_175;
  wire popcount39_ub2f_core_176;
  wire popcount39_ub2f_core_180;
  wire popcount39_ub2f_core_181;
  wire popcount39_ub2f_core_183;
  wire popcount39_ub2f_core_184;
  wire popcount39_ub2f_core_185;
  wire popcount39_ub2f_core_186;
  wire popcount39_ub2f_core_187;
  wire popcount39_ub2f_core_188;
  wire popcount39_ub2f_core_189;
  wire popcount39_ub2f_core_191;
  wire popcount39_ub2f_core_192;
  wire popcount39_ub2f_core_193;
  wire popcount39_ub2f_core_195;
  wire popcount39_ub2f_core_196;
  wire popcount39_ub2f_core_197;
  wire popcount39_ub2f_core_200;
  wire popcount39_ub2f_core_201_not;
  wire popcount39_ub2f_core_202;
  wire popcount39_ub2f_core_206;
  wire popcount39_ub2f_core_207;
  wire popcount39_ub2f_core_208;
  wire popcount39_ub2f_core_209;
  wire popcount39_ub2f_core_210;
  wire popcount39_ub2f_core_212;
  wire popcount39_ub2f_core_213;
  wire popcount39_ub2f_core_215;
  wire popcount39_ub2f_core_216;
  wire popcount39_ub2f_core_218;
  wire popcount39_ub2f_core_219;
  wire popcount39_ub2f_core_220;
  wire popcount39_ub2f_core_225;
  wire popcount39_ub2f_core_226;
  wire popcount39_ub2f_core_227;
  wire popcount39_ub2f_core_228;
  wire popcount39_ub2f_core_229;
  wire popcount39_ub2f_core_232;
  wire popcount39_ub2f_core_235;
  wire popcount39_ub2f_core_236;
  wire popcount39_ub2f_core_241;
  wire popcount39_ub2f_core_244;
  wire popcount39_ub2f_core_245;
  wire popcount39_ub2f_core_247;
  wire popcount39_ub2f_core_248;
  wire popcount39_ub2f_core_249;
  wire popcount39_ub2f_core_250;
  wire popcount39_ub2f_core_251;
  wire popcount39_ub2f_core_252;
  wire popcount39_ub2f_core_256;
  wire popcount39_ub2f_core_258;
  wire popcount39_ub2f_core_259;
  wire popcount39_ub2f_core_261;
  wire popcount39_ub2f_core_262;
  wire popcount39_ub2f_core_264;
  wire popcount39_ub2f_core_266;
  wire popcount39_ub2f_core_268;
  wire popcount39_ub2f_core_269;
  wire popcount39_ub2f_core_271;
  wire popcount39_ub2f_core_273;
  wire popcount39_ub2f_core_274;
  wire popcount39_ub2f_core_277;
  wire popcount39_ub2f_core_278;
  wire popcount39_ub2f_core_279;
  wire popcount39_ub2f_core_280;
  wire popcount39_ub2f_core_281;
  wire popcount39_ub2f_core_282;
  wire popcount39_ub2f_core_283;
  wire popcount39_ub2f_core_284;
  wire popcount39_ub2f_core_285;
  wire popcount39_ub2f_core_287;
  wire popcount39_ub2f_core_288;
  wire popcount39_ub2f_core_290;
  wire popcount39_ub2f_core_292;
  wire popcount39_ub2f_core_293;
  wire popcount39_ub2f_core_294;
  wire popcount39_ub2f_core_295;
  wire popcount39_ub2f_core_296;
  wire popcount39_ub2f_core_299;
  wire popcount39_ub2f_core_300;
  wire popcount39_ub2f_core_304;
  wire popcount39_ub2f_core_305;
  wire popcount39_ub2f_core_306;

  assign popcount39_ub2f_core_041 = ~(input_a[26] ^ input_a[38]);
  assign popcount39_ub2f_core_042 = input_a[38] & input_a[22];
  assign popcount39_ub2f_core_043 = ~input_a[5];
  assign popcount39_ub2f_core_044 = input_a[2] & input_a[21];
  assign popcount39_ub2f_core_045 = input_a[2] & input_a[15];
  assign popcount39_ub2f_core_046 = input_a[16] & input_a[0];
  assign popcount39_ub2f_core_047 = popcount39_ub2f_core_042 | popcount39_ub2f_core_044;
  assign popcount39_ub2f_core_048 = popcount39_ub2f_core_042 & popcount39_ub2f_core_044;
  assign popcount39_ub2f_core_049 = popcount39_ub2f_core_047 | popcount39_ub2f_core_046;
  assign popcount39_ub2f_core_050 = input_a[34] ^ input_a[14];
  assign popcount39_ub2f_core_052 = input_a[4] ^ input_a[5];
  assign popcount39_ub2f_core_053 = input_a[4] & input_a[5];
  assign popcount39_ub2f_core_054 = input_a[12] ^ input_a[7];
  assign popcount39_ub2f_core_055 = input_a[15] & input_a[23];
  assign popcount39_ub2f_core_056 = input_a[28] & input_a[5];
  assign popcount39_ub2f_core_057 = ~input_a[27];
  assign popcount39_ub2f_core_061 = input_a[15] ^ input_a[16];
  assign popcount39_ub2f_core_062 = popcount39_ub2f_core_053 ^ popcount39_ub2f_core_055;
  assign popcount39_ub2f_core_063 = popcount39_ub2f_core_053 & popcount39_ub2f_core_055;
  assign popcount39_ub2f_core_070 = input_a[26] & popcount39_ub2f_core_052;
  assign popcount39_ub2f_core_072 = popcount39_ub2f_core_049 & popcount39_ub2f_core_062;
  assign popcount39_ub2f_core_074 = popcount39_ub2f_core_049 & popcount39_ub2f_core_070;
  assign popcount39_ub2f_core_075 = popcount39_ub2f_core_072 | popcount39_ub2f_core_074;
  assign popcount39_ub2f_core_076 = popcount39_ub2f_core_048 ^ popcount39_ub2f_core_063;
  assign popcount39_ub2f_core_077 = popcount39_ub2f_core_048 & popcount39_ub2f_core_063;
  assign popcount39_ub2f_core_078 = popcount39_ub2f_core_076 | popcount39_ub2f_core_075;
  assign popcount39_ub2f_core_079 = ~input_a[36];
  assign popcount39_ub2f_core_082 = ~input_a[22];
  assign popcount39_ub2f_core_083 = input_a[9] & input_a[14];
  assign popcount39_ub2f_core_084 = input_a[9] & input_a[10];
  assign popcount39_ub2f_core_085 = input_a[12] | input_a[13];
  assign popcount39_ub2f_core_086 = input_a[12] & input_a[13];
  assign popcount39_ub2f_core_087 = ~input_a[10];
  assign popcount39_ub2f_core_088 = input_a[11] & popcount39_ub2f_core_085;
  assign popcount39_ub2f_core_089 = popcount39_ub2f_core_086 | popcount39_ub2f_core_088;
  assign popcount39_ub2f_core_091 = ~input_a[26];
  assign popcount39_ub2f_core_092 = input_a[3] & input_a[1];
  assign popcount39_ub2f_core_093 = popcount39_ub2f_core_084 ^ popcount39_ub2f_core_089;
  assign popcount39_ub2f_core_094 = popcount39_ub2f_core_084 & popcount39_ub2f_core_089;
  assign popcount39_ub2f_core_095 = popcount39_ub2f_core_093 ^ popcount39_ub2f_core_092;
  assign popcount39_ub2f_core_096 = popcount39_ub2f_core_093 & popcount39_ub2f_core_092;
  assign popcount39_ub2f_core_097 = popcount39_ub2f_core_094 | popcount39_ub2f_core_096;
  assign popcount39_ub2f_core_099 = input_a[4] & input_a[17];
  assign popcount39_ub2f_core_101 = input_a[14] & input_a[20];
  assign popcount39_ub2f_core_103 = input_a[6] & input_a[18];
  assign popcount39_ub2f_core_104 = input_a[17] | input_a[31];
  assign popcount39_ub2f_core_105 = input_a[8] & input_a[25];
  assign popcount39_ub2f_core_106 = popcount39_ub2f_core_103 | popcount39_ub2f_core_105;
  assign popcount39_ub2f_core_108 = input_a[4] & input_a[4];
  assign popcount39_ub2f_core_109 = ~(input_a[22] ^ input_a[0]);
  assign popcount39_ub2f_core_110 = popcount39_ub2f_core_101 ^ popcount39_ub2f_core_106;
  assign popcount39_ub2f_core_111 = popcount39_ub2f_core_101 & popcount39_ub2f_core_106;
  assign popcount39_ub2f_core_113 = input_a[24] & input_a[3];
  assign popcount39_ub2f_core_116 = ~(input_a[19] ^ input_a[17]);
  assign popcount39_ub2f_core_118 = input_a[27] & input_a[33];
  assign popcount39_ub2f_core_119 = popcount39_ub2f_core_095 ^ popcount39_ub2f_core_110;
  assign popcount39_ub2f_core_120 = popcount39_ub2f_core_095 & popcount39_ub2f_core_110;
  assign popcount39_ub2f_core_121 = popcount39_ub2f_core_119 ^ popcount39_ub2f_core_118;
  assign popcount39_ub2f_core_122 = popcount39_ub2f_core_119 & popcount39_ub2f_core_118;
  assign popcount39_ub2f_core_123 = popcount39_ub2f_core_120 | popcount39_ub2f_core_122;
  assign popcount39_ub2f_core_124 = popcount39_ub2f_core_097 ^ popcount39_ub2f_core_111;
  assign popcount39_ub2f_core_125 = popcount39_ub2f_core_097 & popcount39_ub2f_core_111;
  assign popcount39_ub2f_core_126 = popcount39_ub2f_core_124 ^ popcount39_ub2f_core_123;
  assign popcount39_ub2f_core_127 = popcount39_ub2f_core_124 & popcount39_ub2f_core_123;
  assign popcount39_ub2f_core_128 = popcount39_ub2f_core_125 | popcount39_ub2f_core_127;
  assign popcount39_ub2f_core_130 = input_a[8] ^ input_a[3];
  assign popcount39_ub2f_core_133 = input_a[17] | input_a[29];
  assign popcount39_ub2f_core_134 = input_a[32] & input_a[13];
  assign popcount39_ub2f_core_135 = input_a[13] ^ input_a[23];
  assign popcount39_ub2f_core_136 = ~(input_a[34] & input_a[28]);
  assign popcount39_ub2f_core_138 = ~input_a[21];
  assign popcount39_ub2f_core_139 = ~(input_a[16] ^ input_a[1]);
  assign popcount39_ub2f_core_141 = popcount39_ub2f_core_078 ^ popcount39_ub2f_core_126;
  assign popcount39_ub2f_core_142 = popcount39_ub2f_core_078 & popcount39_ub2f_core_126;
  assign popcount39_ub2f_core_143 = popcount39_ub2f_core_141 ^ popcount39_ub2f_core_121;
  assign popcount39_ub2f_core_144 = popcount39_ub2f_core_141 & popcount39_ub2f_core_121;
  assign popcount39_ub2f_core_145 = popcount39_ub2f_core_142 | popcount39_ub2f_core_144;
  assign popcount39_ub2f_core_146 = popcount39_ub2f_core_077 ^ popcount39_ub2f_core_128;
  assign popcount39_ub2f_core_147 = popcount39_ub2f_core_077 & popcount39_ub2f_core_128;
  assign popcount39_ub2f_core_148 = popcount39_ub2f_core_146 ^ popcount39_ub2f_core_145;
  assign popcount39_ub2f_core_149 = popcount39_ub2f_core_146 & popcount39_ub2f_core_145;
  assign popcount39_ub2f_core_150 = popcount39_ub2f_core_147 | popcount39_ub2f_core_149;
  assign popcount39_ub2f_core_151 = input_a[34] | popcount39_ub2f_core_133;
  assign popcount39_ub2f_core_153 = popcount39_ub2f_core_151 ^ popcount39_ub2f_core_150;
  assign popcount39_ub2f_core_154 = popcount39_ub2f_core_151 & popcount39_ub2f_core_150;
  assign popcount39_ub2f_core_156 = input_a[34] ^ input_a[35];
  assign popcount39_ub2f_core_157 = ~(input_a[37] ^ input_a[14]);
  assign popcount39_ub2f_core_158 = ~(input_a[30] & input_a[1]);
  assign popcount39_ub2f_core_159 = ~(input_a[22] & input_a[7]);
  assign popcount39_ub2f_core_160 = ~input_a[13];
  assign popcount39_ub2f_core_161 = input_a[22] & input_a[2];
  assign popcount39_ub2f_core_162 = ~(input_a[7] & input_a[27]);
  assign popcount39_ub2f_core_163 = ~(input_a[4] | input_a[17]);
  assign popcount39_ub2f_core_166 = ~input_a[30];
  assign popcount39_ub2f_core_168 = ~(input_a[9] & input_a[21]);
  assign popcount39_ub2f_core_169 = ~(input_a[34] | input_a[5]);
  assign popcount39_ub2f_core_170 = ~(input_a[2] | input_a[10]);
  assign popcount39_ub2f_core_171 = ~(input_a[30] | input_a[26]);
  assign popcount39_ub2f_core_175 = input_a[37] & input_a[25];
  assign popcount39_ub2f_core_176 = input_a[16] ^ input_a[8];
  assign popcount39_ub2f_core_180 = input_a[30] ^ input_a[15];
  assign popcount39_ub2f_core_181 = input_a[18] | input_a[2];
  assign popcount39_ub2f_core_183 = ~input_a[31];
  assign popcount39_ub2f_core_184 = input_a[31] & input_a[38];
  assign popcount39_ub2f_core_185 = input_a[30] ^ input_a[3];
  assign popcount39_ub2f_core_186 = ~input_a[32];
  assign popcount39_ub2f_core_187 = ~(input_a[17] & input_a[15]);
  assign popcount39_ub2f_core_188 = input_a[31] | input_a[36];
  assign popcount39_ub2f_core_189 = input_a[8] ^ input_a[15];
  assign popcount39_ub2f_core_191 = ~input_a[36];
  assign popcount39_ub2f_core_192 = ~(input_a[30] & input_a[23]);
  assign popcount39_ub2f_core_193 = ~(input_a[31] & input_a[1]);
  assign popcount39_ub2f_core_195 = ~(input_a[11] ^ input_a[1]);
  assign popcount39_ub2f_core_196 = ~(input_a[17] ^ input_a[27]);
  assign popcount39_ub2f_core_197 = ~(input_a[16] ^ input_a[8]);
  assign popcount39_ub2f_core_200 = ~(input_a[36] | input_a[37]);
  assign popcount39_ub2f_core_201_not = ~input_a[20];
  assign popcount39_ub2f_core_202 = input_a[20] ^ input_a[3];
  assign popcount39_ub2f_core_206 = ~(input_a[36] | input_a[19]);
  assign popcount39_ub2f_core_207 = input_a[15] ^ input_a[21];
  assign popcount39_ub2f_core_208 = input_a[32] & input_a[37];
  assign popcount39_ub2f_core_209 = input_a[7] | input_a[22];
  assign popcount39_ub2f_core_210 = ~(input_a[13] & input_a[9]);
  assign popcount39_ub2f_core_212 = input_a[26] | input_a[36];
  assign popcount39_ub2f_core_213 = input_a[35] & input_a[24];
  assign popcount39_ub2f_core_215 = ~(input_a[32] ^ input_a[14]);
  assign popcount39_ub2f_core_216 = input_a[28] | input_a[36];
  assign popcount39_ub2f_core_218 = popcount39_ub2f_core_208 & popcount39_ub2f_core_213;
  assign popcount39_ub2f_core_219 = ~(input_a[36] & input_a[17]);
  assign popcount39_ub2f_core_220 = ~input_a[19];
  assign popcount39_ub2f_core_225 = input_a[7] & input_a[36];
  assign popcount39_ub2f_core_226 = input_a[37] ^ input_a[37];
  assign popcount39_ub2f_core_227 = input_a[28] & input_a[30];
  assign popcount39_ub2f_core_228 = ~input_a[13];
  assign popcount39_ub2f_core_229 = input_a[26] | input_a[24];
  assign popcount39_ub2f_core_232 = input_a[26] ^ input_a[11];
  assign popcount39_ub2f_core_235 = popcount39_ub2f_core_225 & popcount39_ub2f_core_227;
  assign popcount39_ub2f_core_236 = ~(input_a[2] ^ input_a[16]);
  assign popcount39_ub2f_core_241 = ~(input_a[31] & input_a[5]);
  assign popcount39_ub2f_core_244 = ~input_a[29];
  assign popcount39_ub2f_core_245 = input_a[15] ^ input_a[24];
  assign popcount39_ub2f_core_247 = input_a[31] | input_a[19];
  assign popcount39_ub2f_core_248 = popcount39_ub2f_core_218 ^ popcount39_ub2f_core_235;
  assign popcount39_ub2f_core_249 = popcount39_ub2f_core_218 & popcount39_ub2f_core_235;
  assign popcount39_ub2f_core_250 = popcount39_ub2f_core_248 ^ popcount39_ub2f_core_247;
  assign popcount39_ub2f_core_251 = popcount39_ub2f_core_248 & popcount39_ub2f_core_247;
  assign popcount39_ub2f_core_252 = popcount39_ub2f_core_249 | popcount39_ub2f_core_251;
  assign popcount39_ub2f_core_256 = input_a[10] ^ input_a[6];
  assign popcount39_ub2f_core_258 = ~(input_a[2] | input_a[17]);
  assign popcount39_ub2f_core_259 = input_a[12] & input_a[30];
  assign popcount39_ub2f_core_261 = ~(input_a[28] & input_a[9]);
  assign popcount39_ub2f_core_262 = input_a[16] | input_a[19];
  assign popcount39_ub2f_core_264 = input_a[16] & input_a[17];
  assign popcount39_ub2f_core_266 = input_a[3] & input_a[2];
  assign popcount39_ub2f_core_268 = input_a[24] | input_a[15];
  assign popcount39_ub2f_core_269 = ~input_a[32];
  assign popcount39_ub2f_core_271 = input_a[4] & input_a[20];
  assign popcount39_ub2f_core_273 = input_a[4] | input_a[14];
  assign popcount39_ub2f_core_274 = input_a[23] & input_a[1];
  assign popcount39_ub2f_core_277 = input_a[25] & input_a[33];
  assign popcount39_ub2f_core_278 = input_a[14] | input_a[26];
  assign popcount39_ub2f_core_279 = input_a[29] | input_a[27];
  assign popcount39_ub2f_core_280 = ~input_a[6];
  assign popcount39_ub2f_core_281 = input_a[6] ^ input_a[32];
  assign popcount39_ub2f_core_282 = ~input_a[22];
  assign popcount39_ub2f_core_283 = ~(input_a[7] | input_a[35]);
  assign popcount39_ub2f_core_284 = ~(input_a[4] & input_a[30]);
  assign popcount39_ub2f_core_285 = input_a[23] & input_a[6];
  assign popcount39_ub2f_core_287 = popcount39_ub2f_core_143 ^ popcount39_ub2f_core_250;
  assign popcount39_ub2f_core_288 = popcount39_ub2f_core_143 & popcount39_ub2f_core_250;
  assign popcount39_ub2f_core_290 = ~(input_a[1] ^ input_a[12]);
  assign popcount39_ub2f_core_292 = popcount39_ub2f_core_148 ^ popcount39_ub2f_core_252;
  assign popcount39_ub2f_core_293 = popcount39_ub2f_core_148 & popcount39_ub2f_core_252;
  assign popcount39_ub2f_core_294 = popcount39_ub2f_core_292 ^ popcount39_ub2f_core_288;
  assign popcount39_ub2f_core_295 = popcount39_ub2f_core_292 & popcount39_ub2f_core_288;
  assign popcount39_ub2f_core_296 = popcount39_ub2f_core_293 | popcount39_ub2f_core_295;
  assign popcount39_ub2f_core_299 = popcount39_ub2f_core_153 ^ popcount39_ub2f_core_296;
  assign popcount39_ub2f_core_300 = popcount39_ub2f_core_153 & popcount39_ub2f_core_296;
  assign popcount39_ub2f_core_304 = popcount39_ub2f_core_154 | popcount39_ub2f_core_300;
  assign popcount39_ub2f_core_305 = ~input_a[31];
  assign popcount39_ub2f_core_306 = input_a[28] ^ input_a[12];

  assign popcount39_ub2f_out[0] = 1'b0;
  assign popcount39_ub2f_out[1] = 1'b0;
  assign popcount39_ub2f_out[2] = popcount39_ub2f_core_287;
  assign popcount39_ub2f_out[3] = popcount39_ub2f_core_294;
  assign popcount39_ub2f_out[4] = popcount39_ub2f_core_299;
  assign popcount39_ub2f_out[5] = popcount39_ub2f_core_304;
endmodule