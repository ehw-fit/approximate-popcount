// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5291
// WCE=44.0
// EP=0.990669%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_mlfx(input [37:0] input_a, output [5:0] popcount38_mlfx_out);
  wire popcount38_mlfx_core_042;
  wire popcount38_mlfx_core_046;
  wire popcount38_mlfx_core_048;
  wire popcount38_mlfx_core_050;
  wire popcount38_mlfx_core_051;
  wire popcount38_mlfx_core_054;
  wire popcount38_mlfx_core_055;
  wire popcount38_mlfx_core_056;
  wire popcount38_mlfx_core_058;
  wire popcount38_mlfx_core_062;
  wire popcount38_mlfx_core_065;
  wire popcount38_mlfx_core_066;
  wire popcount38_mlfx_core_068;
  wire popcount38_mlfx_core_069;
  wire popcount38_mlfx_core_070;
  wire popcount38_mlfx_core_071;
  wire popcount38_mlfx_core_072;
  wire popcount38_mlfx_core_073;
  wire popcount38_mlfx_core_074;
  wire popcount38_mlfx_core_076;
  wire popcount38_mlfx_core_079;
  wire popcount38_mlfx_core_080;
  wire popcount38_mlfx_core_082;
  wire popcount38_mlfx_core_083;
  wire popcount38_mlfx_core_084;
  wire popcount38_mlfx_core_085;
  wire popcount38_mlfx_core_088;
  wire popcount38_mlfx_core_089;
  wire popcount38_mlfx_core_091;
  wire popcount38_mlfx_core_092;
  wire popcount38_mlfx_core_094;
  wire popcount38_mlfx_core_095;
  wire popcount38_mlfx_core_096;
  wire popcount38_mlfx_core_097;
  wire popcount38_mlfx_core_098;
  wire popcount38_mlfx_core_100;
  wire popcount38_mlfx_core_101;
  wire popcount38_mlfx_core_104;
  wire popcount38_mlfx_core_105;
  wire popcount38_mlfx_core_107;
  wire popcount38_mlfx_core_108;
  wire popcount38_mlfx_core_109;
  wire popcount38_mlfx_core_111;
  wire popcount38_mlfx_core_112;
  wire popcount38_mlfx_core_113;
  wire popcount38_mlfx_core_114;
  wire popcount38_mlfx_core_115;
  wire popcount38_mlfx_core_116;
  wire popcount38_mlfx_core_117;
  wire popcount38_mlfx_core_118;
  wire popcount38_mlfx_core_119;
  wire popcount38_mlfx_core_120;
  wire popcount38_mlfx_core_122;
  wire popcount38_mlfx_core_125;
  wire popcount38_mlfx_core_126;
  wire popcount38_mlfx_core_128;
  wire popcount38_mlfx_core_129;
  wire popcount38_mlfx_core_130;
  wire popcount38_mlfx_core_131;
  wire popcount38_mlfx_core_132;
  wire popcount38_mlfx_core_133;
  wire popcount38_mlfx_core_135;
  wire popcount38_mlfx_core_137;
  wire popcount38_mlfx_core_138;
  wire popcount38_mlfx_core_139;
  wire popcount38_mlfx_core_141;
  wire popcount38_mlfx_core_142;
  wire popcount38_mlfx_core_143;
  wire popcount38_mlfx_core_144;
  wire popcount38_mlfx_core_145;
  wire popcount38_mlfx_core_146;
  wire popcount38_mlfx_core_147;
  wire popcount38_mlfx_core_148;
  wire popcount38_mlfx_core_149;
  wire popcount38_mlfx_core_150;
  wire popcount38_mlfx_core_151;
  wire popcount38_mlfx_core_152;
  wire popcount38_mlfx_core_155;
  wire popcount38_mlfx_core_156;
  wire popcount38_mlfx_core_157;
  wire popcount38_mlfx_core_158;
  wire popcount38_mlfx_core_162;
  wire popcount38_mlfx_core_163;
  wire popcount38_mlfx_core_165;
  wire popcount38_mlfx_core_166;
  wire popcount38_mlfx_core_167;
  wire popcount38_mlfx_core_169;
  wire popcount38_mlfx_core_175;
  wire popcount38_mlfx_core_176;
  wire popcount38_mlfx_core_180;
  wire popcount38_mlfx_core_183;
  wire popcount38_mlfx_core_184;
  wire popcount38_mlfx_core_185;
  wire popcount38_mlfx_core_186;
  wire popcount38_mlfx_core_188;
  wire popcount38_mlfx_core_189;
  wire popcount38_mlfx_core_190;
  wire popcount38_mlfx_core_193;
  wire popcount38_mlfx_core_194;
  wire popcount38_mlfx_core_196;
  wire popcount38_mlfx_core_197;
  wire popcount38_mlfx_core_198;
  wire popcount38_mlfx_core_199;
  wire popcount38_mlfx_core_200;
  wire popcount38_mlfx_core_203;
  wire popcount38_mlfx_core_204;
  wire popcount38_mlfx_core_205;
  wire popcount38_mlfx_core_206;
  wire popcount38_mlfx_core_207;
  wire popcount38_mlfx_core_208;
  wire popcount38_mlfx_core_210;
  wire popcount38_mlfx_core_215;
  wire popcount38_mlfx_core_216;
  wire popcount38_mlfx_core_218;
  wire popcount38_mlfx_core_219;
  wire popcount38_mlfx_core_220;
  wire popcount38_mlfx_core_221;
  wire popcount38_mlfx_core_222;
  wire popcount38_mlfx_core_223;
  wire popcount38_mlfx_core_226;
  wire popcount38_mlfx_core_228;
  wire popcount38_mlfx_core_231;
  wire popcount38_mlfx_core_232;
  wire popcount38_mlfx_core_233;
  wire popcount38_mlfx_core_234;
  wire popcount38_mlfx_core_235;
  wire popcount38_mlfx_core_236;
  wire popcount38_mlfx_core_237;
  wire popcount38_mlfx_core_239;
  wire popcount38_mlfx_core_240;
  wire popcount38_mlfx_core_241;
  wire popcount38_mlfx_core_242;
  wire popcount38_mlfx_core_245;
  wire popcount38_mlfx_core_246;
  wire popcount38_mlfx_core_247;
  wire popcount38_mlfx_core_248;
  wire popcount38_mlfx_core_250;
  wire popcount38_mlfx_core_252;
  wire popcount38_mlfx_core_253;
  wire popcount38_mlfx_core_255;
  wire popcount38_mlfx_core_258;
  wire popcount38_mlfx_core_259;
  wire popcount38_mlfx_core_260;
  wire popcount38_mlfx_core_263;
  wire popcount38_mlfx_core_266;
  wire popcount38_mlfx_core_267;
  wire popcount38_mlfx_core_268;
  wire popcount38_mlfx_core_269;
  wire popcount38_mlfx_core_270;
  wire popcount38_mlfx_core_271;
  wire popcount38_mlfx_core_272;
  wire popcount38_mlfx_core_275;
  wire popcount38_mlfx_core_277;
  wire popcount38_mlfx_core_279;
  wire popcount38_mlfx_core_280;
  wire popcount38_mlfx_core_281;
  wire popcount38_mlfx_core_282;
  wire popcount38_mlfx_core_285;
  wire popcount38_mlfx_core_286;
  wire popcount38_mlfx_core_287;
  wire popcount38_mlfx_core_290;
  wire popcount38_mlfx_core_293;
  wire popcount38_mlfx_core_294;

  assign popcount38_mlfx_core_042 = input_a[20] & input_a[9];
  assign popcount38_mlfx_core_046 = input_a[26] | input_a[19];
  assign popcount38_mlfx_core_048 = input_a[27] | input_a[31];
  assign popcount38_mlfx_core_050 = ~input_a[1];
  assign popcount38_mlfx_core_051 = ~(input_a[15] & input_a[23]);
  assign popcount38_mlfx_core_054 = ~(input_a[31] | input_a[21]);
  assign popcount38_mlfx_core_055 = ~(input_a[19] | input_a[3]);
  assign popcount38_mlfx_core_056 = ~(input_a[1] ^ input_a[4]);
  assign popcount38_mlfx_core_058 = ~(input_a[3] ^ input_a[21]);
  assign popcount38_mlfx_core_062 = ~input_a[28];
  assign popcount38_mlfx_core_065 = ~input_a[22];
  assign popcount38_mlfx_core_066 = ~(input_a[37] ^ input_a[33]);
  assign popcount38_mlfx_core_068 = input_a[6] | input_a[32];
  assign popcount38_mlfx_core_069 = ~(input_a[6] | input_a[8]);
  assign popcount38_mlfx_core_070 = ~(input_a[0] | input_a[10]);
  assign popcount38_mlfx_core_071 = ~(input_a[28] ^ input_a[10]);
  assign popcount38_mlfx_core_072 = input_a[3] ^ input_a[37];
  assign popcount38_mlfx_core_073 = ~(input_a[33] & input_a[15]);
  assign popcount38_mlfx_core_074 = input_a[35] | input_a[22];
  assign popcount38_mlfx_core_076 = input_a[0] | input_a[22];
  assign popcount38_mlfx_core_079 = ~(input_a[32] ^ input_a[10]);
  assign popcount38_mlfx_core_080 = ~(input_a[31] | input_a[20]);
  assign popcount38_mlfx_core_082 = ~(input_a[8] & input_a[33]);
  assign popcount38_mlfx_core_083 = ~input_a[4];
  assign popcount38_mlfx_core_084 = ~(input_a[23] ^ input_a[11]);
  assign popcount38_mlfx_core_085 = input_a[2] ^ input_a[12];
  assign popcount38_mlfx_core_088 = input_a[36] ^ input_a[3];
  assign popcount38_mlfx_core_089 = input_a[13] & input_a[37];
  assign popcount38_mlfx_core_091 = input_a[30] & input_a[10];
  assign popcount38_mlfx_core_092 = ~(input_a[5] | input_a[37]);
  assign popcount38_mlfx_core_094 = ~(input_a[22] | input_a[34]);
  assign popcount38_mlfx_core_095 = ~input_a[21];
  assign popcount38_mlfx_core_096 = ~(input_a[33] & input_a[28]);
  assign popcount38_mlfx_core_097 = ~input_a[28];
  assign popcount38_mlfx_core_098 = ~(input_a[3] & input_a[35]);
  assign popcount38_mlfx_core_100 = input_a[24] | input_a[27];
  assign popcount38_mlfx_core_101 = input_a[17] ^ input_a[15];
  assign popcount38_mlfx_core_104 = ~(input_a[26] & input_a[22]);
  assign popcount38_mlfx_core_105 = ~(input_a[26] | input_a[9]);
  assign popcount38_mlfx_core_107 = input_a[20] ^ input_a[30];
  assign popcount38_mlfx_core_108 = input_a[35] ^ input_a[22];
  assign popcount38_mlfx_core_109 = input_a[13] & input_a[4];
  assign popcount38_mlfx_core_111 = ~(input_a[32] ^ input_a[25]);
  assign popcount38_mlfx_core_112 = ~(input_a[18] ^ input_a[35]);
  assign popcount38_mlfx_core_113 = ~input_a[33];
  assign popcount38_mlfx_core_114 = input_a[14] ^ input_a[1];
  assign popcount38_mlfx_core_115 = ~input_a[27];
  assign popcount38_mlfx_core_116 = ~(input_a[19] | input_a[35]);
  assign popcount38_mlfx_core_117 = input_a[10] | input_a[20];
  assign popcount38_mlfx_core_118 = ~(input_a[23] & input_a[15]);
  assign popcount38_mlfx_core_119 = input_a[30] & input_a[4];
  assign popcount38_mlfx_core_120 = input_a[29] & input_a[12];
  assign popcount38_mlfx_core_122 = input_a[26] ^ input_a[35];
  assign popcount38_mlfx_core_125 = input_a[37] ^ input_a[21];
  assign popcount38_mlfx_core_126 = ~(input_a[13] ^ input_a[35]);
  assign popcount38_mlfx_core_128 = ~(input_a[28] & input_a[8]);
  assign popcount38_mlfx_core_129 = ~(input_a[30] | input_a[12]);
  assign popcount38_mlfx_core_130 = input_a[21] ^ input_a[16];
  assign popcount38_mlfx_core_131 = input_a[12] ^ input_a[37];
  assign popcount38_mlfx_core_132 = ~input_a[18];
  assign popcount38_mlfx_core_133 = ~input_a[30];
  assign popcount38_mlfx_core_135 = input_a[3] | input_a[34];
  assign popcount38_mlfx_core_137 = ~(input_a[7] & input_a[16]);
  assign popcount38_mlfx_core_138 = ~input_a[34];
  assign popcount38_mlfx_core_139 = input_a[10] | input_a[28];
  assign popcount38_mlfx_core_141 = input_a[32] | input_a[35];
  assign popcount38_mlfx_core_142 = input_a[33] & input_a[30];
  assign popcount38_mlfx_core_143 = input_a[10] & input_a[23];
  assign popcount38_mlfx_core_144 = ~input_a[25];
  assign popcount38_mlfx_core_145 = input_a[28] & input_a[28];
  assign popcount38_mlfx_core_146 = input_a[20] | input_a[4];
  assign popcount38_mlfx_core_147 = ~(input_a[31] & input_a[0]);
  assign popcount38_mlfx_core_148 = input_a[3] | input_a[13];
  assign popcount38_mlfx_core_149 = ~(input_a[31] ^ input_a[33]);
  assign popcount38_mlfx_core_150 = ~(input_a[35] | input_a[21]);
  assign popcount38_mlfx_core_151 = input_a[37] & input_a[23];
  assign popcount38_mlfx_core_152 = ~(input_a[16] ^ input_a[21]);
  assign popcount38_mlfx_core_155 = input_a[21] | input_a[15];
  assign popcount38_mlfx_core_156 = ~input_a[34];
  assign popcount38_mlfx_core_157 = input_a[33] & input_a[32];
  assign popcount38_mlfx_core_158 = ~input_a[33];
  assign popcount38_mlfx_core_162 = ~(input_a[14] | input_a[37]);
  assign popcount38_mlfx_core_163 = input_a[30] ^ input_a[26];
  assign popcount38_mlfx_core_165 = input_a[23] ^ input_a[31];
  assign popcount38_mlfx_core_166 = ~(input_a[35] | input_a[25]);
  assign popcount38_mlfx_core_167 = input_a[30] & input_a[12];
  assign popcount38_mlfx_core_169 = input_a[0] ^ input_a[14];
  assign popcount38_mlfx_core_175 = ~(input_a[2] ^ input_a[7]);
  assign popcount38_mlfx_core_176 = input_a[2] ^ input_a[35];
  assign popcount38_mlfx_core_180 = input_a[12] ^ input_a[17];
  assign popcount38_mlfx_core_183 = ~(input_a[31] ^ input_a[6]);
  assign popcount38_mlfx_core_184 = ~(input_a[8] ^ input_a[20]);
  assign popcount38_mlfx_core_185 = ~(input_a[8] ^ input_a[14]);
  assign popcount38_mlfx_core_186 = input_a[31] | input_a[19];
  assign popcount38_mlfx_core_188 = ~(input_a[33] ^ input_a[13]);
  assign popcount38_mlfx_core_189 = ~(input_a[4] ^ input_a[7]);
  assign popcount38_mlfx_core_190 = input_a[16] ^ input_a[14];
  assign popcount38_mlfx_core_193 = input_a[1] ^ input_a[6];
  assign popcount38_mlfx_core_194 = ~(input_a[35] & input_a[24]);
  assign popcount38_mlfx_core_196 = ~input_a[26];
  assign popcount38_mlfx_core_197 = ~(input_a[0] ^ input_a[31]);
  assign popcount38_mlfx_core_198 = ~(input_a[19] ^ input_a[7]);
  assign popcount38_mlfx_core_199 = ~(input_a[35] | input_a[6]);
  assign popcount38_mlfx_core_200 = ~(input_a[8] & input_a[17]);
  assign popcount38_mlfx_core_203 = input_a[36] ^ input_a[26];
  assign popcount38_mlfx_core_204 = ~(input_a[4] | input_a[5]);
  assign popcount38_mlfx_core_205 = input_a[18] & input_a[24];
  assign popcount38_mlfx_core_206 = input_a[29] ^ input_a[33];
  assign popcount38_mlfx_core_207 = ~(input_a[8] & input_a[8]);
  assign popcount38_mlfx_core_208 = input_a[25] | input_a[12];
  assign popcount38_mlfx_core_210 = ~(input_a[30] & input_a[0]);
  assign popcount38_mlfx_core_215 = ~(input_a[33] & input_a[3]);
  assign popcount38_mlfx_core_216 = ~(input_a[22] & input_a[4]);
  assign popcount38_mlfx_core_218 = input_a[8] | input_a[28];
  assign popcount38_mlfx_core_219 = ~input_a[1];
  assign popcount38_mlfx_core_220 = input_a[6] ^ input_a[32];
  assign popcount38_mlfx_core_221 = ~(input_a[28] ^ input_a[32]);
  assign popcount38_mlfx_core_222 = ~input_a[33];
  assign popcount38_mlfx_core_223 = ~(input_a[19] | input_a[36]);
  assign popcount38_mlfx_core_226 = input_a[35] | input_a[20];
  assign popcount38_mlfx_core_228 = input_a[29] | input_a[20];
  assign popcount38_mlfx_core_231 = ~input_a[32];
  assign popcount38_mlfx_core_232 = ~input_a[0];
  assign popcount38_mlfx_core_233 = ~input_a[1];
  assign popcount38_mlfx_core_234 = input_a[8] & input_a[20];
  assign popcount38_mlfx_core_235 = ~(input_a[2] & input_a[20]);
  assign popcount38_mlfx_core_236 = input_a[24] & input_a[29];
  assign popcount38_mlfx_core_237 = ~(input_a[9] ^ input_a[35]);
  assign popcount38_mlfx_core_239 = ~input_a[21];
  assign popcount38_mlfx_core_240 = input_a[7] & input_a[34];
  assign popcount38_mlfx_core_241 = ~(input_a[10] | input_a[28]);
  assign popcount38_mlfx_core_242 = ~(input_a[12] & input_a[3]);
  assign popcount38_mlfx_core_245 = ~input_a[7];
  assign popcount38_mlfx_core_246 = ~(input_a[32] | input_a[31]);
  assign popcount38_mlfx_core_247 = input_a[37] ^ input_a[37];
  assign popcount38_mlfx_core_248 = input_a[6] | input_a[6];
  assign popcount38_mlfx_core_250 = ~(input_a[7] | input_a[34]);
  assign popcount38_mlfx_core_252 = input_a[9] | input_a[3];
  assign popcount38_mlfx_core_253 = ~input_a[8];
  assign popcount38_mlfx_core_255 = input_a[9] | input_a[32];
  assign popcount38_mlfx_core_258 = ~(input_a[34] & input_a[28]);
  assign popcount38_mlfx_core_259 = ~(input_a[9] ^ input_a[34]);
  assign popcount38_mlfx_core_260 = ~(input_a[23] ^ input_a[12]);
  assign popcount38_mlfx_core_263 = ~input_a[4];
  assign popcount38_mlfx_core_266 = ~(input_a[24] & input_a[31]);
  assign popcount38_mlfx_core_267 = ~input_a[33];
  assign popcount38_mlfx_core_268 = ~(input_a[29] | input_a[18]);
  assign popcount38_mlfx_core_269 = input_a[34] & input_a[0];
  assign popcount38_mlfx_core_270 = input_a[17] & input_a[11];
  assign popcount38_mlfx_core_271 = ~(input_a[15] | input_a[21]);
  assign popcount38_mlfx_core_272 = ~(input_a[19] & input_a[33]);
  assign popcount38_mlfx_core_275 = ~input_a[35];
  assign popcount38_mlfx_core_277 = ~input_a[31];
  assign popcount38_mlfx_core_279 = ~(input_a[27] ^ input_a[28]);
  assign popcount38_mlfx_core_280 = ~(input_a[1] ^ input_a[32]);
  assign popcount38_mlfx_core_281 = ~(input_a[9] ^ input_a[32]);
  assign popcount38_mlfx_core_282 = ~(input_a[18] | input_a[26]);
  assign popcount38_mlfx_core_285 = input_a[13] | input_a[31];
  assign popcount38_mlfx_core_286 = ~input_a[30];
  assign popcount38_mlfx_core_287 = ~(input_a[25] ^ input_a[22]);
  assign popcount38_mlfx_core_290 = ~(input_a[31] & input_a[35]);
  assign popcount38_mlfx_core_293 = ~(input_a[35] | input_a[36]);
  assign popcount38_mlfx_core_294 = ~(input_a[22] | input_a[32]);

  assign popcount38_mlfx_out[0] = 1'b1;
  assign popcount38_mlfx_out[1] = input_a[28];
  assign popcount38_mlfx_out[2] = input_a[3];
  assign popcount38_mlfx_out[3] = 1'b1;
  assign popcount38_mlfx_out[4] = 1'b0;
  assign popcount38_mlfx_out[5] = input_a[7];
endmodule