// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.23047
// WCE=5.0
// EP=0.753906%
// Printed PDK parameters:
//  Area=38666644.0
//  Delay=57841800.0
//  Power=1944100.0

module popcount25_n4rw(input [24:0] input_a, output [4:0] popcount25_n4rw_out);
  wire popcount25_n4rw_core_027;
  wire popcount25_n4rw_core_028;
  wire popcount25_n4rw_core_030;
  wire popcount25_n4rw_core_031;
  wire popcount25_n4rw_core_032;
  wire popcount25_n4rw_core_034;
  wire popcount25_n4rw_core_038;
  wire popcount25_n4rw_core_039;
  wire popcount25_n4rw_core_040;
  wire popcount25_n4rw_core_041;
  wire popcount25_n4rw_core_042;
  wire popcount25_n4rw_core_044;
  wire popcount25_n4rw_core_047;
  wire popcount25_n4rw_core_048;
  wire popcount25_n4rw_core_050;
  wire popcount25_n4rw_core_051;
  wire popcount25_n4rw_core_052;
  wire popcount25_n4rw_core_053;
  wire popcount25_n4rw_core_054;
  wire popcount25_n4rw_core_055;
  wire popcount25_n4rw_core_057;
  wire popcount25_n4rw_core_058;
  wire popcount25_n4rw_core_060;
  wire popcount25_n4rw_core_061;
  wire popcount25_n4rw_core_062;
  wire popcount25_n4rw_core_064;
  wire popcount25_n4rw_core_065;
  wire popcount25_n4rw_core_066;
  wire popcount25_n4rw_core_067;
  wire popcount25_n4rw_core_068;
  wire popcount25_n4rw_core_069;
  wire popcount25_n4rw_core_071;
  wire popcount25_n4rw_core_073;
  wire popcount25_n4rw_core_077;
  wire popcount25_n4rw_core_078;
  wire popcount25_n4rw_core_080;
  wire popcount25_n4rw_core_082;
  wire popcount25_n4rw_core_083;
  wire popcount25_n4rw_core_084;
  wire popcount25_n4rw_core_085;
  wire popcount25_n4rw_core_086;
  wire popcount25_n4rw_core_088;
  wire popcount25_n4rw_core_091;
  wire popcount25_n4rw_core_092;
  wire popcount25_n4rw_core_093;
  wire popcount25_n4rw_core_094;
  wire popcount25_n4rw_core_095;
  wire popcount25_n4rw_core_096;
  wire popcount25_n4rw_core_097;
  wire popcount25_n4rw_core_098;
  wire popcount25_n4rw_core_099;
  wire popcount25_n4rw_core_100;
  wire popcount25_n4rw_core_101;
  wire popcount25_n4rw_core_102;
  wire popcount25_n4rw_core_104;
  wire popcount25_n4rw_core_105;
  wire popcount25_n4rw_core_106;
  wire popcount25_n4rw_core_107;
  wire popcount25_n4rw_core_108;
  wire popcount25_n4rw_core_109;
  wire popcount25_n4rw_core_110;
  wire popcount25_n4rw_core_112;
  wire popcount25_n4rw_core_114;
  wire popcount25_n4rw_core_115;
  wire popcount25_n4rw_core_116;
  wire popcount25_n4rw_core_117;
  wire popcount25_n4rw_core_118_not;
  wire popcount25_n4rw_core_119;
  wire popcount25_n4rw_core_121;
  wire popcount25_n4rw_core_123;
  wire popcount25_n4rw_core_124;
  wire popcount25_n4rw_core_125;
  wire popcount25_n4rw_core_126;
  wire popcount25_n4rw_core_129;
  wire popcount25_n4rw_core_130;
  wire popcount25_n4rw_core_132;
  wire popcount25_n4rw_core_134;
  wire popcount25_n4rw_core_136;
  wire popcount25_n4rw_core_138;
  wire popcount25_n4rw_core_139;
  wire popcount25_n4rw_core_140;
  wire popcount25_n4rw_core_141;
  wire popcount25_n4rw_core_143;
  wire popcount25_n4rw_core_144;
  wire popcount25_n4rw_core_145;
  wire popcount25_n4rw_core_147;
  wire popcount25_n4rw_core_148;
  wire popcount25_n4rw_core_150;
  wire popcount25_n4rw_core_152;
  wire popcount25_n4rw_core_154;
  wire popcount25_n4rw_core_155;
  wire popcount25_n4rw_core_156;
  wire popcount25_n4rw_core_162;
  wire popcount25_n4rw_core_163;
  wire popcount25_n4rw_core_164;
  wire popcount25_n4rw_core_165;
  wire popcount25_n4rw_core_166;
  wire popcount25_n4rw_core_167;
  wire popcount25_n4rw_core_168;
  wire popcount25_n4rw_core_169;
  wire popcount25_n4rw_core_170;
  wire popcount25_n4rw_core_171;
  wire popcount25_n4rw_core_172;
  wire popcount25_n4rw_core_173;
  wire popcount25_n4rw_core_174;
  wire popcount25_n4rw_core_175;
  wire popcount25_n4rw_core_176;
  wire popcount25_n4rw_core_177;
  wire popcount25_n4rw_core_178;
  wire popcount25_n4rw_core_179;
  wire popcount25_n4rw_core_181;
  wire popcount25_n4rw_core_183;

  assign popcount25_n4rw_core_027 = input_a[19] ^ input_a[21];
  assign popcount25_n4rw_core_028 = input_a[1] & input_a[2];
  assign popcount25_n4rw_core_030 = input_a[0] & input_a[13];
  assign popcount25_n4rw_core_031 = popcount25_n4rw_core_028 ^ popcount25_n4rw_core_030;
  assign popcount25_n4rw_core_032 = popcount25_n4rw_core_028 & popcount25_n4rw_core_030;
  assign popcount25_n4rw_core_034 = input_a[4] & input_a[5];
  assign popcount25_n4rw_core_038 = input_a[12] ^ input_a[13];
  assign popcount25_n4rw_core_039 = input_a[24] ^ input_a[15];
  assign popcount25_n4rw_core_040 = ~(input_a[24] ^ input_a[8]);
  assign popcount25_n4rw_core_041 = popcount25_n4rw_core_031 ^ popcount25_n4rw_core_034;
  assign popcount25_n4rw_core_042 = popcount25_n4rw_core_031 & popcount25_n4rw_core_034;
  assign popcount25_n4rw_core_044 = input_a[12] | input_a[14];
  assign popcount25_n4rw_core_047 = ~(input_a[0] | input_a[20]);
  assign popcount25_n4rw_core_048 = popcount25_n4rw_core_032 | popcount25_n4rw_core_042;
  assign popcount25_n4rw_core_050 = ~(input_a[3] | input_a[6]);
  assign popcount25_n4rw_core_051 = input_a[7] | input_a[8];
  assign popcount25_n4rw_core_052 = input_a[7] & input_a[8];
  assign popcount25_n4rw_core_053 = ~input_a[3];
  assign popcount25_n4rw_core_054 = input_a[6] & popcount25_n4rw_core_051;
  assign popcount25_n4rw_core_055 = popcount25_n4rw_core_052 | popcount25_n4rw_core_054;
  assign popcount25_n4rw_core_057 = input_a[10] | input_a[11];
  assign popcount25_n4rw_core_058 = input_a[10] & input_a[11];
  assign popcount25_n4rw_core_060 = input_a[9] & popcount25_n4rw_core_057;
  assign popcount25_n4rw_core_061 = popcount25_n4rw_core_058 | popcount25_n4rw_core_060;
  assign popcount25_n4rw_core_062 = ~(input_a[11] & input_a[21]);
  assign popcount25_n4rw_core_064 = input_a[22] & input_a[3];
  assign popcount25_n4rw_core_065 = popcount25_n4rw_core_055 ^ popcount25_n4rw_core_061;
  assign popcount25_n4rw_core_066 = popcount25_n4rw_core_055 & popcount25_n4rw_core_061;
  assign popcount25_n4rw_core_067 = popcount25_n4rw_core_065 ^ popcount25_n4rw_core_064;
  assign popcount25_n4rw_core_068 = popcount25_n4rw_core_065 & popcount25_n4rw_core_064;
  assign popcount25_n4rw_core_069 = popcount25_n4rw_core_066 | popcount25_n4rw_core_068;
  assign popcount25_n4rw_core_071 = input_a[21] | input_a[2];
  assign popcount25_n4rw_core_073 = input_a[22] ^ input_a[12];
  assign popcount25_n4rw_core_077 = popcount25_n4rw_core_041 ^ popcount25_n4rw_core_067;
  assign popcount25_n4rw_core_078 = popcount25_n4rw_core_041 & popcount25_n4rw_core_067;
  assign popcount25_n4rw_core_080 = ~input_a[14];
  assign popcount25_n4rw_core_082 = popcount25_n4rw_core_048 ^ popcount25_n4rw_core_069;
  assign popcount25_n4rw_core_083 = popcount25_n4rw_core_048 & popcount25_n4rw_core_069;
  assign popcount25_n4rw_core_084 = popcount25_n4rw_core_082 ^ popcount25_n4rw_core_078;
  assign popcount25_n4rw_core_085 = popcount25_n4rw_core_082 & popcount25_n4rw_core_078;
  assign popcount25_n4rw_core_086 = popcount25_n4rw_core_083 | popcount25_n4rw_core_085;
  assign popcount25_n4rw_core_088 = ~input_a[22];
  assign popcount25_n4rw_core_091 = input_a[7] & input_a[24];
  assign popcount25_n4rw_core_092 = ~(input_a[18] & input_a[2]);
  assign popcount25_n4rw_core_093 = input_a[21] & input_a[14];
  assign popcount25_n4rw_core_094 = ~(input_a[13] | input_a[13]);
  assign popcount25_n4rw_core_095 = input_a[12] & input_a[24];
  assign popcount25_n4rw_core_096 = popcount25_n4rw_core_093 | popcount25_n4rw_core_095;
  assign popcount25_n4rw_core_097 = ~(input_a[17] | input_a[11]);
  assign popcount25_n4rw_core_098 = input_a[16] ^ input_a[17];
  assign popcount25_n4rw_core_099 = input_a[16] & input_a[17];
  assign popcount25_n4rw_core_100 = input_a[15] ^ popcount25_n4rw_core_098;
  assign popcount25_n4rw_core_101 = input_a[15] & popcount25_n4rw_core_098;
  assign popcount25_n4rw_core_102 = popcount25_n4rw_core_099 | popcount25_n4rw_core_101;
  assign popcount25_n4rw_core_104 = input_a[4] ^ input_a[17];
  assign popcount25_n4rw_core_105 = input_a[20] & popcount25_n4rw_core_100;
  assign popcount25_n4rw_core_106 = popcount25_n4rw_core_096 ^ popcount25_n4rw_core_102;
  assign popcount25_n4rw_core_107 = popcount25_n4rw_core_096 & popcount25_n4rw_core_102;
  assign popcount25_n4rw_core_108 = popcount25_n4rw_core_106 ^ popcount25_n4rw_core_105;
  assign popcount25_n4rw_core_109 = popcount25_n4rw_core_106 & popcount25_n4rw_core_105;
  assign popcount25_n4rw_core_110 = popcount25_n4rw_core_107 | popcount25_n4rw_core_109;
  assign popcount25_n4rw_core_112 = ~(input_a[0] & input_a[11]);
  assign popcount25_n4rw_core_114 = input_a[9] ^ input_a[2];
  assign popcount25_n4rw_core_115 = input_a[6] ^ input_a[14];
  assign popcount25_n4rw_core_116 = ~input_a[22];
  assign popcount25_n4rw_core_117 = input_a[19] & input_a[23];
  assign popcount25_n4rw_core_118_not = ~input_a[8];
  assign popcount25_n4rw_core_119 = ~input_a[1];
  assign popcount25_n4rw_core_121 = input_a[11] ^ input_a[8];
  assign popcount25_n4rw_core_123 = ~(input_a[10] | input_a[17]);
  assign popcount25_n4rw_core_124 = ~(input_a[16] & input_a[11]);
  assign popcount25_n4rw_core_125 = ~(input_a[18] & input_a[11]);
  assign popcount25_n4rw_core_126 = ~(input_a[20] ^ input_a[8]);
  assign popcount25_n4rw_core_129 = ~input_a[16];
  assign popcount25_n4rw_core_130 = ~(input_a[4] ^ input_a[18]);
  assign popcount25_n4rw_core_132 = input_a[19] & input_a[14];
  assign popcount25_n4rw_core_134 = ~(input_a[16] | input_a[6]);
  assign popcount25_n4rw_core_136 = input_a[16] ^ input_a[9];
  assign popcount25_n4rw_core_138 = input_a[20] & input_a[3];
  assign popcount25_n4rw_core_139 = ~(input_a[5] & input_a[11]);
  assign popcount25_n4rw_core_140 = input_a[21] & input_a[11];
  assign popcount25_n4rw_core_141 = input_a[15] & input_a[17];
  assign popcount25_n4rw_core_143 = ~(input_a[5] ^ input_a[13]);
  assign popcount25_n4rw_core_144 = input_a[16] & input_a[1];
  assign popcount25_n4rw_core_145 = ~(input_a[14] | input_a[19]);
  assign popcount25_n4rw_core_147 = popcount25_n4rw_core_108 ^ popcount25_n4rw_core_117;
  assign popcount25_n4rw_core_148 = popcount25_n4rw_core_108 & popcount25_n4rw_core_117;
  assign popcount25_n4rw_core_150 = input_a[4] ^ input_a[9];
  assign popcount25_n4rw_core_152 = ~popcount25_n4rw_core_110;
  assign popcount25_n4rw_core_154 = popcount25_n4rw_core_152 ^ popcount25_n4rw_core_148;
  assign popcount25_n4rw_core_155 = input_a[19] & popcount25_n4rw_core_148;
  assign popcount25_n4rw_core_156 = popcount25_n4rw_core_110 | popcount25_n4rw_core_155;
  assign popcount25_n4rw_core_162 = ~input_a[18];
  assign popcount25_n4rw_core_163 = ~input_a[5];
  assign popcount25_n4rw_core_164 = popcount25_n4rw_core_077 ^ popcount25_n4rw_core_147;
  assign popcount25_n4rw_core_165 = popcount25_n4rw_core_077 & popcount25_n4rw_core_147;
  assign popcount25_n4rw_core_166 = popcount25_n4rw_core_164 ^ input_a[18];
  assign popcount25_n4rw_core_167 = popcount25_n4rw_core_164 & input_a[18];
  assign popcount25_n4rw_core_168 = popcount25_n4rw_core_165 | popcount25_n4rw_core_167;
  assign popcount25_n4rw_core_169 = popcount25_n4rw_core_084 ^ popcount25_n4rw_core_154;
  assign popcount25_n4rw_core_170 = popcount25_n4rw_core_084 & popcount25_n4rw_core_154;
  assign popcount25_n4rw_core_171 = popcount25_n4rw_core_169 ^ popcount25_n4rw_core_168;
  assign popcount25_n4rw_core_172 = popcount25_n4rw_core_169 & popcount25_n4rw_core_168;
  assign popcount25_n4rw_core_173 = popcount25_n4rw_core_170 | popcount25_n4rw_core_172;
  assign popcount25_n4rw_core_174 = popcount25_n4rw_core_086 ^ popcount25_n4rw_core_156;
  assign popcount25_n4rw_core_175 = popcount25_n4rw_core_086 & popcount25_n4rw_core_156;
  assign popcount25_n4rw_core_176 = popcount25_n4rw_core_174 ^ popcount25_n4rw_core_173;
  assign popcount25_n4rw_core_177 = popcount25_n4rw_core_174 & popcount25_n4rw_core_173;
  assign popcount25_n4rw_core_178 = popcount25_n4rw_core_175 | popcount25_n4rw_core_177;
  assign popcount25_n4rw_core_179 = ~(input_a[9] & input_a[8]);
  assign popcount25_n4rw_core_181 = input_a[18] | input_a[13];
  assign popcount25_n4rw_core_183 = input_a[17] ^ input_a[19];

  assign popcount25_n4rw_out[0] = popcount25_n4rw_core_162;
  assign popcount25_n4rw_out[1] = popcount25_n4rw_core_166;
  assign popcount25_n4rw_out[2] = popcount25_n4rw_core_171;
  assign popcount25_n4rw_out[3] = popcount25_n4rw_core_176;
  assign popcount25_n4rw_out[4] = popcount25_n4rw_core_178;
endmodule