// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.07994
// WCE=21.0
// EP=0.969959%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_6wfk(input [32:0] input_a, output [5:0] popcount33_6wfk_out);
  wire popcount33_6wfk_core_035;
  wire popcount33_6wfk_core_037;
  wire popcount33_6wfk_core_039;
  wire popcount33_6wfk_core_040;
  wire popcount33_6wfk_core_041;
  wire popcount33_6wfk_core_042_not;
  wire popcount33_6wfk_core_045;
  wire popcount33_6wfk_core_049;
  wire popcount33_6wfk_core_052;
  wire popcount33_6wfk_core_053;
  wire popcount33_6wfk_core_054;
  wire popcount33_6wfk_core_057;
  wire popcount33_6wfk_core_059;
  wire popcount33_6wfk_core_062;
  wire popcount33_6wfk_core_068;
  wire popcount33_6wfk_core_069;
  wire popcount33_6wfk_core_070;
  wire popcount33_6wfk_core_071;
  wire popcount33_6wfk_core_073;
  wire popcount33_6wfk_core_075;
  wire popcount33_6wfk_core_077;
  wire popcount33_6wfk_core_078;
  wire popcount33_6wfk_core_079;
  wire popcount33_6wfk_core_080;
  wire popcount33_6wfk_core_081;
  wire popcount33_6wfk_core_082;
  wire popcount33_6wfk_core_084;
  wire popcount33_6wfk_core_085;
  wire popcount33_6wfk_core_086;
  wire popcount33_6wfk_core_088;
  wire popcount33_6wfk_core_089;
  wire popcount33_6wfk_core_090;
  wire popcount33_6wfk_core_091;
  wire popcount33_6wfk_core_092;
  wire popcount33_6wfk_core_094;
  wire popcount33_6wfk_core_095;
  wire popcount33_6wfk_core_096;
  wire popcount33_6wfk_core_098;
  wire popcount33_6wfk_core_099;
  wire popcount33_6wfk_core_101;
  wire popcount33_6wfk_core_102;
  wire popcount33_6wfk_core_103;
  wire popcount33_6wfk_core_106;
  wire popcount33_6wfk_core_108;
  wire popcount33_6wfk_core_109;
  wire popcount33_6wfk_core_112;
  wire popcount33_6wfk_core_113;
  wire popcount33_6wfk_core_114;
  wire popcount33_6wfk_core_115;
  wire popcount33_6wfk_core_116;
  wire popcount33_6wfk_core_118;
  wire popcount33_6wfk_core_119;
  wire popcount33_6wfk_core_120;
  wire popcount33_6wfk_core_121;
  wire popcount33_6wfk_core_122;
  wire popcount33_6wfk_core_123;
  wire popcount33_6wfk_core_124;
  wire popcount33_6wfk_core_128;
  wire popcount33_6wfk_core_129;
  wire popcount33_6wfk_core_130;
  wire popcount33_6wfk_core_131;
  wire popcount33_6wfk_core_132;
  wire popcount33_6wfk_core_133;
  wire popcount33_6wfk_core_134;
  wire popcount33_6wfk_core_136;
  wire popcount33_6wfk_core_137;
  wire popcount33_6wfk_core_138;
  wire popcount33_6wfk_core_139;
  wire popcount33_6wfk_core_140;
  wire popcount33_6wfk_core_142;
  wire popcount33_6wfk_core_144;
  wire popcount33_6wfk_core_146;
  wire popcount33_6wfk_core_147;
  wire popcount33_6wfk_core_148;
  wire popcount33_6wfk_core_149;
  wire popcount33_6wfk_core_150;
  wire popcount33_6wfk_core_151;
  wire popcount33_6wfk_core_152;
  wire popcount33_6wfk_core_153;
  wire popcount33_6wfk_core_155;
  wire popcount33_6wfk_core_156;
  wire popcount33_6wfk_core_159;
  wire popcount33_6wfk_core_160_not;
  wire popcount33_6wfk_core_161;
  wire popcount33_6wfk_core_162;
  wire popcount33_6wfk_core_163;
  wire popcount33_6wfk_core_165;
  wire popcount33_6wfk_core_167;
  wire popcount33_6wfk_core_168;
  wire popcount33_6wfk_core_169;
  wire popcount33_6wfk_core_170;
  wire popcount33_6wfk_core_173;
  wire popcount33_6wfk_core_177;
  wire popcount33_6wfk_core_181;
  wire popcount33_6wfk_core_183;
  wire popcount33_6wfk_core_185;
  wire popcount33_6wfk_core_186;
  wire popcount33_6wfk_core_187;
  wire popcount33_6wfk_core_189;
  wire popcount33_6wfk_core_190;
  wire popcount33_6wfk_core_191;
  wire popcount33_6wfk_core_192;
  wire popcount33_6wfk_core_194;
  wire popcount33_6wfk_core_195;
  wire popcount33_6wfk_core_196_not;
  wire popcount33_6wfk_core_197;
  wire popcount33_6wfk_core_198;
  wire popcount33_6wfk_core_199;
  wire popcount33_6wfk_core_200;
  wire popcount33_6wfk_core_201;
  wire popcount33_6wfk_core_202;
  wire popcount33_6wfk_core_205;
  wire popcount33_6wfk_core_206;
  wire popcount33_6wfk_core_207;
  wire popcount33_6wfk_core_208;
  wire popcount33_6wfk_core_209;
  wire popcount33_6wfk_core_211;
  wire popcount33_6wfk_core_212;
  wire popcount33_6wfk_core_216;
  wire popcount33_6wfk_core_217;
  wire popcount33_6wfk_core_218;
  wire popcount33_6wfk_core_220;
  wire popcount33_6wfk_core_224;
  wire popcount33_6wfk_core_225;
  wire popcount33_6wfk_core_226;
  wire popcount33_6wfk_core_227;
  wire popcount33_6wfk_core_228;
  wire popcount33_6wfk_core_233;
  wire popcount33_6wfk_core_235;

  assign popcount33_6wfk_core_035 = input_a[28] & input_a[29];
  assign popcount33_6wfk_core_037 = ~(input_a[7] & input_a[29]);
  assign popcount33_6wfk_core_039 = ~input_a[28];
  assign popcount33_6wfk_core_040 = ~(input_a[6] | input_a[11]);
  assign popcount33_6wfk_core_041 = input_a[28] & input_a[14];
  assign popcount33_6wfk_core_042_not = ~input_a[8];
  assign popcount33_6wfk_core_045 = input_a[17] ^ input_a[7];
  assign popcount33_6wfk_core_049 = ~(input_a[18] | input_a[8]);
  assign popcount33_6wfk_core_052 = ~(input_a[2] ^ input_a[11]);
  assign popcount33_6wfk_core_053 = input_a[26] ^ input_a[0];
  assign popcount33_6wfk_core_054 = ~(input_a[4] ^ input_a[3]);
  assign popcount33_6wfk_core_057 = ~input_a[4];
  assign popcount33_6wfk_core_059 = ~(input_a[12] | input_a[32]);
  assign popcount33_6wfk_core_062 = input_a[0] | input_a[24];
  assign popcount33_6wfk_core_068 = input_a[10] | input_a[25];
  assign popcount33_6wfk_core_069 = ~(input_a[13] & input_a[15]);
  assign popcount33_6wfk_core_070 = ~input_a[3];
  assign popcount33_6wfk_core_071 = ~(input_a[20] ^ input_a[22]);
  assign popcount33_6wfk_core_073 = ~(input_a[30] & input_a[25]);
  assign popcount33_6wfk_core_075 = input_a[12] & input_a[18];
  assign popcount33_6wfk_core_077 = input_a[16] ^ input_a[22];
  assign popcount33_6wfk_core_078 = ~input_a[4];
  assign popcount33_6wfk_core_079 = ~input_a[5];
  assign popcount33_6wfk_core_080 = input_a[19] ^ input_a[1];
  assign popcount33_6wfk_core_081 = input_a[14] & input_a[9];
  assign popcount33_6wfk_core_082 = ~input_a[21];
  assign popcount33_6wfk_core_084 = ~(input_a[16] | input_a[30]);
  assign popcount33_6wfk_core_085 = input_a[3] & input_a[32];
  assign popcount33_6wfk_core_086 = ~input_a[6];
  assign popcount33_6wfk_core_088 = input_a[13] | input_a[28];
  assign popcount33_6wfk_core_089 = ~(input_a[10] ^ input_a[0]);
  assign popcount33_6wfk_core_090 = ~(input_a[9] ^ input_a[32]);
  assign popcount33_6wfk_core_091 = ~(input_a[11] | input_a[5]);
  assign popcount33_6wfk_core_092 = ~(input_a[1] & input_a[18]);
  assign popcount33_6wfk_core_094 = ~(input_a[26] ^ input_a[15]);
  assign popcount33_6wfk_core_095 = ~(input_a[15] | input_a[28]);
  assign popcount33_6wfk_core_096 = ~(input_a[11] & input_a[1]);
  assign popcount33_6wfk_core_098 = ~(input_a[19] | input_a[17]);
  assign popcount33_6wfk_core_099 = ~(input_a[30] & input_a[4]);
  assign popcount33_6wfk_core_101 = ~(input_a[3] ^ input_a[25]);
  assign popcount33_6wfk_core_102 = ~input_a[10];
  assign popcount33_6wfk_core_103 = input_a[7] | input_a[20];
  assign popcount33_6wfk_core_106 = ~(input_a[12] | input_a[14]);
  assign popcount33_6wfk_core_108 = input_a[22] | input_a[22];
  assign popcount33_6wfk_core_109 = input_a[26] & input_a[1];
  assign popcount33_6wfk_core_112 = ~(input_a[28] & input_a[12]);
  assign popcount33_6wfk_core_113 = ~(input_a[28] ^ input_a[20]);
  assign popcount33_6wfk_core_114 = ~(input_a[12] | input_a[4]);
  assign popcount33_6wfk_core_115 = input_a[19] ^ input_a[5];
  assign popcount33_6wfk_core_116 = input_a[28] ^ input_a[11];
  assign popcount33_6wfk_core_118 = input_a[18] & input_a[27];
  assign popcount33_6wfk_core_119 = ~(input_a[4] | input_a[18]);
  assign popcount33_6wfk_core_120 = ~(input_a[4] & input_a[1]);
  assign popcount33_6wfk_core_121 = ~(input_a[16] | input_a[30]);
  assign popcount33_6wfk_core_122 = input_a[0] ^ input_a[31];
  assign popcount33_6wfk_core_123 = input_a[18] | input_a[4];
  assign popcount33_6wfk_core_124 = ~(input_a[28] & input_a[5]);
  assign popcount33_6wfk_core_128 = ~input_a[14];
  assign popcount33_6wfk_core_129 = ~input_a[14];
  assign popcount33_6wfk_core_130 = input_a[1] | input_a[0];
  assign popcount33_6wfk_core_131 = ~(input_a[25] ^ input_a[24]);
  assign popcount33_6wfk_core_132 = ~(input_a[18] ^ input_a[11]);
  assign popcount33_6wfk_core_133 = ~input_a[30];
  assign popcount33_6wfk_core_134 = input_a[4] | input_a[18];
  assign popcount33_6wfk_core_136 = input_a[5] | input_a[30];
  assign popcount33_6wfk_core_137 = input_a[10] & input_a[15];
  assign popcount33_6wfk_core_138 = ~(input_a[27] ^ input_a[13]);
  assign popcount33_6wfk_core_139 = ~(input_a[19] | input_a[15]);
  assign popcount33_6wfk_core_140 = ~(input_a[5] ^ input_a[31]);
  assign popcount33_6wfk_core_142 = ~(input_a[10] & input_a[22]);
  assign popcount33_6wfk_core_144 = ~(input_a[5] ^ input_a[6]);
  assign popcount33_6wfk_core_146 = ~(input_a[23] | input_a[31]);
  assign popcount33_6wfk_core_147 = input_a[21] & input_a[4];
  assign popcount33_6wfk_core_148 = input_a[9] & input_a[1];
  assign popcount33_6wfk_core_149 = input_a[18] ^ input_a[6];
  assign popcount33_6wfk_core_150 = input_a[2] | input_a[28];
  assign popcount33_6wfk_core_151 = input_a[24] | input_a[15];
  assign popcount33_6wfk_core_152 = ~(input_a[15] ^ input_a[9]);
  assign popcount33_6wfk_core_153 = ~input_a[1];
  assign popcount33_6wfk_core_155 = ~(input_a[30] ^ input_a[14]);
  assign popcount33_6wfk_core_156 = ~(input_a[30] | input_a[17]);
  assign popcount33_6wfk_core_159 = input_a[4] & input_a[6];
  assign popcount33_6wfk_core_160_not = ~input_a[29];
  assign popcount33_6wfk_core_161 = ~(input_a[21] & input_a[15]);
  assign popcount33_6wfk_core_162 = ~(input_a[2] | input_a[15]);
  assign popcount33_6wfk_core_163 = ~(input_a[16] & input_a[25]);
  assign popcount33_6wfk_core_165 = input_a[21] & input_a[31];
  assign popcount33_6wfk_core_167 = input_a[27] ^ input_a[2];
  assign popcount33_6wfk_core_168 = input_a[22] | input_a[16];
  assign popcount33_6wfk_core_169 = ~input_a[23];
  assign popcount33_6wfk_core_170 = ~(input_a[22] ^ input_a[15]);
  assign popcount33_6wfk_core_173 = ~(input_a[16] & input_a[5]);
  assign popcount33_6wfk_core_177 = input_a[21] ^ input_a[28];
  assign popcount33_6wfk_core_181 = ~(input_a[28] | input_a[22]);
  assign popcount33_6wfk_core_183 = input_a[13] & input_a[26];
  assign popcount33_6wfk_core_185 = input_a[15] & input_a[26];
  assign popcount33_6wfk_core_186 = input_a[17] | input_a[7];
  assign popcount33_6wfk_core_187 = input_a[8] & input_a[20];
  assign popcount33_6wfk_core_189 = input_a[10] ^ input_a[12];
  assign popcount33_6wfk_core_190 = input_a[6] & input_a[22];
  assign popcount33_6wfk_core_191 = input_a[24] | input_a[4];
  assign popcount33_6wfk_core_192 = input_a[32] ^ input_a[26];
  assign popcount33_6wfk_core_194 = input_a[3] & input_a[3];
  assign popcount33_6wfk_core_195 = ~(input_a[22] | input_a[13]);
  assign popcount33_6wfk_core_196_not = ~input_a[18];
  assign popcount33_6wfk_core_197 = ~(input_a[20] & input_a[25]);
  assign popcount33_6wfk_core_198 = ~(input_a[21] & input_a[19]);
  assign popcount33_6wfk_core_199 = input_a[22] | input_a[29];
  assign popcount33_6wfk_core_200 = input_a[22] ^ input_a[23];
  assign popcount33_6wfk_core_201 = ~(input_a[20] | input_a[5]);
  assign popcount33_6wfk_core_202 = input_a[20] & input_a[18];
  assign popcount33_6wfk_core_205 = ~(input_a[10] | input_a[13]);
  assign popcount33_6wfk_core_206 = ~input_a[29];
  assign popcount33_6wfk_core_207 = input_a[16] ^ input_a[31];
  assign popcount33_6wfk_core_208 = input_a[7] & input_a[0];
  assign popcount33_6wfk_core_209 = input_a[9] ^ input_a[4];
  assign popcount33_6wfk_core_211 = input_a[29] & input_a[32];
  assign popcount33_6wfk_core_212 = ~(input_a[18] | input_a[27]);
  assign popcount33_6wfk_core_216 = input_a[30] ^ input_a[14];
  assign popcount33_6wfk_core_217 = input_a[5] & input_a[17];
  assign popcount33_6wfk_core_218 = input_a[29] | input_a[16];
  assign popcount33_6wfk_core_220 = input_a[0] | input_a[15];
  assign popcount33_6wfk_core_224 = ~(input_a[4] | input_a[12]);
  assign popcount33_6wfk_core_225 = input_a[3] & input_a[30];
  assign popcount33_6wfk_core_226 = ~(input_a[23] & input_a[30]);
  assign popcount33_6wfk_core_227 = input_a[24] ^ input_a[10];
  assign popcount33_6wfk_core_228 = ~(input_a[22] | input_a[14]);
  assign popcount33_6wfk_core_233 = ~(input_a[27] | input_a[25]);
  assign popcount33_6wfk_core_235 = ~(input_a[15] & input_a[22]);

  assign popcount33_6wfk_out[0] = input_a[10];
  assign popcount33_6wfk_out[1] = input_a[18];
  assign popcount33_6wfk_out[2] = 1'b1;
  assign popcount33_6wfk_out[3] = 1'b0;
  assign popcount33_6wfk_out[4] = 1'b1;
  assign popcount33_6wfk_out[5] = 1'b0;
endmodule