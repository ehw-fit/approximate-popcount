// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.99895
// WCE=20.0
// EP=0.842421%
// Printed PDK parameters:
//  Area=78870008.0
//  Delay=79433984.0
//  Power=3569100.0

module popcount40_xehm(input [39:0] input_a, output [5:0] popcount40_xehm_out);
  wire popcount40_xehm_core_042;
  wire popcount40_xehm_core_043;
  wire popcount40_xehm_core_044;
  wire popcount40_xehm_core_045;
  wire popcount40_xehm_core_046;
  wire popcount40_xehm_core_051;
  wire popcount40_xehm_core_052;
  wire popcount40_xehm_core_053;
  wire popcount40_xehm_core_054;
  wire popcount40_xehm_core_055;
  wire popcount40_xehm_core_056;
  wire popcount40_xehm_core_058;
  wire popcount40_xehm_core_062;
  wire popcount40_xehm_core_064;
  wire popcount40_xehm_core_065;
  wire popcount40_xehm_core_066;
  wire popcount40_xehm_core_067;
  wire popcount40_xehm_core_073;
  wire popcount40_xehm_core_077;
  wire popcount40_xehm_core_081;
  wire popcount40_xehm_core_082;
  wire popcount40_xehm_core_083_not;
  wire popcount40_xehm_core_089;
  wire popcount40_xehm_core_091;
  wire popcount40_xehm_core_093;
  wire popcount40_xehm_core_094;
  wire popcount40_xehm_core_095;
  wire popcount40_xehm_core_096;
  wire popcount40_xehm_core_097;
  wire popcount40_xehm_core_098;
  wire popcount40_xehm_core_099;
  wire popcount40_xehm_core_100;
  wire popcount40_xehm_core_101;
  wire popcount40_xehm_core_102;
  wire popcount40_xehm_core_103;
  wire popcount40_xehm_core_104;
  wire popcount40_xehm_core_105;
  wire popcount40_xehm_core_106;
  wire popcount40_xehm_core_107;
  wire popcount40_xehm_core_108;
  wire popcount40_xehm_core_109;
  wire popcount40_xehm_core_110;
  wire popcount40_xehm_core_111;
  wire popcount40_xehm_core_114;
  wire popcount40_xehm_core_115;
  wire popcount40_xehm_core_118;
  wire popcount40_xehm_core_119;
  wire popcount40_xehm_core_120;
  wire popcount40_xehm_core_121;
  wire popcount40_xehm_core_122;
  wire popcount40_xehm_core_123;
  wire popcount40_xehm_core_124;
  wire popcount40_xehm_core_126;
  wire popcount40_xehm_core_129;
  wire popcount40_xehm_core_130;
  wire popcount40_xehm_core_134;
  wire popcount40_xehm_core_135;
  wire popcount40_xehm_core_136;
  wire popcount40_xehm_core_140;
  wire popcount40_xehm_core_142;
  wire popcount40_xehm_core_143;
  wire popcount40_xehm_core_144;
  wire popcount40_xehm_core_146;
  wire popcount40_xehm_core_147;
  wire popcount40_xehm_core_151;
  wire popcount40_xehm_core_152;
  wire popcount40_xehm_core_153;
  wire popcount40_xehm_core_154;
  wire popcount40_xehm_core_155;
  wire popcount40_xehm_core_156;
  wire popcount40_xehm_core_157;
  wire popcount40_xehm_core_158;
  wire popcount40_xehm_core_159;
  wire popcount40_xehm_core_160;
  wire popcount40_xehm_core_162;
  wire popcount40_xehm_core_165;
  wire popcount40_xehm_core_166;
  wire popcount40_xehm_core_167;
  wire popcount40_xehm_core_169;
  wire popcount40_xehm_core_174;
  wire popcount40_xehm_core_175;
  wire popcount40_xehm_core_176;
  wire popcount40_xehm_core_177;
  wire popcount40_xehm_core_178;
  wire popcount40_xehm_core_179;
  wire popcount40_xehm_core_180;
  wire popcount40_xehm_core_183;
  wire popcount40_xehm_core_184;
  wire popcount40_xehm_core_185;
  wire popcount40_xehm_core_186;
  wire popcount40_xehm_core_187;
  wire popcount40_xehm_core_188;
  wire popcount40_xehm_core_189;
  wire popcount40_xehm_core_192;
  wire popcount40_xehm_core_193;
  wire popcount40_xehm_core_194;
  wire popcount40_xehm_core_195;
  wire popcount40_xehm_core_196;
  wire popcount40_xehm_core_197;
  wire popcount40_xehm_core_199;
  wire popcount40_xehm_core_200;
  wire popcount40_xehm_core_201;
  wire popcount40_xehm_core_202;
  wire popcount40_xehm_core_203;
  wire popcount40_xehm_core_204;
  wire popcount40_xehm_core_205;
  wire popcount40_xehm_core_206;
  wire popcount40_xehm_core_207;
  wire popcount40_xehm_core_208;
  wire popcount40_xehm_core_209;
  wire popcount40_xehm_core_210;
  wire popcount40_xehm_core_211;
  wire popcount40_xehm_core_213;
  wire popcount40_xehm_core_215_not;
  wire popcount40_xehm_core_216;
  wire popcount40_xehm_core_218;
  wire popcount40_xehm_core_219;
  wire popcount40_xehm_core_220;
  wire popcount40_xehm_core_221;
  wire popcount40_xehm_core_222;
  wire popcount40_xehm_core_223;
  wire popcount40_xehm_core_225;
  wire popcount40_xehm_core_226;
  wire popcount40_xehm_core_227;
  wire popcount40_xehm_core_228;
  wire popcount40_xehm_core_229;
  wire popcount40_xehm_core_230;
  wire popcount40_xehm_core_231;
  wire popcount40_xehm_core_233;
  wire popcount40_xehm_core_235;
  wire popcount40_xehm_core_237;
  wire popcount40_xehm_core_240;
  wire popcount40_xehm_core_242;
  wire popcount40_xehm_core_243;
  wire popcount40_xehm_core_244;
  wire popcount40_xehm_core_245;
  wire popcount40_xehm_core_246;
  wire popcount40_xehm_core_247;
  wire popcount40_xehm_core_248;
  wire popcount40_xehm_core_253;
  wire popcount40_xehm_core_254;
  wire popcount40_xehm_core_258;
  wire popcount40_xehm_core_259;
  wire popcount40_xehm_core_260;
  wire popcount40_xehm_core_261;
  wire popcount40_xehm_core_262;
  wire popcount40_xehm_core_268;
  wire popcount40_xehm_core_269;
  wire popcount40_xehm_core_270;
  wire popcount40_xehm_core_271;
  wire popcount40_xehm_core_273;
  wire popcount40_xehm_core_275;
  wire popcount40_xehm_core_276;
  wire popcount40_xehm_core_277;
  wire popcount40_xehm_core_278;
  wire popcount40_xehm_core_279;
  wire popcount40_xehm_core_280;
  wire popcount40_xehm_core_281;
  wire popcount40_xehm_core_282;
  wire popcount40_xehm_core_283;
  wire popcount40_xehm_core_284;
  wire popcount40_xehm_core_286;
  wire popcount40_xehm_core_288;
  wire popcount40_xehm_core_289;
  wire popcount40_xehm_core_294_not;
  wire popcount40_xehm_core_297;
  wire popcount40_xehm_core_298;
  wire popcount40_xehm_core_299;
  wire popcount40_xehm_core_300;
  wire popcount40_xehm_core_301;
  wire popcount40_xehm_core_302;
  wire popcount40_xehm_core_303;
  wire popcount40_xehm_core_304;
  wire popcount40_xehm_core_305;
  wire popcount40_xehm_core_306;
  wire popcount40_xehm_core_307;
  wire popcount40_xehm_core_309;
  wire popcount40_xehm_core_310;
  wire popcount40_xehm_core_311;
  wire popcount40_xehm_core_312;
  wire popcount40_xehm_core_316;

  assign popcount40_xehm_core_042 = input_a[0] ^ input_a[1];
  assign popcount40_xehm_core_043 = input_a[0] & input_a[1];
  assign popcount40_xehm_core_044 = ~(input_a[23] ^ input_a[21]);
  assign popcount40_xehm_core_045 = input_a[18] & input_a[3];
  assign popcount40_xehm_core_046 = input_a[8] | input_a[32];
  assign popcount40_xehm_core_051 = popcount40_xehm_core_042 & input_a[23];
  assign popcount40_xehm_core_052 = popcount40_xehm_core_043 ^ popcount40_xehm_core_045;
  assign popcount40_xehm_core_053 = popcount40_xehm_core_043 & popcount40_xehm_core_045;
  assign popcount40_xehm_core_054 = popcount40_xehm_core_052 ^ popcount40_xehm_core_051;
  assign popcount40_xehm_core_055 = popcount40_xehm_core_052 & popcount40_xehm_core_051;
  assign popcount40_xehm_core_056 = popcount40_xehm_core_053 | popcount40_xehm_core_055;
  assign popcount40_xehm_core_058 = ~(input_a[7] & input_a[5]);
  assign popcount40_xehm_core_062 = input_a[39] | input_a[22];
  assign popcount40_xehm_core_064 = input_a[23] & input_a[22];
  assign popcount40_xehm_core_065 = ~(input_a[5] ^ input_a[35]);
  assign popcount40_xehm_core_066 = ~(input_a[27] & input_a[38]);
  assign popcount40_xehm_core_067 = ~input_a[18];
  assign popcount40_xehm_core_073 = input_a[7] | input_a[24];
  assign popcount40_xehm_core_077 = input_a[37] & input_a[1];
  assign popcount40_xehm_core_081 = input_a[38] & input_a[4];
  assign popcount40_xehm_core_082 = ~(input_a[11] & input_a[14]);
  assign popcount40_xehm_core_083_not = ~popcount40_xehm_core_056;
  assign popcount40_xehm_core_089 = input_a[22] ^ input_a[24];
  assign popcount40_xehm_core_091 = input_a[13] & input_a[11];
  assign popcount40_xehm_core_093 = input_a[10] ^ input_a[11];
  assign popcount40_xehm_core_094 = input_a[10] & input_a[11];
  assign popcount40_xehm_core_095 = input_a[13] ^ input_a[14];
  assign popcount40_xehm_core_096 = input_a[13] & input_a[14];
  assign popcount40_xehm_core_097 = ~(input_a[12] & popcount40_xehm_core_095);
  assign popcount40_xehm_core_098 = input_a[12] & popcount40_xehm_core_095;
  assign popcount40_xehm_core_099 = popcount40_xehm_core_096 ^ popcount40_xehm_core_098;
  assign popcount40_xehm_core_100 = popcount40_xehm_core_096 & input_a[20];
  assign popcount40_xehm_core_101 = ~(input_a[37] & input_a[29]);
  assign popcount40_xehm_core_102 = popcount40_xehm_core_093 & popcount40_xehm_core_097;
  assign popcount40_xehm_core_103 = popcount40_xehm_core_094 ^ popcount40_xehm_core_099;
  assign popcount40_xehm_core_104 = popcount40_xehm_core_094 & popcount40_xehm_core_099;
  assign popcount40_xehm_core_105 = popcount40_xehm_core_103 ^ popcount40_xehm_core_102;
  assign popcount40_xehm_core_106 = popcount40_xehm_core_103 & popcount40_xehm_core_102;
  assign popcount40_xehm_core_107 = popcount40_xehm_core_104 | popcount40_xehm_core_106;
  assign popcount40_xehm_core_108 = popcount40_xehm_core_100 | popcount40_xehm_core_107;
  assign popcount40_xehm_core_109 = input_a[39] & input_a[12];
  assign popcount40_xehm_core_110 = input_a[15] ^ input_a[16];
  assign popcount40_xehm_core_111 = input_a[15] & input_a[16];
  assign popcount40_xehm_core_114 = ~(input_a[17] & input_a[22]);
  assign popcount40_xehm_core_115 = input_a[17] & input_a[22];
  assign popcount40_xehm_core_118 = ~(input_a[9] & input_a[31]);
  assign popcount40_xehm_core_119 = popcount40_xehm_core_110 & popcount40_xehm_core_114;
  assign popcount40_xehm_core_120 = popcount40_xehm_core_111 ^ popcount40_xehm_core_115;
  assign popcount40_xehm_core_121 = popcount40_xehm_core_111 & popcount40_xehm_core_115;
  assign popcount40_xehm_core_122 = popcount40_xehm_core_120 ^ popcount40_xehm_core_119;
  assign popcount40_xehm_core_123 = popcount40_xehm_core_120 & popcount40_xehm_core_119;
  assign popcount40_xehm_core_124 = popcount40_xehm_core_121 | popcount40_xehm_core_123;
  assign popcount40_xehm_core_126 = input_a[38] | input_a[21];
  assign popcount40_xehm_core_129 = popcount40_xehm_core_105 ^ popcount40_xehm_core_122;
  assign popcount40_xehm_core_130 = popcount40_xehm_core_105 & popcount40_xehm_core_122;
  assign popcount40_xehm_core_134 = popcount40_xehm_core_108 ^ popcount40_xehm_core_124;
  assign popcount40_xehm_core_135 = popcount40_xehm_core_108 & popcount40_xehm_core_124;
  assign popcount40_xehm_core_136 = popcount40_xehm_core_134 | popcount40_xehm_core_130;
  assign popcount40_xehm_core_140 = input_a[11] & input_a[7];
  assign popcount40_xehm_core_142 = input_a[4] & input_a[25];
  assign popcount40_xehm_core_143 = ~input_a[38];
  assign popcount40_xehm_core_144 = input_a[20] | input_a[29];
  assign popcount40_xehm_core_146 = input_a[32] ^ input_a[11];
  assign popcount40_xehm_core_147 = popcount40_xehm_core_054 & popcount40_xehm_core_129;
  assign popcount40_xehm_core_151 = popcount40_xehm_core_083_not ^ popcount40_xehm_core_136;
  assign popcount40_xehm_core_152 = popcount40_xehm_core_083_not & popcount40_xehm_core_136;
  assign popcount40_xehm_core_153 = popcount40_xehm_core_151 ^ popcount40_xehm_core_147;
  assign popcount40_xehm_core_154 = popcount40_xehm_core_151 & popcount40_xehm_core_147;
  assign popcount40_xehm_core_155 = popcount40_xehm_core_152 | popcount40_xehm_core_154;
  assign popcount40_xehm_core_156 = popcount40_xehm_core_056 | popcount40_xehm_core_135;
  assign popcount40_xehm_core_157 = input_a[22] & popcount40_xehm_core_135;
  assign popcount40_xehm_core_158 = popcount40_xehm_core_156 ^ popcount40_xehm_core_155;
  assign popcount40_xehm_core_159 = ~(popcount40_xehm_core_156 | popcount40_xehm_core_155);
  assign popcount40_xehm_core_160 = popcount40_xehm_core_157 & popcount40_xehm_core_159;
  assign popcount40_xehm_core_162 = ~input_a[24];
  assign popcount40_xehm_core_165 = ~(input_a[6] | input_a[0]);
  assign popcount40_xehm_core_166 = input_a[10] ^ input_a[32];
  assign popcount40_xehm_core_167 = input_a[20] & input_a[21];
  assign popcount40_xehm_core_169 = input_a[8] & input_a[24];
  assign popcount40_xehm_core_174 = ~(input_a[8] & input_a[24]);
  assign popcount40_xehm_core_175 = input_a[38] & input_a[24];
  assign popcount40_xehm_core_176 = popcount40_xehm_core_167 ^ popcount40_xehm_core_169;
  assign popcount40_xehm_core_177 = popcount40_xehm_core_167 & popcount40_xehm_core_169;
  assign popcount40_xehm_core_178 = popcount40_xehm_core_176 ^ popcount40_xehm_core_175;
  assign popcount40_xehm_core_179 = popcount40_xehm_core_176 & popcount40_xehm_core_175;
  assign popcount40_xehm_core_180 = popcount40_xehm_core_177 | popcount40_xehm_core_179;
  assign popcount40_xehm_core_183 = input_a[25] ^ input_a[26];
  assign popcount40_xehm_core_184 = input_a[25] & input_a[26];
  assign popcount40_xehm_core_185 = input_a[28] ^ input_a[29];
  assign popcount40_xehm_core_186 = input_a[28] & input_a[29];
  assign popcount40_xehm_core_187 = input_a[27] ^ popcount40_xehm_core_185;
  assign popcount40_xehm_core_188 = input_a[27] & popcount40_xehm_core_185;
  assign popcount40_xehm_core_189 = popcount40_xehm_core_186 | popcount40_xehm_core_188;
  assign popcount40_xehm_core_192 = popcount40_xehm_core_183 & popcount40_xehm_core_187;
  assign popcount40_xehm_core_193 = popcount40_xehm_core_184 ^ popcount40_xehm_core_189;
  assign popcount40_xehm_core_194 = popcount40_xehm_core_184 & popcount40_xehm_core_189;
  assign popcount40_xehm_core_195 = popcount40_xehm_core_193 ^ popcount40_xehm_core_192;
  assign popcount40_xehm_core_196 = popcount40_xehm_core_193 & popcount40_xehm_core_192;
  assign popcount40_xehm_core_197 = popcount40_xehm_core_194 | popcount40_xehm_core_196;
  assign popcount40_xehm_core_199 = ~(input_a[22] | input_a[11]);
  assign popcount40_xehm_core_200 = ~(input_a[20] ^ input_a[31]);
  assign popcount40_xehm_core_201 = popcount40_xehm_core_174 & input_a[8];
  assign popcount40_xehm_core_202 = popcount40_xehm_core_178 ^ popcount40_xehm_core_195;
  assign popcount40_xehm_core_203 = popcount40_xehm_core_178 & popcount40_xehm_core_195;
  assign popcount40_xehm_core_204 = popcount40_xehm_core_202 ^ popcount40_xehm_core_201;
  assign popcount40_xehm_core_205 = popcount40_xehm_core_202 & popcount40_xehm_core_201;
  assign popcount40_xehm_core_206 = popcount40_xehm_core_203 | popcount40_xehm_core_205;
  assign popcount40_xehm_core_207 = popcount40_xehm_core_180 ^ popcount40_xehm_core_197;
  assign popcount40_xehm_core_208 = popcount40_xehm_core_180 & popcount40_xehm_core_197;
  assign popcount40_xehm_core_209 = popcount40_xehm_core_207 ^ popcount40_xehm_core_206;
  assign popcount40_xehm_core_210 = popcount40_xehm_core_207 & popcount40_xehm_core_206;
  assign popcount40_xehm_core_211 = popcount40_xehm_core_208 | popcount40_xehm_core_210;
  assign popcount40_xehm_core_213 = input_a[9] ^ input_a[12];
  assign popcount40_xehm_core_215_not = ~input_a[13];
  assign popcount40_xehm_core_216 = ~(input_a[32] & input_a[0]);
  assign popcount40_xehm_core_218 = input_a[30] & input_a[6];
  assign popcount40_xehm_core_219 = input_a[33] ^ input_a[34];
  assign popcount40_xehm_core_220 = input_a[33] & input_a[34];
  assign popcount40_xehm_core_221 = input_a[32] ^ popcount40_xehm_core_219;
  assign popcount40_xehm_core_222 = input_a[32] & popcount40_xehm_core_219;
  assign popcount40_xehm_core_223 = popcount40_xehm_core_220 | popcount40_xehm_core_222;
  assign popcount40_xehm_core_225 = ~(input_a[36] ^ input_a[0]);
  assign popcount40_xehm_core_226 = input_a[36] & popcount40_xehm_core_221;
  assign popcount40_xehm_core_227 = popcount40_xehm_core_218 ^ popcount40_xehm_core_223;
  assign popcount40_xehm_core_228 = popcount40_xehm_core_218 & popcount40_xehm_core_223;
  assign popcount40_xehm_core_229 = popcount40_xehm_core_227 ^ popcount40_xehm_core_226;
  assign popcount40_xehm_core_230 = popcount40_xehm_core_227 & popcount40_xehm_core_226;
  assign popcount40_xehm_core_231 = popcount40_xehm_core_228 | popcount40_xehm_core_230;
  assign popcount40_xehm_core_233 = ~(input_a[38] & input_a[7]);
  assign popcount40_xehm_core_235 = input_a[35] & input_a[27];
  assign popcount40_xehm_core_237 = input_a[2] & input_a[2];
  assign popcount40_xehm_core_240 = popcount40_xehm_core_237 | input_a[4];
  assign popcount40_xehm_core_242 = ~input_a[35];
  assign popcount40_xehm_core_243 = input_a[7] & input_a[9];
  assign popcount40_xehm_core_244 = popcount40_xehm_core_235 ^ popcount40_xehm_core_240;
  assign popcount40_xehm_core_245 = popcount40_xehm_core_235 & popcount40_xehm_core_240;
  assign popcount40_xehm_core_246 = popcount40_xehm_core_244 ^ popcount40_xehm_core_243;
  assign popcount40_xehm_core_247 = popcount40_xehm_core_244 & popcount40_xehm_core_243;
  assign popcount40_xehm_core_248 = popcount40_xehm_core_245 | popcount40_xehm_core_247;
  assign popcount40_xehm_core_253 = popcount40_xehm_core_229 ^ popcount40_xehm_core_246;
  assign popcount40_xehm_core_254 = popcount40_xehm_core_229 & popcount40_xehm_core_246;
  assign popcount40_xehm_core_258 = popcount40_xehm_core_231 ^ popcount40_xehm_core_248;
  assign popcount40_xehm_core_259 = popcount40_xehm_core_231 & popcount40_xehm_core_248;
  assign popcount40_xehm_core_260 = popcount40_xehm_core_258 ^ popcount40_xehm_core_254;
  assign popcount40_xehm_core_261 = popcount40_xehm_core_258 & popcount40_xehm_core_254;
  assign popcount40_xehm_core_262 = popcount40_xehm_core_259 | popcount40_xehm_core_261;
  assign popcount40_xehm_core_268 = input_a[34] | input_a[5];
  assign popcount40_xehm_core_269 = ~(popcount40_xehm_core_200 ^ input_a[24]);
  assign popcount40_xehm_core_270 = popcount40_xehm_core_204 ^ popcount40_xehm_core_253;
  assign popcount40_xehm_core_271 = popcount40_xehm_core_204 & popcount40_xehm_core_253;
  assign popcount40_xehm_core_273 = input_a[17] ^ input_a[12];
  assign popcount40_xehm_core_275 = popcount40_xehm_core_209 ^ popcount40_xehm_core_260;
  assign popcount40_xehm_core_276 = popcount40_xehm_core_209 & popcount40_xehm_core_260;
  assign popcount40_xehm_core_277 = popcount40_xehm_core_275 ^ popcount40_xehm_core_271;
  assign popcount40_xehm_core_278 = popcount40_xehm_core_275 & popcount40_xehm_core_271;
  assign popcount40_xehm_core_279 = popcount40_xehm_core_276 | popcount40_xehm_core_278;
  assign popcount40_xehm_core_280 = popcount40_xehm_core_211 | popcount40_xehm_core_262;
  assign popcount40_xehm_core_281 = popcount40_xehm_core_211 & popcount40_xehm_core_262;
  assign popcount40_xehm_core_282 = popcount40_xehm_core_280 ^ popcount40_xehm_core_279;
  assign popcount40_xehm_core_283 = popcount40_xehm_core_280 & popcount40_xehm_core_279;
  assign popcount40_xehm_core_284 = popcount40_xehm_core_281 | popcount40_xehm_core_283;
  assign popcount40_xehm_core_286 = ~(input_a[36] & input_a[37]);
  assign popcount40_xehm_core_288 = input_a[2] ^ input_a[21];
  assign popcount40_xehm_core_289 = ~(input_a[9] & input_a[18]);
  assign popcount40_xehm_core_294_not = ~popcount40_xehm_core_270;
  assign popcount40_xehm_core_297 = popcount40_xehm_core_153 ^ popcount40_xehm_core_277;
  assign popcount40_xehm_core_298 = popcount40_xehm_core_153 & popcount40_xehm_core_277;
  assign popcount40_xehm_core_299 = popcount40_xehm_core_297 ^ popcount40_xehm_core_270;
  assign popcount40_xehm_core_300 = popcount40_xehm_core_297 & popcount40_xehm_core_270;
  assign popcount40_xehm_core_301 = popcount40_xehm_core_298 | popcount40_xehm_core_300;
  assign popcount40_xehm_core_302 = popcount40_xehm_core_158 ^ popcount40_xehm_core_282;
  assign popcount40_xehm_core_303 = popcount40_xehm_core_158 & popcount40_xehm_core_282;
  assign popcount40_xehm_core_304 = popcount40_xehm_core_302 ^ popcount40_xehm_core_301;
  assign popcount40_xehm_core_305 = popcount40_xehm_core_302 & popcount40_xehm_core_301;
  assign popcount40_xehm_core_306 = popcount40_xehm_core_303 | popcount40_xehm_core_305;
  assign popcount40_xehm_core_307 = popcount40_xehm_core_160 | popcount40_xehm_core_284;
  assign popcount40_xehm_core_309 = popcount40_xehm_core_307 | popcount40_xehm_core_306;
  assign popcount40_xehm_core_310 = ~(input_a[37] & input_a[29]);
  assign popcount40_xehm_core_311 = input_a[21] | input_a[0];
  assign popcount40_xehm_core_312 = input_a[4] ^ input_a[2];
  assign popcount40_xehm_core_316 = ~(input_a[8] | input_a[6]);

  assign popcount40_xehm_out[0] = 1'b1;
  assign popcount40_xehm_out[1] = popcount40_xehm_core_294_not;
  assign popcount40_xehm_out[2] = popcount40_xehm_core_299;
  assign popcount40_xehm_out[3] = popcount40_xehm_core_304;
  assign popcount40_xehm_out[4] = popcount40_xehm_core_309;
  assign popcount40_xehm_out[5] = 1'b0;
endmodule