// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.47543
// WCE=14.0
// EP=0.875326%
// Printed PDK parameters:
//  Area=7417840.0
//  Delay=15507594.0
//  Power=357240.0

module popcount28_e9p1(input [27:0] input_a, output [4:0] popcount28_e9p1_out);
  wire popcount28_e9p1_core_030;
  wire popcount28_e9p1_core_032;
  wire popcount28_e9p1_core_034;
  wire popcount28_e9p1_core_035_not;
  wire popcount28_e9p1_core_036;
  wire popcount28_e9p1_core_038;
  wire popcount28_e9p1_core_039;
  wire popcount28_e9p1_core_040;
  wire popcount28_e9p1_core_041;
  wire popcount28_e9p1_core_042;
  wire popcount28_e9p1_core_043;
  wire popcount28_e9p1_core_044;
  wire popcount28_e9p1_core_046;
  wire popcount28_e9p1_core_047;
  wire popcount28_e9p1_core_048;
  wire popcount28_e9p1_core_049;
  wire popcount28_e9p1_core_050;
  wire popcount28_e9p1_core_051;
  wire popcount28_e9p1_core_054;
  wire popcount28_e9p1_core_055;
  wire popcount28_e9p1_core_056;
  wire popcount28_e9p1_core_058;
  wire popcount28_e9p1_core_065;
  wire popcount28_e9p1_core_069;
  wire popcount28_e9p1_core_070;
  wire popcount28_e9p1_core_071;
  wire popcount28_e9p1_core_072;
  wire popcount28_e9p1_core_073;
  wire popcount28_e9p1_core_074;
  wire popcount28_e9p1_core_075;
  wire popcount28_e9p1_core_076;
  wire popcount28_e9p1_core_077;
  wire popcount28_e9p1_core_078;
  wire popcount28_e9p1_core_079;
  wire popcount28_e9p1_core_080_not;
  wire popcount28_e9p1_core_081_not;
  wire popcount28_e9p1_core_082;
  wire popcount28_e9p1_core_087;
  wire popcount28_e9p1_core_089;
  wire popcount28_e9p1_core_090;
  wire popcount28_e9p1_core_091;
  wire popcount28_e9p1_core_094;
  wire popcount28_e9p1_core_095;
  wire popcount28_e9p1_core_097;
  wire popcount28_e9p1_core_098;
  wire popcount28_e9p1_core_101;
  wire popcount28_e9p1_core_102;
  wire popcount28_e9p1_core_104;
  wire popcount28_e9p1_core_106;
  wire popcount28_e9p1_core_107;
  wire popcount28_e9p1_core_108;
  wire popcount28_e9p1_core_109;
  wire popcount28_e9p1_core_111;
  wire popcount28_e9p1_core_113;
  wire popcount28_e9p1_core_114;
  wire popcount28_e9p1_core_115;
  wire popcount28_e9p1_core_116;
  wire popcount28_e9p1_core_119;
  wire popcount28_e9p1_core_120;
  wire popcount28_e9p1_core_122;
  wire popcount28_e9p1_core_124;
  wire popcount28_e9p1_core_125;
  wire popcount28_e9p1_core_126;
  wire popcount28_e9p1_core_127;
  wire popcount28_e9p1_core_130;
  wire popcount28_e9p1_core_133;
  wire popcount28_e9p1_core_135;
  wire popcount28_e9p1_core_136;
  wire popcount28_e9p1_core_137;
  wire popcount28_e9p1_core_138;
  wire popcount28_e9p1_core_139;
  wire popcount28_e9p1_core_140;
  wire popcount28_e9p1_core_142;
  wire popcount28_e9p1_core_146;
  wire popcount28_e9p1_core_149;
  wire popcount28_e9p1_core_150;
  wire popcount28_e9p1_core_151;
  wire popcount28_e9p1_core_152;
  wire popcount28_e9p1_core_153;
  wire popcount28_e9p1_core_154;
  wire popcount28_e9p1_core_156;
  wire popcount28_e9p1_core_157_not;
  wire popcount28_e9p1_core_162_not;
  wire popcount28_e9p1_core_163;
  wire popcount28_e9p1_core_164;
  wire popcount28_e9p1_core_169;
  wire popcount28_e9p1_core_170;
  wire popcount28_e9p1_core_171;
  wire popcount28_e9p1_core_173;
  wire popcount28_e9p1_core_178;
  wire popcount28_e9p1_core_179;
  wire popcount28_e9p1_core_183;
  wire popcount28_e9p1_core_184;
  wire popcount28_e9p1_core_186;
  wire popcount28_e9p1_core_187;
  wire popcount28_e9p1_core_188;
  wire popcount28_e9p1_core_189;
  wire popcount28_e9p1_core_190;
  wire popcount28_e9p1_core_192;
  wire popcount28_e9p1_core_193;
  wire popcount28_e9p1_core_194;
  wire popcount28_e9p1_core_195;
  wire popcount28_e9p1_core_196;
  wire popcount28_e9p1_core_198;
  wire popcount28_e9p1_core_201;

  assign popcount28_e9p1_core_030 = input_a[21] & input_a[12];
  assign popcount28_e9p1_core_032 = ~(input_a[1] ^ input_a[10]);
  assign popcount28_e9p1_core_034 = input_a[7] & input_a[5];
  assign popcount28_e9p1_core_035_not = ~input_a[21];
  assign popcount28_e9p1_core_036 = input_a[3] | input_a[21];
  assign popcount28_e9p1_core_038 = ~(input_a[18] & input_a[20]);
  assign popcount28_e9p1_core_039 = ~(input_a[23] | input_a[6]);
  assign popcount28_e9p1_core_040 = ~(input_a[4] & input_a[15]);
  assign popcount28_e9p1_core_041 = input_a[17] & input_a[4];
  assign popcount28_e9p1_core_042 = ~(input_a[12] | input_a[18]);
  assign popcount28_e9p1_core_043 = input_a[25] ^ input_a[15];
  assign popcount28_e9p1_core_044 = input_a[26] ^ input_a[11];
  assign popcount28_e9p1_core_046 = input_a[23] | input_a[21];
  assign popcount28_e9p1_core_047 = ~(input_a[14] ^ input_a[4]);
  assign popcount28_e9p1_core_048 = input_a[22] & input_a[13];
  assign popcount28_e9p1_core_049 = ~(input_a[8] & input_a[10]);
  assign popcount28_e9p1_core_050 = input_a[1] | input_a[17];
  assign popcount28_e9p1_core_051 = ~(input_a[16] | input_a[22]);
  assign popcount28_e9p1_core_054 = input_a[26] | popcount28_e9p1_core_046;
  assign popcount28_e9p1_core_055 = input_a[3] ^ input_a[2];
  assign popcount28_e9p1_core_056 = popcount28_e9p1_core_054 | input_a[17];
  assign popcount28_e9p1_core_058 = ~(input_a[2] & input_a[16]);
  assign popcount28_e9p1_core_065 = input_a[15] & input_a[19];
  assign popcount28_e9p1_core_069 = ~(input_a[2] ^ input_a[6]);
  assign popcount28_e9p1_core_070 = ~input_a[8];
  assign popcount28_e9p1_core_071 = ~(input_a[2] ^ input_a[0]);
  assign popcount28_e9p1_core_072 = ~(input_a[4] ^ input_a[0]);
  assign popcount28_e9p1_core_073 = ~input_a[3];
  assign popcount28_e9p1_core_074 = ~input_a[0];
  assign popcount28_e9p1_core_075 = ~(input_a[27] & input_a[2]);
  assign popcount28_e9p1_core_076 = ~(input_a[13] ^ input_a[15]);
  assign popcount28_e9p1_core_077 = ~input_a[22];
  assign popcount28_e9p1_core_078 = input_a[11] & input_a[3];
  assign popcount28_e9p1_core_079 = ~(input_a[26] | input_a[20]);
  assign popcount28_e9p1_core_080_not = ~input_a[13];
  assign popcount28_e9p1_core_081_not = ~input_a[2];
  assign popcount28_e9p1_core_082 = input_a[17] & input_a[19];
  assign popcount28_e9p1_core_087 = ~(input_a[21] | input_a[6]);
  assign popcount28_e9p1_core_089 = ~(input_a[27] & input_a[7]);
  assign popcount28_e9p1_core_090 = input_a[7] & input_a[23];
  assign popcount28_e9p1_core_091 = input_a[9] ^ input_a[11];
  assign popcount28_e9p1_core_094 = input_a[3] | input_a[7];
  assign popcount28_e9p1_core_095 = ~popcount28_e9p1_core_056;
  assign popcount28_e9p1_core_097 = popcount28_e9p1_core_095 ^ input_a[24];
  assign popcount28_e9p1_core_098 = ~(input_a[26] ^ input_a[7]);
  assign popcount28_e9p1_core_101 = input_a[20] ^ input_a[25];
  assign popcount28_e9p1_core_102 = input_a[24] | popcount28_e9p1_core_056;
  assign popcount28_e9p1_core_104 = ~(input_a[25] & input_a[19]);
  assign popcount28_e9p1_core_106 = ~(input_a[7] ^ input_a[3]);
  assign popcount28_e9p1_core_107 = input_a[11] ^ input_a[24];
  assign popcount28_e9p1_core_108 = ~(input_a[17] | input_a[12]);
  assign popcount28_e9p1_core_109 = ~input_a[25];
  assign popcount28_e9p1_core_111 = input_a[27] ^ input_a[5];
  assign popcount28_e9p1_core_113 = ~(input_a[10] ^ input_a[20]);
  assign popcount28_e9p1_core_114 = input_a[8] & input_a[11];
  assign popcount28_e9p1_core_115 = ~input_a[8];
  assign popcount28_e9p1_core_116 = input_a[20] & input_a[12];
  assign popcount28_e9p1_core_119 = ~(input_a[14] ^ input_a[14]);
  assign popcount28_e9p1_core_120 = popcount28_e9p1_core_114 & popcount28_e9p1_core_116;
  assign popcount28_e9p1_core_122 = ~(input_a[2] & input_a[9]);
  assign popcount28_e9p1_core_124 = ~input_a[14];
  assign popcount28_e9p1_core_125 = ~input_a[18];
  assign popcount28_e9p1_core_126 = ~(input_a[23] | input_a[4]);
  assign popcount28_e9p1_core_127 = ~(input_a[13] | input_a[0]);
  assign popcount28_e9p1_core_130 = ~(input_a[9] & input_a[0]);
  assign popcount28_e9p1_core_133 = input_a[10] ^ input_a[2];
  assign popcount28_e9p1_core_135 = input_a[2] & input_a[14];
  assign popcount28_e9p1_core_136 = input_a[24] ^ input_a[18];
  assign popcount28_e9p1_core_137 = input_a[6] & input_a[15];
  assign popcount28_e9p1_core_138 = ~input_a[17];
  assign popcount28_e9p1_core_139 = popcount28_e9p1_core_135 & popcount28_e9p1_core_137;
  assign popcount28_e9p1_core_140 = input_a[11] | input_a[27];
  assign popcount28_e9p1_core_142 = ~(input_a[1] | input_a[2]);
  assign popcount28_e9p1_core_146 = ~(input_a[3] ^ input_a[22]);
  assign popcount28_e9p1_core_149 = ~(input_a[15] | input_a[23]);
  assign popcount28_e9p1_core_150 = ~input_a[26];
  assign popcount28_e9p1_core_151 = ~(input_a[17] ^ input_a[3]);
  assign popcount28_e9p1_core_152 = ~(input_a[15] & input_a[11]);
  assign popcount28_e9p1_core_153 = ~(input_a[1] | input_a[12]);
  assign popcount28_e9p1_core_154 = ~(input_a[1] ^ input_a[0]);
  assign popcount28_e9p1_core_156 = input_a[18] ^ input_a[24];
  assign popcount28_e9p1_core_157_not = ~input_a[12];
  assign popcount28_e9p1_core_162_not = ~input_a[20];
  assign popcount28_e9p1_core_163 = ~(input_a[7] ^ input_a[22]);
  assign popcount28_e9p1_core_164 = ~(input_a[20] & input_a[17]);
  assign popcount28_e9p1_core_169 = ~(input_a[3] | input_a[9]);
  assign popcount28_e9p1_core_170 = popcount28_e9p1_core_120 ^ popcount28_e9p1_core_139;
  assign popcount28_e9p1_core_171 = popcount28_e9p1_core_120 & popcount28_e9p1_core_139;
  assign popcount28_e9p1_core_173 = ~(input_a[25] ^ input_a[1]);
  assign popcount28_e9p1_core_178 = input_a[20] & input_a[21];
  assign popcount28_e9p1_core_179 = ~input_a[21];
  assign popcount28_e9p1_core_183 = ~input_a[7];
  assign popcount28_e9p1_core_184 = ~(input_a[10] ^ input_a[15]);
  assign popcount28_e9p1_core_186 = input_a[0] ^ input_a[11];
  assign popcount28_e9p1_core_187 = ~(input_a[2] ^ input_a[5]);
  assign popcount28_e9p1_core_188 = popcount28_e9p1_core_097 & popcount28_e9p1_core_170;
  assign popcount28_e9p1_core_189 = input_a[9] ^ input_a[15];
  assign popcount28_e9p1_core_190 = input_a[15] | input_a[13];
  assign popcount28_e9p1_core_192 = popcount28_e9p1_core_102 ^ popcount28_e9p1_core_171;
  assign popcount28_e9p1_core_193 = popcount28_e9p1_core_102 & popcount28_e9p1_core_171;
  assign popcount28_e9p1_core_194 = popcount28_e9p1_core_192 ^ popcount28_e9p1_core_188;
  assign popcount28_e9p1_core_195 = input_a[24] & popcount28_e9p1_core_188;
  assign popcount28_e9p1_core_196 = popcount28_e9p1_core_193 | popcount28_e9p1_core_195;
  assign popcount28_e9p1_core_198 = input_a[12] & input_a[19];
  assign popcount28_e9p1_core_201 = ~(input_a[18] | input_a[26]);

  assign popcount28_e9p1_out[0] = input_a[0];
  assign popcount28_e9p1_out[1] = popcount28_e9p1_core_095;
  assign popcount28_e9p1_out[2] = 1'b1;
  assign popcount28_e9p1_out[3] = popcount28_e9p1_core_194;
  assign popcount28_e9p1_out[4] = popcount28_e9p1_core_196;
endmodule