// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.24722
// WCE=14.0
// EP=0.861624%
// Printed PDK parameters:
//  Area=476280.0
//  Delay=2551099.0
//  Power=3460.8

module popcount27_6onj(input [26:0] input_a, output [4:0] popcount27_6onj_out);
  wire popcount27_6onj_core_029;
  wire popcount27_6onj_core_030;
  wire popcount27_6onj_core_031;
  wire popcount27_6onj_core_033;
  wire popcount27_6onj_core_036;
  wire popcount27_6onj_core_037;
  wire popcount27_6onj_core_038;
  wire popcount27_6onj_core_039;
  wire popcount27_6onj_core_041;
  wire popcount27_6onj_core_042;
  wire popcount27_6onj_core_045;
  wire popcount27_6onj_core_046_not;
  wire popcount27_6onj_core_048;
  wire popcount27_6onj_core_050;
  wire popcount27_6onj_core_052;
  wire popcount27_6onj_core_053;
  wire popcount27_6onj_core_054;
  wire popcount27_6onj_core_055;
  wire popcount27_6onj_core_057;
  wire popcount27_6onj_core_058;
  wire popcount27_6onj_core_060;
  wire popcount27_6onj_core_061;
  wire popcount27_6onj_core_064;
  wire popcount27_6onj_core_065;
  wire popcount27_6onj_core_066;
  wire popcount27_6onj_core_067;
  wire popcount27_6onj_core_069;
  wire popcount27_6onj_core_070;
  wire popcount27_6onj_core_071;
  wire popcount27_6onj_core_072_not;
  wire popcount27_6onj_core_073;
  wire popcount27_6onj_core_074;
  wire popcount27_6onj_core_075;
  wire popcount27_6onj_core_076;
  wire popcount27_6onj_core_077;
  wire popcount27_6onj_core_078;
  wire popcount27_6onj_core_079;
  wire popcount27_6onj_core_082;
  wire popcount27_6onj_core_083_not;
  wire popcount27_6onj_core_084;
  wire popcount27_6onj_core_087;
  wire popcount27_6onj_core_089;
  wire popcount27_6onj_core_090;
  wire popcount27_6onj_core_091;
  wire popcount27_6onj_core_092;
  wire popcount27_6onj_core_093;
  wire popcount27_6onj_core_094;
  wire popcount27_6onj_core_095;
  wire popcount27_6onj_core_096;
  wire popcount27_6onj_core_097;
  wire popcount27_6onj_core_099;
  wire popcount27_6onj_core_102;
  wire popcount27_6onj_core_104;
  wire popcount27_6onj_core_106;
  wire popcount27_6onj_core_107_not;
  wire popcount27_6onj_core_109;
  wire popcount27_6onj_core_110;
  wire popcount27_6onj_core_111;
  wire popcount27_6onj_core_112;
  wire popcount27_6onj_core_113;
  wire popcount27_6onj_core_114;
  wire popcount27_6onj_core_115;
  wire popcount27_6onj_core_116;
  wire popcount27_6onj_core_117;
  wire popcount27_6onj_core_118;
  wire popcount27_6onj_core_119;
  wire popcount27_6onj_core_120;
  wire popcount27_6onj_core_121;
  wire popcount27_6onj_core_122;
  wire popcount27_6onj_core_124;
  wire popcount27_6onj_core_126;
  wire popcount27_6onj_core_127;
  wire popcount27_6onj_core_128;
  wire popcount27_6onj_core_129;
  wire popcount27_6onj_core_130;
  wire popcount27_6onj_core_131;
  wire popcount27_6onj_core_132;
  wire popcount27_6onj_core_133;
  wire popcount27_6onj_core_135;
  wire popcount27_6onj_core_136;
  wire popcount27_6onj_core_138;
  wire popcount27_6onj_core_139;
  wire popcount27_6onj_core_143;
  wire popcount27_6onj_core_146;
  wire popcount27_6onj_core_148;
  wire popcount27_6onj_core_151_not;
  wire popcount27_6onj_core_152;
  wire popcount27_6onj_core_154;
  wire popcount27_6onj_core_156;
  wire popcount27_6onj_core_160;
  wire popcount27_6onj_core_161;
  wire popcount27_6onj_core_164;
  wire popcount27_6onj_core_165;
  wire popcount27_6onj_core_170;
  wire popcount27_6onj_core_173;
  wire popcount27_6onj_core_177;
  wire popcount27_6onj_core_178;
  wire popcount27_6onj_core_179;
  wire popcount27_6onj_core_180;
  wire popcount27_6onj_core_181;
  wire popcount27_6onj_core_182;
  wire popcount27_6onj_core_185;
  wire popcount27_6onj_core_186;
  wire popcount27_6onj_core_187;
  wire popcount27_6onj_core_188;
  wire popcount27_6onj_core_191;
  wire popcount27_6onj_core_194_not;
  wire popcount27_6onj_core_195;

  assign popcount27_6onj_core_029 = input_a[0] | input_a[15];
  assign popcount27_6onj_core_030 = input_a[3] & input_a[9];
  assign popcount27_6onj_core_031 = input_a[9] | input_a[21];
  assign popcount27_6onj_core_033 = input_a[21] & input_a[25];
  assign popcount27_6onj_core_036 = input_a[2] & input_a[22];
  assign popcount27_6onj_core_037 = input_a[15] & input_a[21];
  assign popcount27_6onj_core_038 = ~(input_a[0] & input_a[20]);
  assign popcount27_6onj_core_039 = ~input_a[22];
  assign popcount27_6onj_core_041 = input_a[13] ^ input_a[13];
  assign popcount27_6onj_core_042 = ~(input_a[0] | input_a[16]);
  assign popcount27_6onj_core_045 = input_a[20] & input_a[0];
  assign popcount27_6onj_core_046_not = ~input_a[25];
  assign popcount27_6onj_core_048 = ~(input_a[7] | input_a[25]);
  assign popcount27_6onj_core_050 = input_a[17] ^ input_a[24];
  assign popcount27_6onj_core_052 = input_a[25] | input_a[25];
  assign popcount27_6onj_core_053 = input_a[20] ^ input_a[8];
  assign popcount27_6onj_core_054 = ~(input_a[0] | input_a[15]);
  assign popcount27_6onj_core_055 = ~(input_a[13] ^ input_a[18]);
  assign popcount27_6onj_core_057 = ~(input_a[2] ^ input_a[22]);
  assign popcount27_6onj_core_058 = input_a[2] ^ input_a[15];
  assign popcount27_6onj_core_060 = input_a[11] & input_a[24];
  assign popcount27_6onj_core_061 = input_a[16] | input_a[24];
  assign popcount27_6onj_core_064 = ~input_a[17];
  assign popcount27_6onj_core_065 = input_a[22] | input_a[19];
  assign popcount27_6onj_core_066 = ~(input_a[19] | input_a[10]);
  assign popcount27_6onj_core_067 = ~(input_a[11] | input_a[0]);
  assign popcount27_6onj_core_069 = input_a[24] | input_a[20];
  assign popcount27_6onj_core_070 = ~input_a[9];
  assign popcount27_6onj_core_071 = ~(input_a[22] | input_a[3]);
  assign popcount27_6onj_core_072_not = ~input_a[3];
  assign popcount27_6onj_core_073 = ~(input_a[6] | input_a[15]);
  assign popcount27_6onj_core_074 = ~(input_a[16] ^ input_a[19]);
  assign popcount27_6onj_core_075 = input_a[6] | input_a[14];
  assign popcount27_6onj_core_076 = input_a[6] | input_a[6];
  assign popcount27_6onj_core_077 = ~(input_a[7] ^ input_a[5]);
  assign popcount27_6onj_core_078 = input_a[8] ^ input_a[10];
  assign popcount27_6onj_core_079 = ~(input_a[10] | input_a[6]);
  assign popcount27_6onj_core_082 = ~(input_a[12] | input_a[11]);
  assign popcount27_6onj_core_083_not = ~input_a[1];
  assign popcount27_6onj_core_084 = ~(input_a[2] ^ input_a[26]);
  assign popcount27_6onj_core_087 = ~(input_a[15] | input_a[9]);
  assign popcount27_6onj_core_089 = input_a[16] | input_a[20];
  assign popcount27_6onj_core_090 = ~input_a[21];
  assign popcount27_6onj_core_091 = input_a[15] & input_a[23];
  assign popcount27_6onj_core_092 = input_a[8] ^ input_a[5];
  assign popcount27_6onj_core_093 = input_a[17] & input_a[11];
  assign popcount27_6onj_core_094 = input_a[18] ^ input_a[7];
  assign popcount27_6onj_core_095 = ~(input_a[2] ^ input_a[17]);
  assign popcount27_6onj_core_096 = ~input_a[5];
  assign popcount27_6onj_core_097 = input_a[11] & input_a[19];
  assign popcount27_6onj_core_099 = input_a[3] | input_a[19];
  assign popcount27_6onj_core_102 = ~(input_a[14] | input_a[12]);
  assign popcount27_6onj_core_104 = ~input_a[7];
  assign popcount27_6onj_core_106 = ~(input_a[4] ^ input_a[6]);
  assign popcount27_6onj_core_107_not = ~input_a[26];
  assign popcount27_6onj_core_109 = input_a[26] ^ input_a[20];
  assign popcount27_6onj_core_110 = ~(input_a[17] | input_a[18]);
  assign popcount27_6onj_core_111 = input_a[22] ^ input_a[21];
  assign popcount27_6onj_core_112 = ~input_a[9];
  assign popcount27_6onj_core_113 = input_a[6] | input_a[16];
  assign popcount27_6onj_core_114 = ~input_a[25];
  assign popcount27_6onj_core_115 = ~(input_a[10] & input_a[21]);
  assign popcount27_6onj_core_116 = input_a[0] | input_a[1];
  assign popcount27_6onj_core_117 = ~(input_a[21] ^ input_a[16]);
  assign popcount27_6onj_core_118 = ~(input_a[13] | input_a[26]);
  assign popcount27_6onj_core_119 = ~(input_a[25] ^ input_a[25]);
  assign popcount27_6onj_core_120 = ~(input_a[24] ^ input_a[14]);
  assign popcount27_6onj_core_121 = input_a[22] ^ input_a[0];
  assign popcount27_6onj_core_122 = input_a[0] ^ input_a[9];
  assign popcount27_6onj_core_124 = ~(input_a[1] & input_a[7]);
  assign popcount27_6onj_core_126 = ~(input_a[5] & input_a[24]);
  assign popcount27_6onj_core_127 = input_a[23] ^ input_a[2];
  assign popcount27_6onj_core_128 = ~(input_a[10] ^ input_a[6]);
  assign popcount27_6onj_core_129 = ~(input_a[9] & input_a[2]);
  assign popcount27_6onj_core_130 = ~input_a[19];
  assign popcount27_6onj_core_131 = ~(input_a[2] & input_a[8]);
  assign popcount27_6onj_core_132 = ~(input_a[20] & input_a[20]);
  assign popcount27_6onj_core_133 = input_a[17] ^ input_a[11];
  assign popcount27_6onj_core_135 = input_a[8] & input_a[20];
  assign popcount27_6onj_core_136 = ~(input_a[26] | input_a[9]);
  assign popcount27_6onj_core_138 = ~(input_a[10] ^ input_a[12]);
  assign popcount27_6onj_core_139 = ~(input_a[16] ^ input_a[19]);
  assign popcount27_6onj_core_143 = input_a[23] & input_a[19];
  assign popcount27_6onj_core_146 = input_a[16] & input_a[5];
  assign popcount27_6onj_core_148 = ~input_a[24];
  assign popcount27_6onj_core_151_not = ~input_a[17];
  assign popcount27_6onj_core_152 = ~input_a[1];
  assign popcount27_6onj_core_154 = input_a[8] ^ input_a[4];
  assign popcount27_6onj_core_156 = input_a[8] | input_a[5];
  assign popcount27_6onj_core_160 = input_a[10] ^ input_a[16];
  assign popcount27_6onj_core_161 = ~(input_a[16] | input_a[2]);
  assign popcount27_6onj_core_164 = ~(input_a[13] | input_a[13]);
  assign popcount27_6onj_core_165 = input_a[25] | input_a[15];
  assign popcount27_6onj_core_170 = input_a[24] & input_a[19];
  assign popcount27_6onj_core_173 = input_a[16] & input_a[4];
  assign popcount27_6onj_core_177 = ~(input_a[9] & input_a[15]);
  assign popcount27_6onj_core_178 = ~(input_a[16] & input_a[25]);
  assign popcount27_6onj_core_179 = ~(input_a[18] ^ input_a[18]);
  assign popcount27_6onj_core_180 = ~(input_a[23] | input_a[17]);
  assign popcount27_6onj_core_181 = ~input_a[14];
  assign popcount27_6onj_core_182 = ~(input_a[0] ^ input_a[12]);
  assign popcount27_6onj_core_185 = input_a[13] & input_a[16];
  assign popcount27_6onj_core_186 = ~(input_a[23] | input_a[8]);
  assign popcount27_6onj_core_187 = ~(input_a[24] ^ input_a[25]);
  assign popcount27_6onj_core_188 = ~(input_a[0] & input_a[20]);
  assign popcount27_6onj_core_191 = input_a[19] | input_a[11];
  assign popcount27_6onj_core_194_not = ~input_a[11];
  assign popcount27_6onj_core_195 = ~input_a[26];

  assign popcount27_6onj_out[0] = 1'b0;
  assign popcount27_6onj_out[1] = 1'b0;
  assign popcount27_6onj_out[2] = popcount27_6onj_core_188;
  assign popcount27_6onj_out[3] = popcount27_6onj_core_188;
  assign popcount27_6onj_out[4] = popcount27_6onj_core_045;
endmodule