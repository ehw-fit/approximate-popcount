// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.69417
// WCE=21.0
// EP=0.953061%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_to1t(input [30:0] input_a, output [4:0] popcount31_to1t_out);
  wire popcount31_to1t_core_036;
  wire popcount31_to1t_core_038;
  wire popcount31_to1t_core_039;
  wire popcount31_to1t_core_041;
  wire popcount31_to1t_core_043;
  wire popcount31_to1t_core_045_not;
  wire popcount31_to1t_core_046;
  wire popcount31_to1t_core_050;
  wire popcount31_to1t_core_052;
  wire popcount31_to1t_core_053;
  wire popcount31_to1t_core_054;
  wire popcount31_to1t_core_057;
  wire popcount31_to1t_core_059;
  wire popcount31_to1t_core_060;
  wire popcount31_to1t_core_063;
  wire popcount31_to1t_core_064;
  wire popcount31_to1t_core_065;
  wire popcount31_to1t_core_067;
  wire popcount31_to1t_core_068;
  wire popcount31_to1t_core_069;
  wire popcount31_to1t_core_070;
  wire popcount31_to1t_core_071;
  wire popcount31_to1t_core_073;
  wire popcount31_to1t_core_074;
  wire popcount31_to1t_core_075;
  wire popcount31_to1t_core_076;
  wire popcount31_to1t_core_077;
  wire popcount31_to1t_core_079;
  wire popcount31_to1t_core_080;
  wire popcount31_to1t_core_082;
  wire popcount31_to1t_core_086;
  wire popcount31_to1t_core_088;
  wire popcount31_to1t_core_093;
  wire popcount31_to1t_core_095;
  wire popcount31_to1t_core_096;
  wire popcount31_to1t_core_097;
  wire popcount31_to1t_core_098;
  wire popcount31_to1t_core_099;
  wire popcount31_to1t_core_100;
  wire popcount31_to1t_core_102;
  wire popcount31_to1t_core_104;
  wire popcount31_to1t_core_106;
  wire popcount31_to1t_core_107;
  wire popcount31_to1t_core_115;
  wire popcount31_to1t_core_116;
  wire popcount31_to1t_core_120;
  wire popcount31_to1t_core_121;
  wire popcount31_to1t_core_129;
  wire popcount31_to1t_core_133;
  wire popcount31_to1t_core_134;
  wire popcount31_to1t_core_136;
  wire popcount31_to1t_core_138;
  wire popcount31_to1t_core_139;
  wire popcount31_to1t_core_140;
  wire popcount31_to1t_core_142;
  wire popcount31_to1t_core_143;
  wire popcount31_to1t_core_144;
  wire popcount31_to1t_core_145;
  wire popcount31_to1t_core_146;
  wire popcount31_to1t_core_147;
  wire popcount31_to1t_core_150;
  wire popcount31_to1t_core_151;
  wire popcount31_to1t_core_153;
  wire popcount31_to1t_core_156;
  wire popcount31_to1t_core_158;
  wire popcount31_to1t_core_159;
  wire popcount31_to1t_core_160;
  wire popcount31_to1t_core_161;
  wire popcount31_to1t_core_162;
  wire popcount31_to1t_core_164;
  wire popcount31_to1t_core_166;
  wire popcount31_to1t_core_167;
  wire popcount31_to1t_core_172;
  wire popcount31_to1t_core_173;
  wire popcount31_to1t_core_174;
  wire popcount31_to1t_core_175;
  wire popcount31_to1t_core_177;
  wire popcount31_to1t_core_178;
  wire popcount31_to1t_core_180;
  wire popcount31_to1t_core_181;
  wire popcount31_to1t_core_183;
  wire popcount31_to1t_core_184;
  wire popcount31_to1t_core_186;
  wire popcount31_to1t_core_187;
  wire popcount31_to1t_core_188;
  wire popcount31_to1t_core_189;
  wire popcount31_to1t_core_190;
  wire popcount31_to1t_core_191;
  wire popcount31_to1t_core_192;
  wire popcount31_to1t_core_193;
  wire popcount31_to1t_core_194;
  wire popcount31_to1t_core_195;
  wire popcount31_to1t_core_196;
  wire popcount31_to1t_core_197;
  wire popcount31_to1t_core_200;
  wire popcount31_to1t_core_201_not;
  wire popcount31_to1t_core_203;
  wire popcount31_to1t_core_205;
  wire popcount31_to1t_core_206;
  wire popcount31_to1t_core_207;
  wire popcount31_to1t_core_210;
  wire popcount31_to1t_core_211;
  wire popcount31_to1t_core_213;
  wire popcount31_to1t_core_214;
  wire popcount31_to1t_core_215;
  wire popcount31_to1t_core_218;
  wire popcount31_to1t_core_219;

  assign popcount31_to1t_core_036 = input_a[8] ^ input_a[14];
  assign popcount31_to1t_core_038 = ~(input_a[15] | input_a[2]);
  assign popcount31_to1t_core_039 = ~input_a[9];
  assign popcount31_to1t_core_041 = ~(input_a[22] | input_a[14]);
  assign popcount31_to1t_core_043 = ~(input_a[24] ^ input_a[30]);
  assign popcount31_to1t_core_045_not = ~input_a[8];
  assign popcount31_to1t_core_046 = ~(input_a[23] | input_a[30]);
  assign popcount31_to1t_core_050 = ~(input_a[4] ^ input_a[1]);
  assign popcount31_to1t_core_052 = input_a[27] ^ input_a[24];
  assign popcount31_to1t_core_053 = ~(input_a[22] ^ input_a[9]);
  assign popcount31_to1t_core_054 = input_a[23] & input_a[25];
  assign popcount31_to1t_core_057 = ~(input_a[17] ^ input_a[29]);
  assign popcount31_to1t_core_059 = ~(input_a[28] | input_a[28]);
  assign popcount31_to1t_core_060 = ~(input_a[23] | input_a[18]);
  assign popcount31_to1t_core_063 = input_a[2] ^ input_a[30];
  assign popcount31_to1t_core_064 = ~(input_a[5] ^ input_a[19]);
  assign popcount31_to1t_core_065 = input_a[25] ^ input_a[23];
  assign popcount31_to1t_core_067 = input_a[19] ^ input_a[0];
  assign popcount31_to1t_core_068 = input_a[0] | input_a[14];
  assign popcount31_to1t_core_069 = input_a[17] ^ input_a[30];
  assign popcount31_to1t_core_070 = ~(input_a[12] | input_a[17]);
  assign popcount31_to1t_core_071 = input_a[11] ^ input_a[26];
  assign popcount31_to1t_core_073 = ~(input_a[18] & input_a[22]);
  assign popcount31_to1t_core_074 = ~(input_a[2] | input_a[15]);
  assign popcount31_to1t_core_075 = input_a[20] ^ input_a[6];
  assign popcount31_to1t_core_076 = ~(input_a[12] & input_a[18]);
  assign popcount31_to1t_core_077 = input_a[25] & input_a[6];
  assign popcount31_to1t_core_079 = ~(input_a[9] & input_a[0]);
  assign popcount31_to1t_core_080 = ~(input_a[12] & input_a[10]);
  assign popcount31_to1t_core_082 = input_a[10] ^ input_a[10];
  assign popcount31_to1t_core_086 = ~(input_a[15] & input_a[24]);
  assign popcount31_to1t_core_088 = ~(input_a[2] & input_a[11]);
  assign popcount31_to1t_core_093 = ~(input_a[12] ^ input_a[0]);
  assign popcount31_to1t_core_095 = ~(input_a[5] ^ input_a[29]);
  assign popcount31_to1t_core_096 = input_a[16] & input_a[8];
  assign popcount31_to1t_core_097 = ~(input_a[0] | input_a[22]);
  assign popcount31_to1t_core_098 = input_a[30] ^ input_a[3];
  assign popcount31_to1t_core_099 = ~input_a[9];
  assign popcount31_to1t_core_100 = ~(input_a[22] | input_a[22]);
  assign popcount31_to1t_core_102 = ~input_a[20];
  assign popcount31_to1t_core_104 = ~(input_a[21] ^ input_a[4]);
  assign popcount31_to1t_core_106 = input_a[5] | input_a[18];
  assign popcount31_to1t_core_107 = ~(input_a[13] & input_a[10]);
  assign popcount31_to1t_core_115 = ~(input_a[28] | input_a[28]);
  assign popcount31_to1t_core_116 = input_a[11] | input_a[15];
  assign popcount31_to1t_core_120 = input_a[27] | input_a[25];
  assign popcount31_to1t_core_121 = ~input_a[10];
  assign popcount31_to1t_core_129 = input_a[30] & input_a[11];
  assign popcount31_to1t_core_133 = input_a[10] | input_a[5];
  assign popcount31_to1t_core_134 = input_a[10] & input_a[16];
  assign popcount31_to1t_core_136 = ~(input_a[10] ^ input_a[30]);
  assign popcount31_to1t_core_138 = input_a[12] & input_a[19];
  assign popcount31_to1t_core_139 = input_a[20] ^ input_a[14];
  assign popcount31_to1t_core_140 = ~(input_a[26] | input_a[2]);
  assign popcount31_to1t_core_142 = ~(input_a[30] & input_a[21]);
  assign popcount31_to1t_core_143 = input_a[27] | input_a[30];
  assign popcount31_to1t_core_144 = input_a[17] | input_a[18];
  assign popcount31_to1t_core_145 = ~(input_a[9] | input_a[18]);
  assign popcount31_to1t_core_146 = input_a[18] ^ input_a[22];
  assign popcount31_to1t_core_147 = input_a[4] | input_a[6];
  assign popcount31_to1t_core_150 = ~(input_a[12] ^ input_a[20]);
  assign popcount31_to1t_core_151 = ~(input_a[29] ^ input_a[2]);
  assign popcount31_to1t_core_153 = ~(input_a[22] | input_a[1]);
  assign popcount31_to1t_core_156 = ~(input_a[18] & input_a[26]);
  assign popcount31_to1t_core_158 = input_a[11] ^ input_a[26];
  assign popcount31_to1t_core_159 = input_a[22] | input_a[14];
  assign popcount31_to1t_core_160 = input_a[20] ^ input_a[11];
  assign popcount31_to1t_core_161 = ~(input_a[25] | input_a[7]);
  assign popcount31_to1t_core_162 = input_a[8] & input_a[27];
  assign popcount31_to1t_core_164 = ~input_a[0];
  assign popcount31_to1t_core_166 = input_a[10] & input_a[20];
  assign popcount31_to1t_core_167 = input_a[30] ^ input_a[17];
  assign popcount31_to1t_core_172 = ~(input_a[4] & input_a[6]);
  assign popcount31_to1t_core_173 = ~(input_a[8] ^ input_a[28]);
  assign popcount31_to1t_core_174 = ~(input_a[21] | input_a[3]);
  assign popcount31_to1t_core_175 = ~(input_a[19] | input_a[6]);
  assign popcount31_to1t_core_177 = input_a[13] ^ input_a[1];
  assign popcount31_to1t_core_178 = input_a[15] & input_a[28];
  assign popcount31_to1t_core_180 = ~input_a[6];
  assign popcount31_to1t_core_181 = input_a[18] & input_a[0];
  assign popcount31_to1t_core_183 = input_a[0] & input_a[27];
  assign popcount31_to1t_core_184 = ~(input_a[20] & input_a[5]);
  assign popcount31_to1t_core_186 = input_a[6] & input_a[15];
  assign popcount31_to1t_core_187 = input_a[9] & input_a[23];
  assign popcount31_to1t_core_188 = input_a[0] & input_a[7];
  assign popcount31_to1t_core_189 = ~input_a[1];
  assign popcount31_to1t_core_190 = ~(input_a[7] & input_a[28]);
  assign popcount31_to1t_core_191 = input_a[12] | input_a[11];
  assign popcount31_to1t_core_192 = ~(input_a[25] | input_a[4]);
  assign popcount31_to1t_core_193 = input_a[9] & input_a[2];
  assign popcount31_to1t_core_194 = ~(input_a[14] | input_a[5]);
  assign popcount31_to1t_core_195 = ~(input_a[22] ^ input_a[30]);
  assign popcount31_to1t_core_196 = input_a[9] | input_a[17];
  assign popcount31_to1t_core_197 = input_a[7] | input_a[11];
  assign popcount31_to1t_core_200 = ~input_a[26];
  assign popcount31_to1t_core_201_not = ~input_a[28];
  assign popcount31_to1t_core_203 = ~(input_a[11] & input_a[7]);
  assign popcount31_to1t_core_205 = ~(input_a[3] | input_a[29]);
  assign popcount31_to1t_core_206 = input_a[26] ^ input_a[15];
  assign popcount31_to1t_core_207 = input_a[8] & input_a[12];
  assign popcount31_to1t_core_210 = ~input_a[25];
  assign popcount31_to1t_core_211 = ~input_a[14];
  assign popcount31_to1t_core_213 = input_a[13] ^ input_a[23];
  assign popcount31_to1t_core_214 = ~input_a[21];
  assign popcount31_to1t_core_215 = input_a[25] | input_a[0];
  assign popcount31_to1t_core_218 = input_a[23] | input_a[9];
  assign popcount31_to1t_core_219 = ~(input_a[23] ^ input_a[30]);

  assign popcount31_to1t_out[0] = 1'b0;
  assign popcount31_to1t_out[1] = input_a[1];
  assign popcount31_to1t_out[2] = input_a[23];
  assign popcount31_to1t_out[3] = 1'b1;
  assign popcount31_to1t_out[4] = 1'b0;
endmodule