// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.48658
// WCE=11.0
// EP=0.790412%
// Printed PDK parameters:
//  Area=45176751.0
//  Delay=69366280.0
//  Power=2540700.0

module popcount30_lnxq(input [29:0] input_a, output [4:0] popcount30_lnxq_out);
  wire popcount30_lnxq_core_032;
  wire popcount30_lnxq_core_033;
  wire popcount30_lnxq_core_035;
  wire popcount30_lnxq_core_036;
  wire popcount30_lnxq_core_037;
  wire popcount30_lnxq_core_038;
  wire popcount30_lnxq_core_039;
  wire popcount30_lnxq_core_040;
  wire popcount30_lnxq_core_041;
  wire popcount30_lnxq_core_044;
  wire popcount30_lnxq_core_045;
  wire popcount30_lnxq_core_047;
  wire popcount30_lnxq_core_048;
  wire popcount30_lnxq_core_051;
  wire popcount30_lnxq_core_052;
  wire popcount30_lnxq_core_054;
  wire popcount30_lnxq_core_057_not;
  wire popcount30_lnxq_core_058;
  wire popcount30_lnxq_core_059;
  wire popcount30_lnxq_core_062;
  wire popcount30_lnxq_core_063;
  wire popcount30_lnxq_core_064;
  wire popcount30_lnxq_core_067;
  wire popcount30_lnxq_core_068;
  wire popcount30_lnxq_core_069;
  wire popcount30_lnxq_core_070;
  wire popcount30_lnxq_core_071;
  wire popcount30_lnxq_core_072;
  wire popcount30_lnxq_core_075;
  wire popcount30_lnxq_core_076;
  wire popcount30_lnxq_core_078;
  wire popcount30_lnxq_core_079;
  wire popcount30_lnxq_core_080;
  wire popcount30_lnxq_core_081;
  wire popcount30_lnxq_core_083;
  wire popcount30_lnxq_core_084;
  wire popcount30_lnxq_core_085;
  wire popcount30_lnxq_core_086;
  wire popcount30_lnxq_core_087;
  wire popcount30_lnxq_core_088;
  wire popcount30_lnxq_core_089;
  wire popcount30_lnxq_core_090;
  wire popcount30_lnxq_core_091;
  wire popcount30_lnxq_core_092;
  wire popcount30_lnxq_core_093;
  wire popcount30_lnxq_core_094;
  wire popcount30_lnxq_core_096;
  wire popcount30_lnxq_core_097;
  wire popcount30_lnxq_core_098;
  wire popcount30_lnxq_core_099;
  wire popcount30_lnxq_core_100;
  wire popcount30_lnxq_core_101;
  wire popcount30_lnxq_core_102;
  wire popcount30_lnxq_core_103;
  wire popcount30_lnxq_core_104;
  wire popcount30_lnxq_core_105;
  wire popcount30_lnxq_core_106;
  wire popcount30_lnxq_core_108;
  wire popcount30_lnxq_core_109;
  wire popcount30_lnxq_core_111;
  wire popcount30_lnxq_core_112;
  wire popcount30_lnxq_core_113;
  wire popcount30_lnxq_core_114;
  wire popcount30_lnxq_core_115;
  wire popcount30_lnxq_core_118;
  wire popcount30_lnxq_core_120;
  wire popcount30_lnxq_core_121;
  wire popcount30_lnxq_core_122;
  wire popcount30_lnxq_core_124;
  wire popcount30_lnxq_core_126;
  wire popcount30_lnxq_core_127;
  wire popcount30_lnxq_core_128;
  wire popcount30_lnxq_core_129;
  wire popcount30_lnxq_core_130;
  wire popcount30_lnxq_core_131_not;
  wire popcount30_lnxq_core_133;
  wire popcount30_lnxq_core_134;
  wire popcount30_lnxq_core_136;
  wire popcount30_lnxq_core_137;
  wire popcount30_lnxq_core_138;
  wire popcount30_lnxq_core_143;
  wire popcount30_lnxq_core_144;
  wire popcount30_lnxq_core_146;
  wire popcount30_lnxq_core_147;
  wire popcount30_lnxq_core_148;
  wire popcount30_lnxq_core_152;
  wire popcount30_lnxq_core_153;
  wire popcount30_lnxq_core_156;
  wire popcount30_lnxq_core_157;
  wire popcount30_lnxq_core_158;
  wire popcount30_lnxq_core_159;
  wire popcount30_lnxq_core_160;
  wire popcount30_lnxq_core_161;
  wire popcount30_lnxq_core_162;
  wire popcount30_lnxq_core_164;
  wire popcount30_lnxq_core_165;
  wire popcount30_lnxq_core_166;
  wire popcount30_lnxq_core_169;
  wire popcount30_lnxq_core_170;
  wire popcount30_lnxq_core_172;
  wire popcount30_lnxq_core_173;
  wire popcount30_lnxq_core_174;
  wire popcount30_lnxq_core_176;
  wire popcount30_lnxq_core_177;
  wire popcount30_lnxq_core_178;
  wire popcount30_lnxq_core_179;
  wire popcount30_lnxq_core_180;
  wire popcount30_lnxq_core_181;
  wire popcount30_lnxq_core_182;
  wire popcount30_lnxq_core_183;
  wire popcount30_lnxq_core_184;
  wire popcount30_lnxq_core_185;
  wire popcount30_lnxq_core_186;
  wire popcount30_lnxq_core_188;
  wire popcount30_lnxq_core_194;
  wire popcount30_lnxq_core_195;
  wire popcount30_lnxq_core_197;
  wire popcount30_lnxq_core_199;
  wire popcount30_lnxq_core_200;
  wire popcount30_lnxq_core_201;
  wire popcount30_lnxq_core_202;
  wire popcount30_lnxq_core_203;
  wire popcount30_lnxq_core_204;
  wire popcount30_lnxq_core_205;
  wire popcount30_lnxq_core_206;
  wire popcount30_lnxq_core_207;
  wire popcount30_lnxq_core_208;
  wire popcount30_lnxq_core_210;
  wire popcount30_lnxq_core_211;
  wire popcount30_lnxq_core_212;

  assign popcount30_lnxq_core_032 = input_a[13] | input_a[6];
  assign popcount30_lnxq_core_033 = input_a[28] & input_a[27];
  assign popcount30_lnxq_core_035 = input_a[4] & input_a[25];
  assign popcount30_lnxq_core_036 = popcount30_lnxq_core_033 ^ popcount30_lnxq_core_035;
  assign popcount30_lnxq_core_037 = popcount30_lnxq_core_033 & popcount30_lnxq_core_035;
  assign popcount30_lnxq_core_038 = input_a[26] & input_a[18];
  assign popcount30_lnxq_core_039 = input_a[22] & input_a[26];
  assign popcount30_lnxq_core_040 = input_a[29] & input_a[6];
  assign popcount30_lnxq_core_041 = input_a[19] & input_a[6];
  assign popcount30_lnxq_core_044 = popcount30_lnxq_core_039 | popcount30_lnxq_core_041;
  assign popcount30_lnxq_core_045 = ~(input_a[8] | input_a[15]);
  assign popcount30_lnxq_core_047 = input_a[17] ^ input_a[22];
  assign popcount30_lnxq_core_048 = ~(input_a[6] ^ input_a[22]);
  assign popcount30_lnxq_core_051 = popcount30_lnxq_core_036 ^ popcount30_lnxq_core_044;
  assign popcount30_lnxq_core_052 = popcount30_lnxq_core_036 & popcount30_lnxq_core_044;
  assign popcount30_lnxq_core_054 = ~input_a[24];
  assign popcount30_lnxq_core_057_not = ~input_a[5];
  assign popcount30_lnxq_core_058 = popcount30_lnxq_core_037 | popcount30_lnxq_core_052;
  assign popcount30_lnxq_core_059 = ~(input_a[2] | input_a[29]);
  assign popcount30_lnxq_core_062 = input_a[18] & input_a[3];
  assign popcount30_lnxq_core_063 = input_a[9] ^ input_a[10];
  assign popcount30_lnxq_core_064 = input_a[9] & input_a[10];
  assign popcount30_lnxq_core_067 = popcount30_lnxq_core_062 ^ popcount30_lnxq_core_064;
  assign popcount30_lnxq_core_068 = popcount30_lnxq_core_062 & input_a[9];
  assign popcount30_lnxq_core_069 = popcount30_lnxq_core_067 ^ popcount30_lnxq_core_063;
  assign popcount30_lnxq_core_070 = popcount30_lnxq_core_067 & popcount30_lnxq_core_063;
  assign popcount30_lnxq_core_071 = popcount30_lnxq_core_068 | popcount30_lnxq_core_070;
  assign popcount30_lnxq_core_072 = input_a[12] ^ input_a[16];
  assign popcount30_lnxq_core_075 = input_a[17] & input_a[5];
  assign popcount30_lnxq_core_076 = input_a[8] | input_a[5];
  assign popcount30_lnxq_core_078 = input_a[11] ^ popcount30_lnxq_core_075;
  assign popcount30_lnxq_core_079 = input_a[11] & popcount30_lnxq_core_075;
  assign popcount30_lnxq_core_080 = popcount30_lnxq_core_078 | input_a[1];
  assign popcount30_lnxq_core_081 = input_a[9] & input_a[21];
  assign popcount30_lnxq_core_083 = input_a[26] & input_a[25];
  assign popcount30_lnxq_core_084 = input_a[0] & input_a[12];
  assign popcount30_lnxq_core_085 = popcount30_lnxq_core_069 ^ popcount30_lnxq_core_080;
  assign popcount30_lnxq_core_086 = popcount30_lnxq_core_069 & popcount30_lnxq_core_080;
  assign popcount30_lnxq_core_087 = popcount30_lnxq_core_085 ^ popcount30_lnxq_core_084;
  assign popcount30_lnxq_core_088 = popcount30_lnxq_core_085 & popcount30_lnxq_core_084;
  assign popcount30_lnxq_core_089 = popcount30_lnxq_core_086 | popcount30_lnxq_core_088;
  assign popcount30_lnxq_core_090 = popcount30_lnxq_core_071 ^ popcount30_lnxq_core_079;
  assign popcount30_lnxq_core_091 = popcount30_lnxq_core_071 & popcount30_lnxq_core_079;
  assign popcount30_lnxq_core_092 = popcount30_lnxq_core_090 ^ popcount30_lnxq_core_089;
  assign popcount30_lnxq_core_093 = popcount30_lnxq_core_090 & popcount30_lnxq_core_089;
  assign popcount30_lnxq_core_094 = popcount30_lnxq_core_091 | popcount30_lnxq_core_093;
  assign popcount30_lnxq_core_096 = input_a[23] & input_a[13];
  assign popcount30_lnxq_core_097 = popcount30_lnxq_core_051 ^ popcount30_lnxq_core_087;
  assign popcount30_lnxq_core_098 = popcount30_lnxq_core_051 & popcount30_lnxq_core_087;
  assign popcount30_lnxq_core_099 = popcount30_lnxq_core_097 ^ popcount30_lnxq_core_096;
  assign popcount30_lnxq_core_100 = popcount30_lnxq_core_097 & popcount30_lnxq_core_096;
  assign popcount30_lnxq_core_101 = popcount30_lnxq_core_098 | popcount30_lnxq_core_100;
  assign popcount30_lnxq_core_102 = popcount30_lnxq_core_058 ^ popcount30_lnxq_core_092;
  assign popcount30_lnxq_core_103 = popcount30_lnxq_core_058 & popcount30_lnxq_core_092;
  assign popcount30_lnxq_core_104 = popcount30_lnxq_core_102 ^ popcount30_lnxq_core_101;
  assign popcount30_lnxq_core_105 = popcount30_lnxq_core_102 & popcount30_lnxq_core_101;
  assign popcount30_lnxq_core_106 = popcount30_lnxq_core_103 | popcount30_lnxq_core_105;
  assign popcount30_lnxq_core_108 = input_a[27] ^ input_a[19];
  assign popcount30_lnxq_core_109 = popcount30_lnxq_core_094 | popcount30_lnxq_core_106;
  assign popcount30_lnxq_core_111 = ~(input_a[5] & input_a[8]);
  assign popcount30_lnxq_core_112 = ~input_a[17];
  assign popcount30_lnxq_core_113 = ~(input_a[18] ^ input_a[1]);
  assign popcount30_lnxq_core_114 = ~input_a[26];
  assign popcount30_lnxq_core_115 = input_a[14] | input_a[20];
  assign popcount30_lnxq_core_118 = input_a[7] ^ input_a[2];
  assign popcount30_lnxq_core_120 = ~(input_a[20] & input_a[21]);
  assign popcount30_lnxq_core_121 = input_a[20] & input_a[21];
  assign popcount30_lnxq_core_122 = popcount30_lnxq_core_118 ^ popcount30_lnxq_core_120;
  assign popcount30_lnxq_core_124 = input_a[2] ^ popcount30_lnxq_core_121;
  assign popcount30_lnxq_core_126 = popcount30_lnxq_core_124 | popcount30_lnxq_core_118;
  assign popcount30_lnxq_core_127 = ~(input_a[6] ^ input_a[4]);
  assign popcount30_lnxq_core_128 = ~(input_a[18] & input_a[11]);
  assign popcount30_lnxq_core_129 = ~(input_a[17] | input_a[21]);
  assign popcount30_lnxq_core_130 = input_a[15] & popcount30_lnxq_core_122;
  assign popcount30_lnxq_core_131_not = ~popcount30_lnxq_core_126;
  assign popcount30_lnxq_core_133 = popcount30_lnxq_core_131_not ^ popcount30_lnxq_core_130;
  assign popcount30_lnxq_core_134 = ~(input_a[27] ^ input_a[20]);
  assign popcount30_lnxq_core_136 = input_a[15] | input_a[7];
  assign popcount30_lnxq_core_137 = ~(input_a[19] & input_a[27]);
  assign popcount30_lnxq_core_138 = popcount30_lnxq_core_136 | popcount30_lnxq_core_126;
  assign popcount30_lnxq_core_143 = ~input_a[5];
  assign popcount30_lnxq_core_144 = ~(input_a[18] & input_a[18]);
  assign popcount30_lnxq_core_146 = ~input_a[19];
  assign popcount30_lnxq_core_147 = ~(input_a[4] | input_a[29]);
  assign popcount30_lnxq_core_148 = input_a[20] | input_a[19];
  assign popcount30_lnxq_core_152 = ~(input_a[4] | input_a[25]);
  assign popcount30_lnxq_core_153 = ~(input_a[15] | input_a[16]);
  assign popcount30_lnxq_core_156 = ~(input_a[13] & input_a[0]);
  assign popcount30_lnxq_core_157 = ~(input_a[1] ^ input_a[1]);
  assign popcount30_lnxq_core_158 = ~(input_a[3] | input_a[10]);
  assign popcount30_lnxq_core_159 = ~(input_a[11] | input_a[18]);
  assign popcount30_lnxq_core_160 = ~(input_a[11] & input_a[8]);
  assign popcount30_lnxq_core_161 = input_a[8] ^ input_a[7];
  assign popcount30_lnxq_core_162 = input_a[19] | input_a[5];
  assign popcount30_lnxq_core_164 = ~(input_a[16] | input_a[23]);
  assign popcount30_lnxq_core_165 = ~input_a[29];
  assign popcount30_lnxq_core_166 = ~(input_a[15] | input_a[8]);
  assign popcount30_lnxq_core_169 = input_a[10] & input_a[27];
  assign popcount30_lnxq_core_170 = ~(input_a[21] | input_a[21]);
  assign popcount30_lnxq_core_172 = input_a[10] | input_a[25];
  assign popcount30_lnxq_core_173 = input_a[9] ^ input_a[5];
  assign popcount30_lnxq_core_174 = input_a[27] ^ input_a[1];
  assign popcount30_lnxq_core_176 = input_a[8] & input_a[14];
  assign popcount30_lnxq_core_177 = popcount30_lnxq_core_133 ^ popcount30_lnxq_core_165;
  assign popcount30_lnxq_core_178 = popcount30_lnxq_core_133 & popcount30_lnxq_core_165;
  assign popcount30_lnxq_core_179 = popcount30_lnxq_core_177 ^ popcount30_lnxq_core_176;
  assign popcount30_lnxq_core_180 = popcount30_lnxq_core_177 & popcount30_lnxq_core_176;
  assign popcount30_lnxq_core_181 = popcount30_lnxq_core_178 | popcount30_lnxq_core_180;
  assign popcount30_lnxq_core_182 = popcount30_lnxq_core_138 ^ input_a[29];
  assign popcount30_lnxq_core_183 = popcount30_lnxq_core_138 & input_a[29];
  assign popcount30_lnxq_core_184 = popcount30_lnxq_core_182 ^ popcount30_lnxq_core_181;
  assign popcount30_lnxq_core_185 = popcount30_lnxq_core_182 & popcount30_lnxq_core_181;
  assign popcount30_lnxq_core_186 = popcount30_lnxq_core_183 | popcount30_lnxq_core_185;
  assign popcount30_lnxq_core_188 = ~(input_a[17] ^ input_a[6]);
  assign popcount30_lnxq_core_194 = popcount30_lnxq_core_099 ^ popcount30_lnxq_core_179;
  assign popcount30_lnxq_core_195 = popcount30_lnxq_core_099 & popcount30_lnxq_core_179;
  assign popcount30_lnxq_core_197 = input_a[2] & input_a[28];
  assign popcount30_lnxq_core_199 = popcount30_lnxq_core_104 ^ popcount30_lnxq_core_184;
  assign popcount30_lnxq_core_200 = popcount30_lnxq_core_104 & popcount30_lnxq_core_184;
  assign popcount30_lnxq_core_201 = popcount30_lnxq_core_199 ^ popcount30_lnxq_core_195;
  assign popcount30_lnxq_core_202 = popcount30_lnxq_core_199 & popcount30_lnxq_core_195;
  assign popcount30_lnxq_core_203 = popcount30_lnxq_core_200 | popcount30_lnxq_core_202;
  assign popcount30_lnxq_core_204 = popcount30_lnxq_core_109 ^ popcount30_lnxq_core_186;
  assign popcount30_lnxq_core_205 = popcount30_lnxq_core_109 & popcount30_lnxq_core_186;
  assign popcount30_lnxq_core_206 = popcount30_lnxq_core_204 ^ popcount30_lnxq_core_203;
  assign popcount30_lnxq_core_207 = popcount30_lnxq_core_204 & popcount30_lnxq_core_203;
  assign popcount30_lnxq_core_208 = popcount30_lnxq_core_205 | popcount30_lnxq_core_207;
  assign popcount30_lnxq_core_210 = ~(input_a[2] | input_a[1]);
  assign popcount30_lnxq_core_211 = ~(input_a[26] & input_a[2]);
  assign popcount30_lnxq_core_212 = ~input_a[14];

  assign popcount30_lnxq_out[0] = popcount30_lnxq_core_206;
  assign popcount30_lnxq_out[1] = popcount30_lnxq_core_194;
  assign popcount30_lnxq_out[2] = popcount30_lnxq_core_201;
  assign popcount30_lnxq_out[3] = popcount30_lnxq_core_206;
  assign popcount30_lnxq_out[4] = popcount30_lnxq_core_208;
endmodule