// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.25652
// WCE=13.0
// EP=0.863617%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_bpx5(input [22:0] input_a, output [4:0] popcount23_bpx5_out);
  wire popcount23_bpx5_core_026;
  wire popcount23_bpx5_core_027;
  wire popcount23_bpx5_core_028;
  wire popcount23_bpx5_core_029;
  wire popcount23_bpx5_core_030;
  wire popcount23_bpx5_core_031;
  wire popcount23_bpx5_core_033;
  wire popcount23_bpx5_core_035;
  wire popcount23_bpx5_core_036;
  wire popcount23_bpx5_core_038;
  wire popcount23_bpx5_core_040;
  wire popcount23_bpx5_core_042;
  wire popcount23_bpx5_core_043;
  wire popcount23_bpx5_core_044_not;
  wire popcount23_bpx5_core_047;
  wire popcount23_bpx5_core_048;
  wire popcount23_bpx5_core_049;
  wire popcount23_bpx5_core_052;
  wire popcount23_bpx5_core_056;
  wire popcount23_bpx5_core_058;
  wire popcount23_bpx5_core_059;
  wire popcount23_bpx5_core_061;
  wire popcount23_bpx5_core_063;
  wire popcount23_bpx5_core_065_not;
  wire popcount23_bpx5_core_066;
  wire popcount23_bpx5_core_067;
  wire popcount23_bpx5_core_069;
  wire popcount23_bpx5_core_070;
  wire popcount23_bpx5_core_071;
  wire popcount23_bpx5_core_072_not;
  wire popcount23_bpx5_core_073;
  wire popcount23_bpx5_core_074;
  wire popcount23_bpx5_core_075;
  wire popcount23_bpx5_core_076;
  wire popcount23_bpx5_core_077;
  wire popcount23_bpx5_core_078;
  wire popcount23_bpx5_core_081;
  wire popcount23_bpx5_core_084;
  wire popcount23_bpx5_core_085;
  wire popcount23_bpx5_core_086;
  wire popcount23_bpx5_core_087;
  wire popcount23_bpx5_core_090;
  wire popcount23_bpx5_core_093_not;
  wire popcount23_bpx5_core_094;
  wire popcount23_bpx5_core_095;
  wire popcount23_bpx5_core_096;
  wire popcount23_bpx5_core_097;
  wire popcount23_bpx5_core_098;
  wire popcount23_bpx5_core_100;
  wire popcount23_bpx5_core_101;
  wire popcount23_bpx5_core_102;
  wire popcount23_bpx5_core_104;
  wire popcount23_bpx5_core_107;
  wire popcount23_bpx5_core_110;
  wire popcount23_bpx5_core_111;
  wire popcount23_bpx5_core_112;
  wire popcount23_bpx5_core_114;
  wire popcount23_bpx5_core_120;
  wire popcount23_bpx5_core_122;
  wire popcount23_bpx5_core_123;
  wire popcount23_bpx5_core_125;
  wire popcount23_bpx5_core_126;
  wire popcount23_bpx5_core_127;
  wire popcount23_bpx5_core_130;
  wire popcount23_bpx5_core_131;
  wire popcount23_bpx5_core_133;
  wire popcount23_bpx5_core_134;
  wire popcount23_bpx5_core_135;
  wire popcount23_bpx5_core_136;
  wire popcount23_bpx5_core_138;
  wire popcount23_bpx5_core_139;
  wire popcount23_bpx5_core_141;
  wire popcount23_bpx5_core_143;
  wire popcount23_bpx5_core_145;
  wire popcount23_bpx5_core_146;
  wire popcount23_bpx5_core_147;
  wire popcount23_bpx5_core_148;
  wire popcount23_bpx5_core_151;
  wire popcount23_bpx5_core_153;
  wire popcount23_bpx5_core_155;
  wire popcount23_bpx5_core_156;
  wire popcount23_bpx5_core_159;
  wire popcount23_bpx5_core_160;
  wire popcount23_bpx5_core_161_not;
  wire popcount23_bpx5_core_166;
  wire popcount23_bpx5_core_167;

  assign popcount23_bpx5_core_026 = input_a[8] ^ input_a[7];
  assign popcount23_bpx5_core_027 = input_a[3] | input_a[2];
  assign popcount23_bpx5_core_028 = ~(input_a[14] ^ input_a[7]);
  assign popcount23_bpx5_core_029 = input_a[11] ^ input_a[0];
  assign popcount23_bpx5_core_030 = ~input_a[18];
  assign popcount23_bpx5_core_031 = ~(input_a[20] & input_a[3]);
  assign popcount23_bpx5_core_033 = input_a[13] ^ input_a[14];
  assign popcount23_bpx5_core_035 = ~(input_a[22] & input_a[10]);
  assign popcount23_bpx5_core_036 = ~input_a[4];
  assign popcount23_bpx5_core_038 = input_a[22] ^ input_a[11];
  assign popcount23_bpx5_core_040 = input_a[21] & input_a[5];
  assign popcount23_bpx5_core_042 = ~(input_a[3] ^ input_a[11]);
  assign popcount23_bpx5_core_043 = ~input_a[14];
  assign popcount23_bpx5_core_044_not = ~input_a[22];
  assign popcount23_bpx5_core_047 = input_a[13] & input_a[0];
  assign popcount23_bpx5_core_048 = ~(input_a[10] | input_a[15]);
  assign popcount23_bpx5_core_049 = input_a[16] | input_a[18];
  assign popcount23_bpx5_core_052 = input_a[7] ^ input_a[9];
  assign popcount23_bpx5_core_056 = input_a[6] ^ input_a[16];
  assign popcount23_bpx5_core_058 = input_a[1] & input_a[1];
  assign popcount23_bpx5_core_059 = input_a[20] ^ input_a[14];
  assign popcount23_bpx5_core_061 = input_a[22] & input_a[5];
  assign popcount23_bpx5_core_063 = ~input_a[6];
  assign popcount23_bpx5_core_065_not = ~input_a[0];
  assign popcount23_bpx5_core_066 = ~(input_a[4] | input_a[11]);
  assign popcount23_bpx5_core_067 = input_a[3] | input_a[15];
  assign popcount23_bpx5_core_069 = ~(input_a[7] & input_a[7]);
  assign popcount23_bpx5_core_070 = input_a[4] & input_a[17];
  assign popcount23_bpx5_core_071 = ~(input_a[0] & input_a[15]);
  assign popcount23_bpx5_core_072_not = ~input_a[0];
  assign popcount23_bpx5_core_073 = ~(input_a[16] & input_a[15]);
  assign popcount23_bpx5_core_074 = input_a[7] ^ input_a[19];
  assign popcount23_bpx5_core_075 = input_a[11] | input_a[21];
  assign popcount23_bpx5_core_076 = ~input_a[16];
  assign popcount23_bpx5_core_077 = input_a[12] ^ input_a[1];
  assign popcount23_bpx5_core_078 = ~(input_a[21] ^ input_a[18]);
  assign popcount23_bpx5_core_081 = input_a[21] ^ input_a[18];
  assign popcount23_bpx5_core_084 = ~(input_a[4] & input_a[22]);
  assign popcount23_bpx5_core_085 = input_a[20] & input_a[6];
  assign popcount23_bpx5_core_086 = input_a[8] ^ input_a[21];
  assign popcount23_bpx5_core_087 = input_a[12] & input_a[5];
  assign popcount23_bpx5_core_090 = ~(input_a[11] & input_a[22]);
  assign popcount23_bpx5_core_093_not = ~input_a[13];
  assign popcount23_bpx5_core_094 = ~(input_a[6] & input_a[14]);
  assign popcount23_bpx5_core_095 = ~input_a[17];
  assign popcount23_bpx5_core_096 = input_a[22] ^ input_a[5];
  assign popcount23_bpx5_core_097 = input_a[15] & input_a[11];
  assign popcount23_bpx5_core_098 = ~(input_a[12] | input_a[14]);
  assign popcount23_bpx5_core_100 = input_a[9] ^ input_a[13];
  assign popcount23_bpx5_core_101 = input_a[16] & input_a[12];
  assign popcount23_bpx5_core_102 = ~(input_a[13] ^ input_a[14]);
  assign popcount23_bpx5_core_104 = input_a[6] & input_a[15];
  assign popcount23_bpx5_core_107 = ~(input_a[10] ^ input_a[8]);
  assign popcount23_bpx5_core_110 = input_a[1] ^ input_a[15];
  assign popcount23_bpx5_core_111 = ~(input_a[16] ^ input_a[3]);
  assign popcount23_bpx5_core_112 = input_a[4] ^ input_a[5];
  assign popcount23_bpx5_core_114 = input_a[4] | input_a[8];
  assign popcount23_bpx5_core_120 = input_a[22] ^ input_a[2];
  assign popcount23_bpx5_core_122 = ~(input_a[18] & input_a[0]);
  assign popcount23_bpx5_core_123 = ~(input_a[10] & input_a[22]);
  assign popcount23_bpx5_core_125 = input_a[11] & input_a[18];
  assign popcount23_bpx5_core_126 = ~(input_a[18] | input_a[13]);
  assign popcount23_bpx5_core_127 = ~input_a[6];
  assign popcount23_bpx5_core_130 = ~input_a[16];
  assign popcount23_bpx5_core_131 = ~(input_a[0] ^ input_a[16]);
  assign popcount23_bpx5_core_133 = input_a[15] | input_a[1];
  assign popcount23_bpx5_core_134 = input_a[13] ^ input_a[2];
  assign popcount23_bpx5_core_135 = ~(input_a[0] & input_a[3]);
  assign popcount23_bpx5_core_136 = input_a[17] & input_a[13];
  assign popcount23_bpx5_core_138 = ~(input_a[12] | input_a[6]);
  assign popcount23_bpx5_core_139 = ~input_a[12];
  assign popcount23_bpx5_core_141 = input_a[5] ^ input_a[20];
  assign popcount23_bpx5_core_143 = ~input_a[22];
  assign popcount23_bpx5_core_145 = ~(input_a[13] & input_a[5]);
  assign popcount23_bpx5_core_146 = ~(input_a[10] & input_a[15]);
  assign popcount23_bpx5_core_147 = ~input_a[13];
  assign popcount23_bpx5_core_148 = ~input_a[16];
  assign popcount23_bpx5_core_151 = ~(input_a[1] | input_a[10]);
  assign popcount23_bpx5_core_153 = input_a[19] | input_a[17];
  assign popcount23_bpx5_core_155 = input_a[4] | input_a[5];
  assign popcount23_bpx5_core_156 = input_a[11] | input_a[8];
  assign popcount23_bpx5_core_159 = input_a[15] & input_a[2];
  assign popcount23_bpx5_core_160 = input_a[21] & input_a[5];
  assign popcount23_bpx5_core_161_not = ~input_a[14];
  assign popcount23_bpx5_core_166 = input_a[22] ^ input_a[9];
  assign popcount23_bpx5_core_167 = ~(input_a[4] & input_a[19]);

  assign popcount23_bpx5_out[0] = 1'b1;
  assign popcount23_bpx5_out[1] = input_a[16];
  assign popcount23_bpx5_out[2] = input_a[3];
  assign popcount23_bpx5_out[3] = 1'b1;
  assign popcount23_bpx5_out[4] = 1'b0;
endmodule