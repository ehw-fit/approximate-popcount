// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.9251
// WCE=24.0
// EP=0.892746%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount47_hhto(input [46:0] input_a, output [5:0] popcount47_hhto_out);
  wire popcount47_hhto_core_050;
  wire popcount47_hhto_core_051;
  wire popcount47_hhto_core_052;
  wire popcount47_hhto_core_053;
  wire popcount47_hhto_core_056;
  wire popcount47_hhto_core_058;
  wire popcount47_hhto_core_061;
  wire popcount47_hhto_core_062;
  wire popcount47_hhto_core_063;
  wire popcount47_hhto_core_064;
  wire popcount47_hhto_core_065;
  wire popcount47_hhto_core_066;
  wire popcount47_hhto_core_070;
  wire popcount47_hhto_core_071;
  wire popcount47_hhto_core_072;
  wire popcount47_hhto_core_074;
  wire popcount47_hhto_core_075;
  wire popcount47_hhto_core_076;
  wire popcount47_hhto_core_078;
  wire popcount47_hhto_core_079;
  wire popcount47_hhto_core_081;
  wire popcount47_hhto_core_083;
  wire popcount47_hhto_core_084;
  wire popcount47_hhto_core_085;
  wire popcount47_hhto_core_086;
  wire popcount47_hhto_core_088;
  wire popcount47_hhto_core_089;
  wire popcount47_hhto_core_090;
  wire popcount47_hhto_core_092;
  wire popcount47_hhto_core_094;
  wire popcount47_hhto_core_096;
  wire popcount47_hhto_core_097;
  wire popcount47_hhto_core_098;
  wire popcount47_hhto_core_099;
  wire popcount47_hhto_core_100;
  wire popcount47_hhto_core_101;
  wire popcount47_hhto_core_102;
  wire popcount47_hhto_core_103;
  wire popcount47_hhto_core_106;
  wire popcount47_hhto_core_107;
  wire popcount47_hhto_core_108;
  wire popcount47_hhto_core_112;
  wire popcount47_hhto_core_114;
  wire popcount47_hhto_core_115;
  wire popcount47_hhto_core_116;
  wire popcount47_hhto_core_119;
  wire popcount47_hhto_core_121;
  wire popcount47_hhto_core_123;
  wire popcount47_hhto_core_124;
  wire popcount47_hhto_core_125;
  wire popcount47_hhto_core_126;
  wire popcount47_hhto_core_127;
  wire popcount47_hhto_core_128;
  wire popcount47_hhto_core_131;
  wire popcount47_hhto_core_133;
  wire popcount47_hhto_core_134;
  wire popcount47_hhto_core_135;
  wire popcount47_hhto_core_136;
  wire popcount47_hhto_core_140;
  wire popcount47_hhto_core_142;
  wire popcount47_hhto_core_143;
  wire popcount47_hhto_core_144;
  wire popcount47_hhto_core_147;
  wire popcount47_hhto_core_149;
  wire popcount47_hhto_core_150;
  wire popcount47_hhto_core_152;
  wire popcount47_hhto_core_154;
  wire popcount47_hhto_core_156;
  wire popcount47_hhto_core_161;
  wire popcount47_hhto_core_162;
  wire popcount47_hhto_core_165;
  wire popcount47_hhto_core_166_not;
  wire popcount47_hhto_core_167;
  wire popcount47_hhto_core_168;
  wire popcount47_hhto_core_170;
  wire popcount47_hhto_core_172_not;
  wire popcount47_hhto_core_173;
  wire popcount47_hhto_core_174;
  wire popcount47_hhto_core_175;
  wire popcount47_hhto_core_176;
  wire popcount47_hhto_core_177;
  wire popcount47_hhto_core_182;
  wire popcount47_hhto_core_183;
  wire popcount47_hhto_core_184;
  wire popcount47_hhto_core_185;
  wire popcount47_hhto_core_187;
  wire popcount47_hhto_core_188;
  wire popcount47_hhto_core_189;
  wire popcount47_hhto_core_194;
  wire popcount47_hhto_core_195;
  wire popcount47_hhto_core_196;
  wire popcount47_hhto_core_198;
  wire popcount47_hhto_core_199;
  wire popcount47_hhto_core_200;
  wire popcount47_hhto_core_201;
  wire popcount47_hhto_core_202;
  wire popcount47_hhto_core_203;
  wire popcount47_hhto_core_205;
  wire popcount47_hhto_core_206;
  wire popcount47_hhto_core_208;
  wire popcount47_hhto_core_210;
  wire popcount47_hhto_core_216;
  wire popcount47_hhto_core_219;
  wire popcount47_hhto_core_220;
  wire popcount47_hhto_core_221;
  wire popcount47_hhto_core_222;
  wire popcount47_hhto_core_224;
  wire popcount47_hhto_core_226;
  wire popcount47_hhto_core_227;
  wire popcount47_hhto_core_228;
  wire popcount47_hhto_core_229;
  wire popcount47_hhto_core_231;
  wire popcount47_hhto_core_232;
  wire popcount47_hhto_core_233;
  wire popcount47_hhto_core_234;
  wire popcount47_hhto_core_235;
  wire popcount47_hhto_core_237;
  wire popcount47_hhto_core_239;
  wire popcount47_hhto_core_241;
  wire popcount47_hhto_core_243;
  wire popcount47_hhto_core_244;
  wire popcount47_hhto_core_245;
  wire popcount47_hhto_core_246;
  wire popcount47_hhto_core_247;
  wire popcount47_hhto_core_249;
  wire popcount47_hhto_core_250;
  wire popcount47_hhto_core_251;
  wire popcount47_hhto_core_252;
  wire popcount47_hhto_core_255;
  wire popcount47_hhto_core_256;
  wire popcount47_hhto_core_257;
  wire popcount47_hhto_core_258;
  wire popcount47_hhto_core_260;
  wire popcount47_hhto_core_261;
  wire popcount47_hhto_core_262_not;
  wire popcount47_hhto_core_263;
  wire popcount47_hhto_core_266;
  wire popcount47_hhto_core_268;
  wire popcount47_hhto_core_270;
  wire popcount47_hhto_core_272;
  wire popcount47_hhto_core_273;
  wire popcount47_hhto_core_274;
  wire popcount47_hhto_core_277;
  wire popcount47_hhto_core_278;
  wire popcount47_hhto_core_280;
  wire popcount47_hhto_core_281;
  wire popcount47_hhto_core_282;
  wire popcount47_hhto_core_283;
  wire popcount47_hhto_core_284;
  wire popcount47_hhto_core_285;
  wire popcount47_hhto_core_286;
  wire popcount47_hhto_core_287;
  wire popcount47_hhto_core_289;
  wire popcount47_hhto_core_291;
  wire popcount47_hhto_core_292;
  wire popcount47_hhto_core_294;
  wire popcount47_hhto_core_297;
  wire popcount47_hhto_core_299_not;
  wire popcount47_hhto_core_301;
  wire popcount47_hhto_core_302;
  wire popcount47_hhto_core_304;
  wire popcount47_hhto_core_305;
  wire popcount47_hhto_core_307;
  wire popcount47_hhto_core_309;
  wire popcount47_hhto_core_310;
  wire popcount47_hhto_core_311;
  wire popcount47_hhto_core_312;
  wire popcount47_hhto_core_313;
  wire popcount47_hhto_core_314;
  wire popcount47_hhto_core_316;
  wire popcount47_hhto_core_317_not;
  wire popcount47_hhto_core_320;
  wire popcount47_hhto_core_321;
  wire popcount47_hhto_core_322;
  wire popcount47_hhto_core_324_not;
  wire popcount47_hhto_core_326;
  wire popcount47_hhto_core_328;
  wire popcount47_hhto_core_330;
  wire popcount47_hhto_core_332;
  wire popcount47_hhto_core_336;
  wire popcount47_hhto_core_337;
  wire popcount47_hhto_core_338;
  wire popcount47_hhto_core_340;
  wire popcount47_hhto_core_342;
  wire popcount47_hhto_core_343;
  wire popcount47_hhto_core_345;
  wire popcount47_hhto_core_346;
  wire popcount47_hhto_core_347;
  wire popcount47_hhto_core_349;
  wire popcount47_hhto_core_350_not;
  wire popcount47_hhto_core_351;
  wire popcount47_hhto_core_352;
  wire popcount47_hhto_core_354;
  wire popcount47_hhto_core_356;
  wire popcount47_hhto_core_357;
  wire popcount47_hhto_core_361;
  wire popcount47_hhto_core_364;
  wire popcount47_hhto_core_370;
  wire popcount47_hhto_core_371;
  wire popcount47_hhto_core_372;

  assign popcount47_hhto_core_050 = input_a[5] ^ input_a[18];
  assign popcount47_hhto_core_051 = input_a[19] | input_a[40];
  assign popcount47_hhto_core_052 = ~(input_a[29] | input_a[43]);
  assign popcount47_hhto_core_053 = ~input_a[5];
  assign popcount47_hhto_core_056 = ~input_a[38];
  assign popcount47_hhto_core_058 = ~(input_a[34] ^ input_a[34]);
  assign popcount47_hhto_core_061 = input_a[3] | input_a[29];
  assign popcount47_hhto_core_062 = ~(input_a[26] | input_a[20]);
  assign popcount47_hhto_core_063 = input_a[16] | input_a[5];
  assign popcount47_hhto_core_064 = input_a[37] | input_a[31];
  assign popcount47_hhto_core_065 = ~(input_a[37] & input_a[1]);
  assign popcount47_hhto_core_066 = input_a[13] & input_a[33];
  assign popcount47_hhto_core_070 = ~input_a[45];
  assign popcount47_hhto_core_071 = ~(input_a[28] & input_a[39]);
  assign popcount47_hhto_core_072 = input_a[23] & input_a[34];
  assign popcount47_hhto_core_074 = input_a[4] ^ input_a[12];
  assign popcount47_hhto_core_075 = input_a[32] & input_a[34];
  assign popcount47_hhto_core_076 = input_a[46] ^ input_a[12];
  assign popcount47_hhto_core_078 = input_a[3] & input_a[12];
  assign popcount47_hhto_core_079 = ~(input_a[2] | input_a[5]);
  assign popcount47_hhto_core_081 = input_a[22] & input_a[43];
  assign popcount47_hhto_core_083 = input_a[26] | input_a[19];
  assign popcount47_hhto_core_084 = ~(input_a[33] ^ input_a[17]);
  assign popcount47_hhto_core_085 = ~(input_a[16] ^ input_a[7]);
  assign popcount47_hhto_core_086 = ~input_a[30];
  assign popcount47_hhto_core_088 = ~input_a[14];
  assign popcount47_hhto_core_089 = ~(input_a[22] & input_a[15]);
  assign popcount47_hhto_core_090 = ~(input_a[45] & input_a[17]);
  assign popcount47_hhto_core_092 = ~input_a[13];
  assign popcount47_hhto_core_094 = input_a[27] & input_a[23];
  assign popcount47_hhto_core_096 = input_a[45] ^ input_a[26];
  assign popcount47_hhto_core_097 = input_a[2] ^ input_a[44];
  assign popcount47_hhto_core_098 = input_a[42] & input_a[5];
  assign popcount47_hhto_core_099 = ~(input_a[40] ^ input_a[9]);
  assign popcount47_hhto_core_100 = ~(input_a[44] ^ input_a[19]);
  assign popcount47_hhto_core_101 = ~(input_a[32] | input_a[45]);
  assign popcount47_hhto_core_102 = ~(input_a[7] ^ input_a[46]);
  assign popcount47_hhto_core_103 = ~(input_a[12] ^ input_a[7]);
  assign popcount47_hhto_core_106 = ~(input_a[11] ^ input_a[20]);
  assign popcount47_hhto_core_107 = ~(input_a[19] & input_a[21]);
  assign popcount47_hhto_core_108 = input_a[8] | input_a[39];
  assign popcount47_hhto_core_112 = input_a[18] | input_a[6];
  assign popcount47_hhto_core_114 = ~input_a[17];
  assign popcount47_hhto_core_115 = input_a[29] & input_a[8];
  assign popcount47_hhto_core_116 = ~(input_a[0] ^ input_a[29]);
  assign popcount47_hhto_core_119 = input_a[36] & input_a[9];
  assign popcount47_hhto_core_121 = ~(input_a[29] & input_a[31]);
  assign popcount47_hhto_core_123 = input_a[2] ^ input_a[16];
  assign popcount47_hhto_core_124 = input_a[38] ^ input_a[30];
  assign popcount47_hhto_core_125 = ~(input_a[39] ^ input_a[20]);
  assign popcount47_hhto_core_126 = ~(input_a[18] & input_a[24]);
  assign popcount47_hhto_core_127 = input_a[30] & input_a[46];
  assign popcount47_hhto_core_128 = ~input_a[25];
  assign popcount47_hhto_core_131 = ~input_a[29];
  assign popcount47_hhto_core_133 = ~(input_a[12] & input_a[45]);
  assign popcount47_hhto_core_134 = ~(input_a[16] & input_a[36]);
  assign popcount47_hhto_core_135 = input_a[24] ^ input_a[45];
  assign popcount47_hhto_core_136 = ~input_a[32];
  assign popcount47_hhto_core_140 = ~input_a[26];
  assign popcount47_hhto_core_142 = ~(input_a[29] & input_a[39]);
  assign popcount47_hhto_core_143 = ~(input_a[31] & input_a[7]);
  assign popcount47_hhto_core_144 = input_a[9] | input_a[7];
  assign popcount47_hhto_core_147 = input_a[6] ^ input_a[5];
  assign popcount47_hhto_core_149 = input_a[11] & input_a[14];
  assign popcount47_hhto_core_150 = ~input_a[7];
  assign popcount47_hhto_core_152 = ~(input_a[34] ^ input_a[12]);
  assign popcount47_hhto_core_154 = ~(input_a[13] ^ input_a[20]);
  assign popcount47_hhto_core_156 = input_a[41] | input_a[18];
  assign popcount47_hhto_core_161 = input_a[44] | input_a[12];
  assign popcount47_hhto_core_162 = ~(input_a[14] & input_a[0]);
  assign popcount47_hhto_core_165 = ~(input_a[0] & input_a[26]);
  assign popcount47_hhto_core_166_not = ~input_a[16];
  assign popcount47_hhto_core_167 = input_a[4] ^ input_a[18];
  assign popcount47_hhto_core_168 = input_a[31] | input_a[44];
  assign popcount47_hhto_core_170 = input_a[22] & input_a[38];
  assign popcount47_hhto_core_172_not = ~input_a[45];
  assign popcount47_hhto_core_173 = input_a[18] & input_a[11];
  assign popcount47_hhto_core_174 = ~input_a[8];
  assign popcount47_hhto_core_175 = input_a[29] & input_a[28];
  assign popcount47_hhto_core_176 = ~input_a[20];
  assign popcount47_hhto_core_177 = input_a[41] & input_a[10];
  assign popcount47_hhto_core_182 = ~(input_a[24] | input_a[16]);
  assign popcount47_hhto_core_183 = input_a[27] ^ input_a[33];
  assign popcount47_hhto_core_184 = ~(input_a[46] ^ input_a[40]);
  assign popcount47_hhto_core_185 = ~input_a[2];
  assign popcount47_hhto_core_187 = input_a[31] & input_a[40];
  assign popcount47_hhto_core_188 = input_a[9] | input_a[16];
  assign popcount47_hhto_core_189 = ~(input_a[41] & input_a[32]);
  assign popcount47_hhto_core_194 = ~(input_a[26] ^ input_a[27]);
  assign popcount47_hhto_core_195 = input_a[0] & input_a[16];
  assign popcount47_hhto_core_196 = input_a[13] ^ input_a[21];
  assign popcount47_hhto_core_198 = ~(input_a[19] | input_a[16]);
  assign popcount47_hhto_core_199 = input_a[40] ^ input_a[2];
  assign popcount47_hhto_core_200 = ~(input_a[15] | input_a[5]);
  assign popcount47_hhto_core_201 = ~(input_a[38] & input_a[43]);
  assign popcount47_hhto_core_202 = input_a[35] | input_a[20];
  assign popcount47_hhto_core_203 = input_a[23] ^ input_a[9];
  assign popcount47_hhto_core_205 = ~input_a[25];
  assign popcount47_hhto_core_206 = ~(input_a[0] | input_a[14]);
  assign popcount47_hhto_core_208 = ~(input_a[44] & input_a[32]);
  assign popcount47_hhto_core_210 = input_a[2] ^ input_a[41];
  assign popcount47_hhto_core_216 = ~input_a[14];
  assign popcount47_hhto_core_219 = ~(input_a[14] & input_a[43]);
  assign popcount47_hhto_core_220 = ~(input_a[29] & input_a[29]);
  assign popcount47_hhto_core_221 = ~input_a[8];
  assign popcount47_hhto_core_222 = input_a[10] | input_a[30];
  assign popcount47_hhto_core_224 = input_a[5] & input_a[33];
  assign popcount47_hhto_core_226 = input_a[3] ^ input_a[5];
  assign popcount47_hhto_core_227 = ~(input_a[3] & input_a[14]);
  assign popcount47_hhto_core_228 = input_a[40] & input_a[29];
  assign popcount47_hhto_core_229 = ~(input_a[41] | input_a[32]);
  assign popcount47_hhto_core_231 = ~(input_a[6] | input_a[23]);
  assign popcount47_hhto_core_232 = ~(input_a[0] & input_a[29]);
  assign popcount47_hhto_core_233 = ~(input_a[17] ^ input_a[28]);
  assign popcount47_hhto_core_234 = ~(input_a[38] & input_a[2]);
  assign popcount47_hhto_core_235 = ~(input_a[0] | input_a[1]);
  assign popcount47_hhto_core_237 = ~(input_a[32] | input_a[5]);
  assign popcount47_hhto_core_239 = input_a[44] ^ input_a[9];
  assign popcount47_hhto_core_241 = ~(input_a[28] | input_a[35]);
  assign popcount47_hhto_core_243 = ~input_a[5];
  assign popcount47_hhto_core_244 = ~(input_a[16] | input_a[9]);
  assign popcount47_hhto_core_245 = ~(input_a[41] & input_a[28]);
  assign popcount47_hhto_core_246 = input_a[14] & input_a[8];
  assign popcount47_hhto_core_247 = ~(input_a[26] ^ input_a[20]);
  assign popcount47_hhto_core_249 = ~(input_a[39] & input_a[15]);
  assign popcount47_hhto_core_250 = input_a[26] | input_a[12];
  assign popcount47_hhto_core_251 = ~(input_a[17] & input_a[42]);
  assign popcount47_hhto_core_252 = input_a[35] & input_a[25];
  assign popcount47_hhto_core_255 = input_a[14] | input_a[28];
  assign popcount47_hhto_core_256 = input_a[23] ^ input_a[6];
  assign popcount47_hhto_core_257 = input_a[35] & input_a[13];
  assign popcount47_hhto_core_258 = input_a[42] | input_a[43];
  assign popcount47_hhto_core_260 = ~(input_a[36] | input_a[8]);
  assign popcount47_hhto_core_261 = ~(input_a[3] ^ input_a[0]);
  assign popcount47_hhto_core_262_not = ~input_a[24];
  assign popcount47_hhto_core_263 = ~(input_a[41] ^ input_a[25]);
  assign popcount47_hhto_core_266 = ~input_a[44];
  assign popcount47_hhto_core_268 = ~(input_a[21] | input_a[17]);
  assign popcount47_hhto_core_270 = ~(input_a[2] & input_a[16]);
  assign popcount47_hhto_core_272 = ~input_a[14];
  assign popcount47_hhto_core_273 = ~(input_a[46] & input_a[30]);
  assign popcount47_hhto_core_274 = ~(input_a[10] | input_a[30]);
  assign popcount47_hhto_core_277 = input_a[20] ^ input_a[35];
  assign popcount47_hhto_core_278 = ~(input_a[4] ^ input_a[8]);
  assign popcount47_hhto_core_280 = input_a[4] & input_a[40];
  assign popcount47_hhto_core_281 = ~(input_a[22] | input_a[6]);
  assign popcount47_hhto_core_282 = ~input_a[7];
  assign popcount47_hhto_core_283 = ~(input_a[32] ^ input_a[2]);
  assign popcount47_hhto_core_284 = input_a[10] & input_a[6];
  assign popcount47_hhto_core_285 = ~(input_a[30] & input_a[24]);
  assign popcount47_hhto_core_286 = ~(input_a[46] & input_a[10]);
  assign popcount47_hhto_core_287 = ~(input_a[8] & input_a[20]);
  assign popcount47_hhto_core_289 = ~(input_a[0] ^ input_a[16]);
  assign popcount47_hhto_core_291 = input_a[34] ^ input_a[10];
  assign popcount47_hhto_core_292 = ~(input_a[43] ^ input_a[10]);
  assign popcount47_hhto_core_294 = ~(input_a[10] & input_a[46]);
  assign popcount47_hhto_core_297 = ~(input_a[27] | input_a[14]);
  assign popcount47_hhto_core_299_not = ~input_a[39];
  assign popcount47_hhto_core_301 = ~input_a[35];
  assign popcount47_hhto_core_302 = input_a[17] & input_a[42];
  assign popcount47_hhto_core_304 = input_a[26] | input_a[44];
  assign popcount47_hhto_core_305 = ~(input_a[24] | input_a[35]);
  assign popcount47_hhto_core_307 = input_a[42] ^ input_a[38];
  assign popcount47_hhto_core_309 = input_a[18] & input_a[42];
  assign popcount47_hhto_core_310 = ~(input_a[43] | input_a[46]);
  assign popcount47_hhto_core_311 = input_a[37] | input_a[20];
  assign popcount47_hhto_core_312 = ~(input_a[8] | input_a[20]);
  assign popcount47_hhto_core_313 = input_a[21] | input_a[25];
  assign popcount47_hhto_core_314 = ~input_a[5];
  assign popcount47_hhto_core_316 = ~(input_a[45] | input_a[41]);
  assign popcount47_hhto_core_317_not = ~input_a[41];
  assign popcount47_hhto_core_320 = input_a[40] & input_a[12];
  assign popcount47_hhto_core_321 = ~(input_a[4] & input_a[40]);
  assign popcount47_hhto_core_322 = input_a[42] ^ input_a[2];
  assign popcount47_hhto_core_324_not = ~input_a[31];
  assign popcount47_hhto_core_326 = ~input_a[23];
  assign popcount47_hhto_core_328 = ~(input_a[15] & input_a[27]);
  assign popcount47_hhto_core_330 = ~(input_a[39] & input_a[39]);
  assign popcount47_hhto_core_332 = ~(input_a[19] | input_a[11]);
  assign popcount47_hhto_core_336 = ~(input_a[5] | input_a[8]);
  assign popcount47_hhto_core_337 = input_a[18] | input_a[13];
  assign popcount47_hhto_core_338 = input_a[37] | input_a[16];
  assign popcount47_hhto_core_340 = input_a[30] | input_a[20];
  assign popcount47_hhto_core_342 = ~(input_a[17] | input_a[23]);
  assign popcount47_hhto_core_343 = input_a[14] & input_a[44];
  assign popcount47_hhto_core_345 = ~(input_a[18] | input_a[16]);
  assign popcount47_hhto_core_346 = input_a[24] ^ input_a[37];
  assign popcount47_hhto_core_347 = ~(input_a[26] & input_a[34]);
  assign popcount47_hhto_core_349 = input_a[9] | input_a[37];
  assign popcount47_hhto_core_350_not = ~input_a[45];
  assign popcount47_hhto_core_351 = input_a[1] & input_a[35];
  assign popcount47_hhto_core_352 = ~(input_a[1] & input_a[42]);
  assign popcount47_hhto_core_354 = ~input_a[39];
  assign popcount47_hhto_core_356 = input_a[33] | input_a[27];
  assign popcount47_hhto_core_357 = ~(input_a[7] & input_a[40]);
  assign popcount47_hhto_core_361 = ~(input_a[4] ^ input_a[19]);
  assign popcount47_hhto_core_364 = input_a[41] & input_a[44];
  assign popcount47_hhto_core_370 = input_a[23] & input_a[25];
  assign popcount47_hhto_core_371 = input_a[11] ^ input_a[24];
  assign popcount47_hhto_core_372 = input_a[36] | input_a[1];

  assign popcount47_hhto_out[0] = input_a[25];
  assign popcount47_hhto_out[1] = input_a[12];
  assign popcount47_hhto_out[2] = popcount47_hhto_core_272;
  assign popcount47_hhto_out[3] = input_a[14];
  assign popcount47_hhto_out[4] = 1'b1;
  assign popcount47_hhto_out[5] = 1'b0;
endmodule