// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.75805
// WCE=15.0
// EP=0.931616%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount20_dajg(input [19:0] input_a, output [4:0] popcount20_dajg_out);
  wire popcount20_dajg_core_023;
  wire popcount20_dajg_core_024;
  wire popcount20_dajg_core_032;
  wire popcount20_dajg_core_033;
  wire popcount20_dajg_core_035;
  wire popcount20_dajg_core_036;
  wire popcount20_dajg_core_040;
  wire popcount20_dajg_core_041;
  wire popcount20_dajg_core_042;
  wire popcount20_dajg_core_044;
  wire popcount20_dajg_core_046;
  wire popcount20_dajg_core_047;
  wire popcount20_dajg_core_049;
  wire popcount20_dajg_core_051;
  wire popcount20_dajg_core_053;
  wire popcount20_dajg_core_054;
  wire popcount20_dajg_core_055;
  wire popcount20_dajg_core_058;
  wire popcount20_dajg_core_060;
  wire popcount20_dajg_core_062;
  wire popcount20_dajg_core_063_not;
  wire popcount20_dajg_core_064;
  wire popcount20_dajg_core_065;
  wire popcount20_dajg_core_066;
  wire popcount20_dajg_core_067;
  wire popcount20_dajg_core_068;
  wire popcount20_dajg_core_069;
  wire popcount20_dajg_core_070;
  wire popcount20_dajg_core_071_not;
  wire popcount20_dajg_core_072;
  wire popcount20_dajg_core_073;
  wire popcount20_dajg_core_074;
  wire popcount20_dajg_core_076;
  wire popcount20_dajg_core_078;
  wire popcount20_dajg_core_079;
  wire popcount20_dajg_core_081;
  wire popcount20_dajg_core_082;
  wire popcount20_dajg_core_083;
  wire popcount20_dajg_core_085;
  wire popcount20_dajg_core_087;
  wire popcount20_dajg_core_088;
  wire popcount20_dajg_core_089;
  wire popcount20_dajg_core_090;
  wire popcount20_dajg_core_093;
  wire popcount20_dajg_core_094;
  wire popcount20_dajg_core_095;
  wire popcount20_dajg_core_096;
  wire popcount20_dajg_core_097;
  wire popcount20_dajg_core_100;
  wire popcount20_dajg_core_103;
  wire popcount20_dajg_core_109;
  wire popcount20_dajg_core_111;
  wire popcount20_dajg_core_112;
  wire popcount20_dajg_core_114;
  wire popcount20_dajg_core_115_not;
  wire popcount20_dajg_core_116;
  wire popcount20_dajg_core_117;
  wire popcount20_dajg_core_118;
  wire popcount20_dajg_core_119;
  wire popcount20_dajg_core_120;
  wire popcount20_dajg_core_121;
  wire popcount20_dajg_core_122;
  wire popcount20_dajg_core_123;
  wire popcount20_dajg_core_125;
  wire popcount20_dajg_core_126;
  wire popcount20_dajg_core_127;
  wire popcount20_dajg_core_128;
  wire popcount20_dajg_core_131;
  wire popcount20_dajg_core_132;
  wire popcount20_dajg_core_133;
  wire popcount20_dajg_core_135;
  wire popcount20_dajg_core_136;
  wire popcount20_dajg_core_138;
  wire popcount20_dajg_core_140;
  wire popcount20_dajg_core_142;
  wire popcount20_dajg_core_144;

  assign popcount20_dajg_core_023 = input_a[15] | input_a[7];
  assign popcount20_dajg_core_024 = input_a[16] & input_a[1];
  assign popcount20_dajg_core_032 = ~(input_a[3] | input_a[15]);
  assign popcount20_dajg_core_033 = ~(input_a[8] | input_a[9]);
  assign popcount20_dajg_core_035 = ~(input_a[19] | input_a[18]);
  assign popcount20_dajg_core_036 = input_a[0] & input_a[5];
  assign popcount20_dajg_core_040 = ~input_a[12];
  assign popcount20_dajg_core_041 = ~(input_a[14] & input_a[0]);
  assign popcount20_dajg_core_042 = input_a[1] ^ input_a[9];
  assign popcount20_dajg_core_044 = input_a[16] ^ input_a[7];
  assign popcount20_dajg_core_046 = ~(input_a[3] & input_a[10]);
  assign popcount20_dajg_core_047 = ~(input_a[1] ^ input_a[9]);
  assign popcount20_dajg_core_049 = input_a[1] | input_a[6];
  assign popcount20_dajg_core_051 = ~(input_a[14] & input_a[13]);
  assign popcount20_dajg_core_053 = ~(input_a[14] ^ input_a[11]);
  assign popcount20_dajg_core_054 = input_a[14] & input_a[10];
  assign popcount20_dajg_core_055 = input_a[17] & input_a[16];
  assign popcount20_dajg_core_058 = ~input_a[10];
  assign popcount20_dajg_core_060 = input_a[16] & input_a[19];
  assign popcount20_dajg_core_062 = ~(input_a[13] & input_a[2]);
  assign popcount20_dajg_core_063_not = ~input_a[0];
  assign popcount20_dajg_core_064 = input_a[17] | input_a[1];
  assign popcount20_dajg_core_065 = ~(input_a[19] & input_a[7]);
  assign popcount20_dajg_core_066 = ~(input_a[8] | input_a[8]);
  assign popcount20_dajg_core_067 = ~(input_a[3] & input_a[16]);
  assign popcount20_dajg_core_068 = ~(input_a[14] & input_a[10]);
  assign popcount20_dajg_core_069 = input_a[7] | input_a[2];
  assign popcount20_dajg_core_070 = ~(input_a[8] ^ input_a[5]);
  assign popcount20_dajg_core_071_not = ~input_a[16];
  assign popcount20_dajg_core_072 = ~(input_a[6] | input_a[6]);
  assign popcount20_dajg_core_073 = ~(input_a[14] & input_a[3]);
  assign popcount20_dajg_core_074 = ~(input_a[9] ^ input_a[10]);
  assign popcount20_dajg_core_076 = ~(input_a[10] & input_a[16]);
  assign popcount20_dajg_core_078 = ~(input_a[11] | input_a[12]);
  assign popcount20_dajg_core_079 = ~(input_a[1] & input_a[19]);
  assign popcount20_dajg_core_081 = ~(input_a[7] ^ input_a[8]);
  assign popcount20_dajg_core_082 = input_a[2] | input_a[7];
  assign popcount20_dajg_core_083 = input_a[14] ^ input_a[2];
  assign popcount20_dajg_core_085 = ~(input_a[10] ^ input_a[15]);
  assign popcount20_dajg_core_087 = input_a[13] ^ input_a[11];
  assign popcount20_dajg_core_088 = input_a[16] ^ input_a[17];
  assign popcount20_dajg_core_089 = ~(input_a[8] | input_a[5]);
  assign popcount20_dajg_core_090 = input_a[10] | input_a[14];
  assign popcount20_dajg_core_093 = input_a[4] & input_a[18];
  assign popcount20_dajg_core_094 = ~(input_a[17] ^ input_a[10]);
  assign popcount20_dajg_core_095 = ~input_a[9];
  assign popcount20_dajg_core_096 = ~(input_a[10] | input_a[7]);
  assign popcount20_dajg_core_097 = input_a[18] ^ input_a[9];
  assign popcount20_dajg_core_100 = ~input_a[15];
  assign popcount20_dajg_core_103 = ~input_a[3];
  assign popcount20_dajg_core_109 = input_a[3] ^ input_a[5];
  assign popcount20_dajg_core_111 = ~(input_a[17] | input_a[10]);
  assign popcount20_dajg_core_112 = input_a[9] ^ input_a[17];
  assign popcount20_dajg_core_114 = input_a[1] & input_a[7];
  assign popcount20_dajg_core_115_not = ~input_a[3];
  assign popcount20_dajg_core_116 = ~(input_a[5] | input_a[14]);
  assign popcount20_dajg_core_117 = input_a[2] & input_a[4];
  assign popcount20_dajg_core_118 = ~(input_a[19] ^ input_a[15]);
  assign popcount20_dajg_core_119 = input_a[1] ^ input_a[7];
  assign popcount20_dajg_core_120 = ~(input_a[5] & input_a[10]);
  assign popcount20_dajg_core_121 = ~(input_a[16] ^ input_a[4]);
  assign popcount20_dajg_core_122 = ~(input_a[5] | input_a[17]);
  assign popcount20_dajg_core_123 = ~(input_a[4] | input_a[6]);
  assign popcount20_dajg_core_125 = ~(input_a[16] | input_a[5]);
  assign popcount20_dajg_core_126 = input_a[5] | input_a[17];
  assign popcount20_dajg_core_127 = ~(input_a[5] | input_a[2]);
  assign popcount20_dajg_core_128 = ~input_a[3];
  assign popcount20_dajg_core_131 = ~(input_a[16] ^ input_a[9]);
  assign popcount20_dajg_core_132 = input_a[2] | input_a[8];
  assign popcount20_dajg_core_133 = input_a[11] ^ input_a[0];
  assign popcount20_dajg_core_135 = input_a[6] ^ input_a[14];
  assign popcount20_dajg_core_136 = input_a[7] ^ input_a[4];
  assign popcount20_dajg_core_138 = ~(input_a[19] & input_a[2]);
  assign popcount20_dajg_core_140 = ~(input_a[15] & input_a[3]);
  assign popcount20_dajg_core_142 = ~(input_a[10] | input_a[6]);
  assign popcount20_dajg_core_144 = input_a[8] ^ input_a[10];

  assign popcount20_dajg_out[0] = 1'b1;
  assign popcount20_dajg_out[1] = 1'b1;
  assign popcount20_dajg_out[2] = input_a[19];
  assign popcount20_dajg_out[3] = input_a[0];
  assign popcount20_dajg_out[4] = 1'b0;
endmodule