// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.63899
// WCE=12.0
// EP=0.808142%
// Printed PDK parameters:
//  Area=44775968.0
//  Delay=67857376.0
//  Power=2030100.0

module popcount33_5ac0(input [32:0] input_a, output [5:0] popcount33_5ac0_out);
  wire popcount33_5ac0_core_035;
  wire popcount33_5ac0_core_036;
  wire popcount33_5ac0_core_037;
  wire popcount33_5ac0_core_038;
  wire popcount33_5ac0_core_039;
  wire popcount33_5ac0_core_040;
  wire popcount33_5ac0_core_041;
  wire popcount33_5ac0_core_042;
  wire popcount33_5ac0_core_043;
  wire popcount33_5ac0_core_047;
  wire popcount33_5ac0_core_048;
  wire popcount33_5ac0_core_051;
  wire popcount33_5ac0_core_052;
  wire popcount33_5ac0_core_054;
  wire popcount33_5ac0_core_055;
  wire popcount33_5ac0_core_056;
  wire popcount33_5ac0_core_058;
  wire popcount33_5ac0_core_059;
  wire popcount33_5ac0_core_060;
  wire popcount33_5ac0_core_061;
  wire popcount33_5ac0_core_062;
  wire popcount33_5ac0_core_063;
  wire popcount33_5ac0_core_068;
  wire popcount33_5ac0_core_070;
  wire popcount33_5ac0_core_071;
  wire popcount33_5ac0_core_072;
  wire popcount33_5ac0_core_073;
  wire popcount33_5ac0_core_074;
  wire popcount33_5ac0_core_075;
  wire popcount33_5ac0_core_076;
  wire popcount33_5ac0_core_080;
  wire popcount33_5ac0_core_081;
  wire popcount33_5ac0_core_083;
  wire popcount33_5ac0_core_084;
  wire popcount33_5ac0_core_085;
  wire popcount33_5ac0_core_086;
  wire popcount33_5ac0_core_087;
  wire popcount33_5ac0_core_088;
  wire popcount33_5ac0_core_090;
  wire popcount33_5ac0_core_092;
  wire popcount33_5ac0_core_093;
  wire popcount33_5ac0_core_096;
  wire popcount33_5ac0_core_103;
  wire popcount33_5ac0_core_104;
  wire popcount33_5ac0_core_105;
  wire popcount33_5ac0_core_106;
  wire popcount33_5ac0_core_110;
  wire popcount33_5ac0_core_111;
  wire popcount33_5ac0_core_112;
  wire popcount33_5ac0_core_113;
  wire popcount33_5ac0_core_114;
  wire popcount33_5ac0_core_116;
  wire popcount33_5ac0_core_118;
  wire popcount33_5ac0_core_121;
  wire popcount33_5ac0_core_122;
  wire popcount33_5ac0_core_123;
  wire popcount33_5ac0_core_124;
  wire popcount33_5ac0_core_127;
  wire popcount33_5ac0_core_128;
  wire popcount33_5ac0_core_129;
  wire popcount33_5ac0_core_130;
  wire popcount33_5ac0_core_131;
  wire popcount33_5ac0_core_132;
  wire popcount33_5ac0_core_134;
  wire popcount33_5ac0_core_136;
  wire popcount33_5ac0_core_137;
  wire popcount33_5ac0_core_138;
  wire popcount33_5ac0_core_139;
  wire popcount33_5ac0_core_141;
  wire popcount33_5ac0_core_143;
  wire popcount33_5ac0_core_144;
  wire popcount33_5ac0_core_145;
  wire popcount33_5ac0_core_146;
  wire popcount33_5ac0_core_147;
  wire popcount33_5ac0_core_148;
  wire popcount33_5ac0_core_152;
  wire popcount33_5ac0_core_155;
  wire popcount33_5ac0_core_156_not;
  wire popcount33_5ac0_core_157;
  wire popcount33_5ac0_core_158;
  wire popcount33_5ac0_core_159;
  wire popcount33_5ac0_core_160;
  wire popcount33_5ac0_core_161;
  wire popcount33_5ac0_core_162;
  wire popcount33_5ac0_core_163;
  wire popcount33_5ac0_core_164;
  wire popcount33_5ac0_core_167;
  wire popcount33_5ac0_core_168;
  wire popcount33_5ac0_core_169;
  wire popcount33_5ac0_core_171;
  wire popcount33_5ac0_core_172;
  wire popcount33_5ac0_core_173;
  wire popcount33_5ac0_core_175;
  wire popcount33_5ac0_core_176;
  wire popcount33_5ac0_core_180;
  wire popcount33_5ac0_core_182;
  wire popcount33_5ac0_core_184;
  wire popcount33_5ac0_core_185;
  wire popcount33_5ac0_core_187;
  wire popcount33_5ac0_core_189;
  wire popcount33_5ac0_core_190;
  wire popcount33_5ac0_core_191;
  wire popcount33_5ac0_core_192;
  wire popcount33_5ac0_core_193;
  wire popcount33_5ac0_core_196;
  wire popcount33_5ac0_core_197;
  wire popcount33_5ac0_core_198;
  wire popcount33_5ac0_core_199;
  wire popcount33_5ac0_core_200;
  wire popcount33_5ac0_core_201;
  wire popcount33_5ac0_core_202;
  wire popcount33_5ac0_core_203;
  wire popcount33_5ac0_core_204;
  wire popcount33_5ac0_core_205;
  wire popcount33_5ac0_core_206;
  wire popcount33_5ac0_core_207;
  wire popcount33_5ac0_core_210;
  wire popcount33_5ac0_core_211;
  wire popcount33_5ac0_core_215;
  wire popcount33_5ac0_core_217;
  wire popcount33_5ac0_core_218;
  wire popcount33_5ac0_core_219;
  wire popcount33_5ac0_core_220;
  wire popcount33_5ac0_core_222;
  wire popcount33_5ac0_core_223;
  wire popcount33_5ac0_core_224;
  wire popcount33_5ac0_core_225;
  wire popcount33_5ac0_core_226;
  wire popcount33_5ac0_core_227;
  wire popcount33_5ac0_core_228;
  wire popcount33_5ac0_core_229;
  wire popcount33_5ac0_core_230;
  wire popcount33_5ac0_core_231;
  wire popcount33_5ac0_core_233;
  wire popcount33_5ac0_core_234;
  wire popcount33_5ac0_core_235;
  wire popcount33_5ac0_core_236;
  wire popcount33_5ac0_core_237;

  assign popcount33_5ac0_core_035 = input_a[3] | input_a[17];
  assign popcount33_5ac0_core_036 = input_a[18] | input_a[5];
  assign popcount33_5ac0_core_037 = input_a[13] | input_a[14];
  assign popcount33_5ac0_core_038 = input_a[28] ^ input_a[10];
  assign popcount33_5ac0_core_039 = ~(input_a[23] | input_a[4]);
  assign popcount33_5ac0_core_040 = popcount33_5ac0_core_035 & popcount33_5ac0_core_037;
  assign popcount33_5ac0_core_041 = ~(input_a[9] | input_a[29]);
  assign popcount33_5ac0_core_042 = ~input_a[23];
  assign popcount33_5ac0_core_043 = input_a[24] | popcount33_5ac0_core_040;
  assign popcount33_5ac0_core_047 = ~input_a[18];
  assign popcount33_5ac0_core_048 = ~(input_a[17] & input_a[16]);
  assign popcount33_5ac0_core_051 = ~input_a[11];
  assign popcount33_5ac0_core_052 = ~(input_a[20] | input_a[31]);
  assign popcount33_5ac0_core_054 = input_a[29] | input_a[22];
  assign popcount33_5ac0_core_055 = input_a[2] | input_a[31];
  assign popcount33_5ac0_core_056 = ~input_a[12];
  assign popcount33_5ac0_core_058 = input_a[4] & input_a[31];
  assign popcount33_5ac0_core_059 = popcount33_5ac0_core_043 ^ popcount33_5ac0_core_054;
  assign popcount33_5ac0_core_060 = popcount33_5ac0_core_043 & popcount33_5ac0_core_054;
  assign popcount33_5ac0_core_061 = popcount33_5ac0_core_059 ^ popcount33_5ac0_core_058;
  assign popcount33_5ac0_core_062 = popcount33_5ac0_core_059 & popcount33_5ac0_core_058;
  assign popcount33_5ac0_core_063 = popcount33_5ac0_core_060 | popcount33_5ac0_core_062;
  assign popcount33_5ac0_core_068 = ~(input_a[7] ^ input_a[17]);
  assign popcount33_5ac0_core_070 = input_a[0] & input_a[27];
  assign popcount33_5ac0_core_071 = ~(input_a[10] ^ input_a[6]);
  assign popcount33_5ac0_core_072 = input_a[1] & input_a[7];
  assign popcount33_5ac0_core_073 = ~(input_a[31] ^ input_a[26]);
  assign popcount33_5ac0_core_074 = ~(input_a[22] | input_a[5]);
  assign popcount33_5ac0_core_075 = popcount33_5ac0_core_070 | popcount33_5ac0_core_072;
  assign popcount33_5ac0_core_076 = input_a[18] | input_a[24];
  assign popcount33_5ac0_core_080 = ~(input_a[29] & input_a[0]);
  assign popcount33_5ac0_core_081 = input_a[29] & input_a[23];
  assign popcount33_5ac0_core_083 = input_a[0] ^ input_a[26];
  assign popcount33_5ac0_core_084 = ~input_a[4];
  assign popcount33_5ac0_core_085 = input_a[8] | input_a[14];
  assign popcount33_5ac0_core_086 = ~input_a[29];
  assign popcount33_5ac0_core_087 = ~(input_a[13] | input_a[26]);
  assign popcount33_5ac0_core_088 = ~(input_a[20] ^ input_a[15]);
  assign popcount33_5ac0_core_090 = ~(input_a[24] & input_a[27]);
  assign popcount33_5ac0_core_092 = ~(input_a[32] | input_a[14]);
  assign popcount33_5ac0_core_093 = ~popcount33_5ac0_core_075;
  assign popcount33_5ac0_core_096 = ~(input_a[4] & input_a[3]);
  assign popcount33_5ac0_core_103 = ~(input_a[22] | input_a[15]);
  assign popcount33_5ac0_core_104 = ~(input_a[14] & input_a[0]);
  assign popcount33_5ac0_core_105 = popcount33_5ac0_core_061 ^ popcount33_5ac0_core_093;
  assign popcount33_5ac0_core_106 = popcount33_5ac0_core_061 & popcount33_5ac0_core_093;
  assign popcount33_5ac0_core_110 = popcount33_5ac0_core_063 ^ popcount33_5ac0_core_075;
  assign popcount33_5ac0_core_111 = popcount33_5ac0_core_063 & popcount33_5ac0_core_075;
  assign popcount33_5ac0_core_112 = popcount33_5ac0_core_110 ^ popcount33_5ac0_core_106;
  assign popcount33_5ac0_core_113 = popcount33_5ac0_core_110 & popcount33_5ac0_core_106;
  assign popcount33_5ac0_core_114 = popcount33_5ac0_core_111 | popcount33_5ac0_core_113;
  assign popcount33_5ac0_core_116 = ~(input_a[9] ^ input_a[19]);
  assign popcount33_5ac0_core_118 = ~(input_a[4] ^ input_a[12]);
  assign popcount33_5ac0_core_121 = ~(input_a[4] | input_a[22]);
  assign popcount33_5ac0_core_122 = input_a[5] ^ input_a[8];
  assign popcount33_5ac0_core_123 = ~input_a[12];
  assign popcount33_5ac0_core_124 = ~(input_a[11] ^ input_a[14]);
  assign popcount33_5ac0_core_127 = ~(input_a[20] ^ input_a[16]);
  assign popcount33_5ac0_core_128 = input_a[18] | input_a[6];
  assign popcount33_5ac0_core_129 = ~input_a[25];
  assign popcount33_5ac0_core_130 = input_a[31] | input_a[4];
  assign popcount33_5ac0_core_131 = input_a[15] | input_a[4];
  assign popcount33_5ac0_core_132 = input_a[20] & input_a[5];
  assign popcount33_5ac0_core_134 = input_a[23] & input_a[9];
  assign popcount33_5ac0_core_136 = input_a[15] & input_a[11];
  assign popcount33_5ac0_core_137 = popcount33_5ac0_core_132 | popcount33_5ac0_core_134;
  assign popcount33_5ac0_core_138 = ~(input_a[21] & input_a[29]);
  assign popcount33_5ac0_core_139 = popcount33_5ac0_core_137 | popcount33_5ac0_core_136;
  assign popcount33_5ac0_core_141 = input_a[9] & input_a[24];
  assign popcount33_5ac0_core_143 = input_a[21] & input_a[25];
  assign popcount33_5ac0_core_144 = popcount33_5ac0_core_128 ^ popcount33_5ac0_core_139;
  assign popcount33_5ac0_core_145 = popcount33_5ac0_core_128 & popcount33_5ac0_core_139;
  assign popcount33_5ac0_core_146 = popcount33_5ac0_core_144 ^ popcount33_5ac0_core_143;
  assign popcount33_5ac0_core_147 = popcount33_5ac0_core_144 & popcount33_5ac0_core_143;
  assign popcount33_5ac0_core_148 = popcount33_5ac0_core_145 | popcount33_5ac0_core_147;
  assign popcount33_5ac0_core_152 = input_a[6] | input_a[13];
  assign popcount33_5ac0_core_155 = input_a[10] & input_a[8];
  assign popcount33_5ac0_core_156_not = ~input_a[22];
  assign popcount33_5ac0_core_157 = input_a[2] & input_a[26];
  assign popcount33_5ac0_core_158 = ~(input_a[10] | input_a[21]);
  assign popcount33_5ac0_core_159 = input_a[28] & input_a[16];
  assign popcount33_5ac0_core_160 = popcount33_5ac0_core_155 ^ popcount33_5ac0_core_157;
  assign popcount33_5ac0_core_161 = popcount33_5ac0_core_155 & popcount33_5ac0_core_157;
  assign popcount33_5ac0_core_162 = popcount33_5ac0_core_160 ^ popcount33_5ac0_core_159;
  assign popcount33_5ac0_core_163 = popcount33_5ac0_core_160 & popcount33_5ac0_core_159;
  assign popcount33_5ac0_core_164 = popcount33_5ac0_core_161 | popcount33_5ac0_core_163;
  assign popcount33_5ac0_core_167 = ~(input_a[23] | input_a[5]);
  assign popcount33_5ac0_core_168 = ~input_a[13];
  assign popcount33_5ac0_core_169 = ~(input_a[4] & input_a[24]);
  assign popcount33_5ac0_core_171 = ~(input_a[12] & input_a[30]);
  assign popcount33_5ac0_core_172 = input_a[12] & input_a[30];
  assign popcount33_5ac0_core_173 = input_a[16] ^ input_a[18];
  assign popcount33_5ac0_core_175 = input_a[19] ^ popcount33_5ac0_core_171;
  assign popcount33_5ac0_core_176 = input_a[25] | input_a[17];
  assign popcount33_5ac0_core_180 = popcount33_5ac0_core_172 | input_a[19];
  assign popcount33_5ac0_core_182 = ~(input_a[0] & input_a[24]);
  assign popcount33_5ac0_core_184 = popcount33_5ac0_core_162 ^ popcount33_5ac0_core_175;
  assign popcount33_5ac0_core_185 = popcount33_5ac0_core_162 & popcount33_5ac0_core_175;
  assign popcount33_5ac0_core_187 = input_a[30] & input_a[25];
  assign popcount33_5ac0_core_189 = popcount33_5ac0_core_164 ^ popcount33_5ac0_core_180;
  assign popcount33_5ac0_core_190 = popcount33_5ac0_core_164 & popcount33_5ac0_core_180;
  assign popcount33_5ac0_core_191 = popcount33_5ac0_core_189 ^ popcount33_5ac0_core_185;
  assign popcount33_5ac0_core_192 = popcount33_5ac0_core_189 & popcount33_5ac0_core_185;
  assign popcount33_5ac0_core_193 = popcount33_5ac0_core_190 | popcount33_5ac0_core_192;
  assign popcount33_5ac0_core_196 = ~(input_a[13] ^ input_a[18]);
  assign popcount33_5ac0_core_197 = input_a[10] ^ input_a[28];
  assign popcount33_5ac0_core_198 = popcount33_5ac0_core_146 ^ popcount33_5ac0_core_184;
  assign popcount33_5ac0_core_199 = popcount33_5ac0_core_146 & popcount33_5ac0_core_184;
  assign popcount33_5ac0_core_200 = ~(popcount33_5ac0_core_198 & input_a[32]);
  assign popcount33_5ac0_core_201 = popcount33_5ac0_core_198 & input_a[32];
  assign popcount33_5ac0_core_202 = popcount33_5ac0_core_199 | popcount33_5ac0_core_201;
  assign popcount33_5ac0_core_203 = popcount33_5ac0_core_148 ^ popcount33_5ac0_core_191;
  assign popcount33_5ac0_core_204 = popcount33_5ac0_core_148 & popcount33_5ac0_core_191;
  assign popcount33_5ac0_core_205 = popcount33_5ac0_core_203 ^ popcount33_5ac0_core_202;
  assign popcount33_5ac0_core_206 = popcount33_5ac0_core_203 & popcount33_5ac0_core_202;
  assign popcount33_5ac0_core_207 = popcount33_5ac0_core_204 | popcount33_5ac0_core_206;
  assign popcount33_5ac0_core_210 = popcount33_5ac0_core_193 ^ popcount33_5ac0_core_207;
  assign popcount33_5ac0_core_211 = popcount33_5ac0_core_193 & popcount33_5ac0_core_207;
  assign popcount33_5ac0_core_215 = input_a[6] & input_a[5];
  assign popcount33_5ac0_core_217 = ~(popcount33_5ac0_core_105 & popcount33_5ac0_core_200);
  assign popcount33_5ac0_core_218 = popcount33_5ac0_core_105 & popcount33_5ac0_core_200;
  assign popcount33_5ac0_core_219 = input_a[3] | input_a[19];
  assign popcount33_5ac0_core_220 = ~(input_a[21] | input_a[28]);
  assign popcount33_5ac0_core_222 = popcount33_5ac0_core_112 ^ popcount33_5ac0_core_205;
  assign popcount33_5ac0_core_223 = popcount33_5ac0_core_112 & popcount33_5ac0_core_205;
  assign popcount33_5ac0_core_224 = popcount33_5ac0_core_222 ^ popcount33_5ac0_core_218;
  assign popcount33_5ac0_core_225 = popcount33_5ac0_core_222 & popcount33_5ac0_core_218;
  assign popcount33_5ac0_core_226 = popcount33_5ac0_core_223 | popcount33_5ac0_core_225;
  assign popcount33_5ac0_core_227 = popcount33_5ac0_core_114 ^ popcount33_5ac0_core_210;
  assign popcount33_5ac0_core_228 = popcount33_5ac0_core_114 & popcount33_5ac0_core_210;
  assign popcount33_5ac0_core_229 = popcount33_5ac0_core_227 ^ popcount33_5ac0_core_226;
  assign popcount33_5ac0_core_230 = popcount33_5ac0_core_227 & popcount33_5ac0_core_226;
  assign popcount33_5ac0_core_231 = popcount33_5ac0_core_228 | popcount33_5ac0_core_230;
  assign popcount33_5ac0_core_233 = input_a[23] ^ input_a[8];
  assign popcount33_5ac0_core_234 = popcount33_5ac0_core_211 | popcount33_5ac0_core_231;
  assign popcount33_5ac0_core_235 = input_a[5] ^ input_a[10];
  assign popcount33_5ac0_core_236 = ~(input_a[6] & input_a[19]);
  assign popcount33_5ac0_core_237 = ~input_a[1];

  assign popcount33_5ac0_out[0] = popcount33_5ac0_core_217;
  assign popcount33_5ac0_out[1] = popcount33_5ac0_core_229;
  assign popcount33_5ac0_out[2] = popcount33_5ac0_core_224;
  assign popcount33_5ac0_out[3] = popcount33_5ac0_core_229;
  assign popcount33_5ac0_out[4] = popcount33_5ac0_core_234;
  assign popcount33_5ac0_out[5] = 1'b0;
endmodule