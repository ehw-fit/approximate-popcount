// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.66364
// WCE=26.0
// EP=0.943107%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_hnxw(input [33:0] input_a, output [5:0] popcount34_hnxw_out);
  wire popcount34_hnxw_core_037;
  wire popcount34_hnxw_core_038;
  wire popcount34_hnxw_core_040;
  wire popcount34_hnxw_core_041;
  wire popcount34_hnxw_core_042;
  wire popcount34_hnxw_core_043;
  wire popcount34_hnxw_core_044;
  wire popcount34_hnxw_core_048;
  wire popcount34_hnxw_core_049;
  wire popcount34_hnxw_core_050;
  wire popcount34_hnxw_core_052;
  wire popcount34_hnxw_core_053;
  wire popcount34_hnxw_core_054;
  wire popcount34_hnxw_core_056;
  wire popcount34_hnxw_core_057;
  wire popcount34_hnxw_core_059;
  wire popcount34_hnxw_core_060;
  wire popcount34_hnxw_core_061;
  wire popcount34_hnxw_core_062;
  wire popcount34_hnxw_core_063;
  wire popcount34_hnxw_core_064;
  wire popcount34_hnxw_core_065;
  wire popcount34_hnxw_core_066;
  wire popcount34_hnxw_core_067;
  wire popcount34_hnxw_core_068;
  wire popcount34_hnxw_core_069;
  wire popcount34_hnxw_core_070;
  wire popcount34_hnxw_core_072;
  wire popcount34_hnxw_core_073;
  wire popcount34_hnxw_core_076;
  wire popcount34_hnxw_core_079;
  wire popcount34_hnxw_core_080;
  wire popcount34_hnxw_core_082;
  wire popcount34_hnxw_core_083;
  wire popcount34_hnxw_core_084;
  wire popcount34_hnxw_core_086_not;
  wire popcount34_hnxw_core_087;
  wire popcount34_hnxw_core_088_not;
  wire popcount34_hnxw_core_089;
  wire popcount34_hnxw_core_090;
  wire popcount34_hnxw_core_092;
  wire popcount34_hnxw_core_093;
  wire popcount34_hnxw_core_094;
  wire popcount34_hnxw_core_095;
  wire popcount34_hnxw_core_097;
  wire popcount34_hnxw_core_098;
  wire popcount34_hnxw_core_099;
  wire popcount34_hnxw_core_100;
  wire popcount34_hnxw_core_101;
  wire popcount34_hnxw_core_102;
  wire popcount34_hnxw_core_105;
  wire popcount34_hnxw_core_107;
  wire popcount34_hnxw_core_109;
  wire popcount34_hnxw_core_113;
  wire popcount34_hnxw_core_114;
  wire popcount34_hnxw_core_116;
  wire popcount34_hnxw_core_117;
  wire popcount34_hnxw_core_118;
  wire popcount34_hnxw_core_119;
  wire popcount34_hnxw_core_121;
  wire popcount34_hnxw_core_124;
  wire popcount34_hnxw_core_125;
  wire popcount34_hnxw_core_126;
  wire popcount34_hnxw_core_128;
  wire popcount34_hnxw_core_130;
  wire popcount34_hnxw_core_131;
  wire popcount34_hnxw_core_134;
  wire popcount34_hnxw_core_136;
  wire popcount34_hnxw_core_137;
  wire popcount34_hnxw_core_138;
  wire popcount34_hnxw_core_139;
  wire popcount34_hnxw_core_142;
  wire popcount34_hnxw_core_144;
  wire popcount34_hnxw_core_145;
  wire popcount34_hnxw_core_149;
  wire popcount34_hnxw_core_150;
  wire popcount34_hnxw_core_153;
  wire popcount34_hnxw_core_156;
  wire popcount34_hnxw_core_157;
  wire popcount34_hnxw_core_158;
  wire popcount34_hnxw_core_159;
  wire popcount34_hnxw_core_160;
  wire popcount34_hnxw_core_164;
  wire popcount34_hnxw_core_167;
  wire popcount34_hnxw_core_169_not;
  wire popcount34_hnxw_core_170;
  wire popcount34_hnxw_core_171;
  wire popcount34_hnxw_core_172;
  wire popcount34_hnxw_core_173;
  wire popcount34_hnxw_core_175;
  wire popcount34_hnxw_core_176;
  wire popcount34_hnxw_core_177;
  wire popcount34_hnxw_core_178;
  wire popcount34_hnxw_core_179;
  wire popcount34_hnxw_core_180;
  wire popcount34_hnxw_core_181;
  wire popcount34_hnxw_core_183;
  wire popcount34_hnxw_core_184;
  wire popcount34_hnxw_core_185;
  wire popcount34_hnxw_core_188;
  wire popcount34_hnxw_core_189;
  wire popcount34_hnxw_core_190;
  wire popcount34_hnxw_core_191;
  wire popcount34_hnxw_core_192;
  wire popcount34_hnxw_core_193;
  wire popcount34_hnxw_core_194;
  wire popcount34_hnxw_core_196;
  wire popcount34_hnxw_core_197;
  wire popcount34_hnxw_core_202;
  wire popcount34_hnxw_core_203;
  wire popcount34_hnxw_core_204_not;
  wire popcount34_hnxw_core_205;
  wire popcount34_hnxw_core_207;
  wire popcount34_hnxw_core_208;
  wire popcount34_hnxw_core_209;
  wire popcount34_hnxw_core_212;
  wire popcount34_hnxw_core_213;
  wire popcount34_hnxw_core_214;
  wire popcount34_hnxw_core_216;
  wire popcount34_hnxw_core_217;
  wire popcount34_hnxw_core_219;
  wire popcount34_hnxw_core_221;
  wire popcount34_hnxw_core_222;
  wire popcount34_hnxw_core_224;
  wire popcount34_hnxw_core_225;
  wire popcount34_hnxw_core_226;
  wire popcount34_hnxw_core_228;
  wire popcount34_hnxw_core_229;
  wire popcount34_hnxw_core_230;
  wire popcount34_hnxw_core_231;
  wire popcount34_hnxw_core_232;
  wire popcount34_hnxw_core_234;
  wire popcount34_hnxw_core_237;
  wire popcount34_hnxw_core_238;
  wire popcount34_hnxw_core_239;
  wire popcount34_hnxw_core_244;
  wire popcount34_hnxw_core_246;
  wire popcount34_hnxw_core_247;
  wire popcount34_hnxw_core_248;
  wire popcount34_hnxw_core_249;
  wire popcount34_hnxw_core_250;

  assign popcount34_hnxw_core_037 = ~input_a[1];
  assign popcount34_hnxw_core_038 = input_a[11] | input_a[26];
  assign popcount34_hnxw_core_040 = ~(input_a[1] | input_a[9]);
  assign popcount34_hnxw_core_041 = input_a[8] | input_a[29];
  assign popcount34_hnxw_core_042 = ~(input_a[25] | input_a[5]);
  assign popcount34_hnxw_core_043 = input_a[23] ^ input_a[6];
  assign popcount34_hnxw_core_044 = input_a[4] ^ input_a[20];
  assign popcount34_hnxw_core_048 = ~input_a[1];
  assign popcount34_hnxw_core_049 = ~input_a[31];
  assign popcount34_hnxw_core_050 = ~(input_a[8] | input_a[13]);
  assign popcount34_hnxw_core_052 = ~input_a[27];
  assign popcount34_hnxw_core_053 = input_a[25] & input_a[28];
  assign popcount34_hnxw_core_054 = input_a[28] & input_a[10];
  assign popcount34_hnxw_core_056 = ~(input_a[27] | input_a[18]);
  assign popcount34_hnxw_core_057 = ~(input_a[20] & input_a[9]);
  assign popcount34_hnxw_core_059 = ~input_a[33];
  assign popcount34_hnxw_core_060 = ~(input_a[19] | input_a[30]);
  assign popcount34_hnxw_core_061 = ~input_a[3];
  assign popcount34_hnxw_core_062 = input_a[25] & input_a[32];
  assign popcount34_hnxw_core_063 = ~(input_a[28] ^ input_a[17]);
  assign popcount34_hnxw_core_064 = input_a[7] ^ input_a[16];
  assign popcount34_hnxw_core_065 = input_a[26] | input_a[30];
  assign popcount34_hnxw_core_066 = ~(input_a[22] | input_a[28]);
  assign popcount34_hnxw_core_067 = input_a[9] ^ input_a[2];
  assign popcount34_hnxw_core_068 = input_a[32] ^ input_a[6];
  assign popcount34_hnxw_core_069 = input_a[28] ^ input_a[19];
  assign popcount34_hnxw_core_070 = ~input_a[4];
  assign popcount34_hnxw_core_072 = ~(input_a[9] ^ input_a[31]);
  assign popcount34_hnxw_core_073 = input_a[22] ^ input_a[9];
  assign popcount34_hnxw_core_076 = input_a[32] & input_a[23];
  assign popcount34_hnxw_core_079 = ~(input_a[6] & input_a[14]);
  assign popcount34_hnxw_core_080 = input_a[30] | input_a[27];
  assign popcount34_hnxw_core_082 = input_a[0] & input_a[32];
  assign popcount34_hnxw_core_083 = ~(input_a[20] ^ input_a[20]);
  assign popcount34_hnxw_core_084 = input_a[32] ^ input_a[24];
  assign popcount34_hnxw_core_086_not = ~input_a[27];
  assign popcount34_hnxw_core_087 = ~(input_a[4] | input_a[6]);
  assign popcount34_hnxw_core_088_not = ~input_a[22];
  assign popcount34_hnxw_core_089 = ~(input_a[0] & input_a[26]);
  assign popcount34_hnxw_core_090 = ~(input_a[9] | input_a[24]);
  assign popcount34_hnxw_core_092 = ~(input_a[27] | input_a[17]);
  assign popcount34_hnxw_core_093 = input_a[21] | input_a[9];
  assign popcount34_hnxw_core_094 = ~(input_a[33] & input_a[25]);
  assign popcount34_hnxw_core_095 = input_a[32] & input_a[17];
  assign popcount34_hnxw_core_097 = input_a[21] ^ input_a[33];
  assign popcount34_hnxw_core_098 = ~input_a[20];
  assign popcount34_hnxw_core_099 = input_a[19] ^ input_a[12];
  assign popcount34_hnxw_core_100 = ~(input_a[27] & input_a[30]);
  assign popcount34_hnxw_core_101 = ~input_a[33];
  assign popcount34_hnxw_core_102 = input_a[23] & input_a[13];
  assign popcount34_hnxw_core_105 = input_a[25] | input_a[27];
  assign popcount34_hnxw_core_107 = input_a[16] | input_a[27];
  assign popcount34_hnxw_core_109 = ~(input_a[17] ^ input_a[22]);
  assign popcount34_hnxw_core_113 = ~(input_a[14] & input_a[5]);
  assign popcount34_hnxw_core_114 = ~input_a[20];
  assign popcount34_hnxw_core_116 = ~(input_a[19] & input_a[22]);
  assign popcount34_hnxw_core_117 = ~(input_a[23] & input_a[26]);
  assign popcount34_hnxw_core_118 = ~(input_a[8] | input_a[18]);
  assign popcount34_hnxw_core_119 = ~(input_a[24] | input_a[29]);
  assign popcount34_hnxw_core_121 = ~(input_a[2] | input_a[11]);
  assign popcount34_hnxw_core_124 = input_a[8] | input_a[28];
  assign popcount34_hnxw_core_125 = ~(input_a[16] ^ input_a[11]);
  assign popcount34_hnxw_core_126 = ~(input_a[26] & input_a[29]);
  assign popcount34_hnxw_core_128 = ~(input_a[24] ^ input_a[2]);
  assign popcount34_hnxw_core_130 = ~(input_a[1] & input_a[20]);
  assign popcount34_hnxw_core_131 = ~(input_a[5] | input_a[14]);
  assign popcount34_hnxw_core_134 = ~(input_a[1] ^ input_a[18]);
  assign popcount34_hnxw_core_136 = input_a[9] ^ input_a[21];
  assign popcount34_hnxw_core_137 = ~(input_a[5] & input_a[4]);
  assign popcount34_hnxw_core_138 = ~(input_a[12] | input_a[25]);
  assign popcount34_hnxw_core_139 = input_a[32] | input_a[0];
  assign popcount34_hnxw_core_142 = ~(input_a[4] ^ input_a[26]);
  assign popcount34_hnxw_core_144 = ~input_a[11];
  assign popcount34_hnxw_core_145 = ~input_a[13];
  assign popcount34_hnxw_core_149 = ~(input_a[32] ^ input_a[3]);
  assign popcount34_hnxw_core_150 = ~input_a[21];
  assign popcount34_hnxw_core_153 = input_a[11] | input_a[13];
  assign popcount34_hnxw_core_156 = ~(input_a[27] & input_a[23]);
  assign popcount34_hnxw_core_157 = ~input_a[16];
  assign popcount34_hnxw_core_158 = input_a[19] ^ input_a[4];
  assign popcount34_hnxw_core_159 = ~input_a[21];
  assign popcount34_hnxw_core_160 = ~input_a[19];
  assign popcount34_hnxw_core_164 = input_a[31] ^ input_a[3];
  assign popcount34_hnxw_core_167 = ~(input_a[20] | input_a[22]);
  assign popcount34_hnxw_core_169_not = ~input_a[3];
  assign popcount34_hnxw_core_170 = ~input_a[30];
  assign popcount34_hnxw_core_171 = ~(input_a[24] | input_a[32]);
  assign popcount34_hnxw_core_172 = input_a[18] | input_a[10];
  assign popcount34_hnxw_core_173 = ~(input_a[0] | input_a[8]);
  assign popcount34_hnxw_core_175 = ~input_a[26];
  assign popcount34_hnxw_core_176 = ~input_a[27];
  assign popcount34_hnxw_core_177 = ~(input_a[33] ^ input_a[18]);
  assign popcount34_hnxw_core_178 = input_a[11] | input_a[32];
  assign popcount34_hnxw_core_179 = ~(input_a[29] & input_a[12]);
  assign popcount34_hnxw_core_180 = ~(input_a[5] & input_a[22]);
  assign popcount34_hnxw_core_181 = input_a[11] & input_a[32];
  assign popcount34_hnxw_core_183 = ~(input_a[1] | input_a[3]);
  assign popcount34_hnxw_core_184 = ~(input_a[28] & input_a[15]);
  assign popcount34_hnxw_core_185 = ~(input_a[22] ^ input_a[30]);
  assign popcount34_hnxw_core_188 = ~input_a[24];
  assign popcount34_hnxw_core_189 = ~input_a[23];
  assign popcount34_hnxw_core_190 = ~(input_a[5] & input_a[0]);
  assign popcount34_hnxw_core_191 = ~(input_a[1] & input_a[28]);
  assign popcount34_hnxw_core_192 = ~input_a[33];
  assign popcount34_hnxw_core_193 = ~(input_a[8] ^ input_a[15]);
  assign popcount34_hnxw_core_194 = input_a[6] & input_a[9];
  assign popcount34_hnxw_core_196 = input_a[8] & input_a[20];
  assign popcount34_hnxw_core_197 = ~(input_a[17] ^ input_a[7]);
  assign popcount34_hnxw_core_202 = input_a[0] | input_a[9];
  assign popcount34_hnxw_core_203 = input_a[25] ^ input_a[22];
  assign popcount34_hnxw_core_204_not = ~input_a[1];
  assign popcount34_hnxw_core_205 = ~(input_a[20] | input_a[7]);
  assign popcount34_hnxw_core_207 = input_a[4] & input_a[28];
  assign popcount34_hnxw_core_208 = ~(input_a[20] & input_a[29]);
  assign popcount34_hnxw_core_209 = input_a[29] & input_a[8];
  assign popcount34_hnxw_core_212 = input_a[30] | input_a[28];
  assign popcount34_hnxw_core_213 = ~(input_a[0] & input_a[5]);
  assign popcount34_hnxw_core_214 = input_a[21] & input_a[13];
  assign popcount34_hnxw_core_216 = ~input_a[28];
  assign popcount34_hnxw_core_217 = ~(input_a[9] ^ input_a[5]);
  assign popcount34_hnxw_core_219 = ~(input_a[0] & input_a[9]);
  assign popcount34_hnxw_core_221 = ~input_a[25];
  assign popcount34_hnxw_core_222 = input_a[22] & input_a[14];
  assign popcount34_hnxw_core_224 = ~input_a[24];
  assign popcount34_hnxw_core_225 = input_a[9] & input_a[13];
  assign popcount34_hnxw_core_226 = ~input_a[13];
  assign popcount34_hnxw_core_228 = ~(input_a[3] & input_a[9]);
  assign popcount34_hnxw_core_229 = ~(input_a[5] ^ input_a[8]);
  assign popcount34_hnxw_core_230 = ~(input_a[20] | input_a[9]);
  assign popcount34_hnxw_core_231 = input_a[13] & input_a[2];
  assign popcount34_hnxw_core_232 = ~(input_a[1] & input_a[8]);
  assign popcount34_hnxw_core_234 = ~(input_a[23] ^ input_a[0]);
  assign popcount34_hnxw_core_237 = ~(input_a[16] & input_a[22]);
  assign popcount34_hnxw_core_238 = ~(input_a[33] ^ input_a[6]);
  assign popcount34_hnxw_core_239 = ~input_a[13];
  assign popcount34_hnxw_core_244 = ~(input_a[5] & input_a[6]);
  assign popcount34_hnxw_core_246 = ~(input_a[3] ^ input_a[3]);
  assign popcount34_hnxw_core_247 = ~(input_a[22] ^ input_a[5]);
  assign popcount34_hnxw_core_248 = ~(input_a[20] | input_a[0]);
  assign popcount34_hnxw_core_249 = input_a[23] | input_a[30];
  assign popcount34_hnxw_core_250 = ~(input_a[3] ^ input_a[9]);

  assign popcount34_hnxw_out[0] = 1'b0;
  assign popcount34_hnxw_out[1] = 1'b0;
  assign popcount34_hnxw_out[2] = input_a[33];
  assign popcount34_hnxw_out[3] = input_a[12];
  assign popcount34_hnxw_out[4] = 1'b1;
  assign popcount34_hnxw_out[5] = 1'b0;
endmodule