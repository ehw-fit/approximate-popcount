// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=11.5008
// WCE=28.0
// EP=0.99899%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_h47o(input [24:0] input_a, output [4:0] popcount25_h47o_out);
  wire popcount25_h47o_core_027;
  wire popcount25_h47o_core_028_not;
  wire popcount25_h47o_core_029;
  wire popcount25_h47o_core_030;
  wire popcount25_h47o_core_031;
  wire popcount25_h47o_core_032;
  wire popcount25_h47o_core_035;
  wire popcount25_h47o_core_038;
  wire popcount25_h47o_core_041;
  wire popcount25_h47o_core_042;
  wire popcount25_h47o_core_047;
  wire popcount25_h47o_core_048;
  wire popcount25_h47o_core_049;
  wire popcount25_h47o_core_052;
  wire popcount25_h47o_core_053;
  wire popcount25_h47o_core_054;
  wire popcount25_h47o_core_057;
  wire popcount25_h47o_core_059;
  wire popcount25_h47o_core_060;
  wire popcount25_h47o_core_062;
  wire popcount25_h47o_core_063;
  wire popcount25_h47o_core_064;
  wire popcount25_h47o_core_065;
  wire popcount25_h47o_core_066;
  wire popcount25_h47o_core_067;
  wire popcount25_h47o_core_068;
  wire popcount25_h47o_core_069;
  wire popcount25_h47o_core_072;
  wire popcount25_h47o_core_073;
  wire popcount25_h47o_core_074;
  wire popcount25_h47o_core_075;
  wire popcount25_h47o_core_076;
  wire popcount25_h47o_core_077;
  wire popcount25_h47o_core_078;
  wire popcount25_h47o_core_079;
  wire popcount25_h47o_core_080;
  wire popcount25_h47o_core_082;
  wire popcount25_h47o_core_084_not;
  wire popcount25_h47o_core_086;
  wire popcount25_h47o_core_087;
  wire popcount25_h47o_core_089;
  wire popcount25_h47o_core_090_not;
  wire popcount25_h47o_core_092;
  wire popcount25_h47o_core_093;
  wire popcount25_h47o_core_094;
  wire popcount25_h47o_core_095_not;
  wire popcount25_h47o_core_097;
  wire popcount25_h47o_core_098;
  wire popcount25_h47o_core_099;
  wire popcount25_h47o_core_100;
  wire popcount25_h47o_core_103;
  wire popcount25_h47o_core_104;
  wire popcount25_h47o_core_109;
  wire popcount25_h47o_core_110;
  wire popcount25_h47o_core_111_not;
  wire popcount25_h47o_core_112;
  wire popcount25_h47o_core_113;
  wire popcount25_h47o_core_116;
  wire popcount25_h47o_core_118;
  wire popcount25_h47o_core_120;
  wire popcount25_h47o_core_124;
  wire popcount25_h47o_core_125;
  wire popcount25_h47o_core_127;
  wire popcount25_h47o_core_128;
  wire popcount25_h47o_core_129;
  wire popcount25_h47o_core_130_not;
  wire popcount25_h47o_core_134;
  wire popcount25_h47o_core_137;
  wire popcount25_h47o_core_138_not;
  wire popcount25_h47o_core_139;
  wire popcount25_h47o_core_141;
  wire popcount25_h47o_core_142;
  wire popcount25_h47o_core_143;
  wire popcount25_h47o_core_144;
  wire popcount25_h47o_core_146;
  wire popcount25_h47o_core_147;
  wire popcount25_h47o_core_148;
  wire popcount25_h47o_core_149;
  wire popcount25_h47o_core_152;
  wire popcount25_h47o_core_156;
  wire popcount25_h47o_core_157;
  wire popcount25_h47o_core_158;
  wire popcount25_h47o_core_161;
  wire popcount25_h47o_core_162;
  wire popcount25_h47o_core_165;
  wire popcount25_h47o_core_166;
  wire popcount25_h47o_core_170;
  wire popcount25_h47o_core_172;
  wire popcount25_h47o_core_173;
  wire popcount25_h47o_core_176;
  wire popcount25_h47o_core_177;
  wire popcount25_h47o_core_179;
  wire popcount25_h47o_core_180;
  wire popcount25_h47o_core_181;
  wire popcount25_h47o_core_182;
  wire popcount25_h47o_core_183_not;

  assign popcount25_h47o_core_027 = input_a[13] & input_a[22];
  assign popcount25_h47o_core_028_not = ~input_a[20];
  assign popcount25_h47o_core_029 = ~input_a[18];
  assign popcount25_h47o_core_030 = ~(input_a[0] & input_a[22]);
  assign popcount25_h47o_core_031 = input_a[5] & input_a[22];
  assign popcount25_h47o_core_032 = ~(input_a[17] ^ input_a[8]);
  assign popcount25_h47o_core_035 = ~(input_a[12] ^ input_a[7]);
  assign popcount25_h47o_core_038 = input_a[3] & input_a[24];
  assign popcount25_h47o_core_041 = input_a[4] ^ input_a[9];
  assign popcount25_h47o_core_042 = input_a[3] | input_a[22];
  assign popcount25_h47o_core_047 = input_a[21] | input_a[3];
  assign popcount25_h47o_core_048 = ~(input_a[10] ^ input_a[14]);
  assign popcount25_h47o_core_049 = input_a[5] ^ input_a[16];
  assign popcount25_h47o_core_052 = ~(input_a[10] ^ input_a[7]);
  assign popcount25_h47o_core_053 = ~(input_a[4] | input_a[7]);
  assign popcount25_h47o_core_054 = input_a[20] | input_a[17];
  assign popcount25_h47o_core_057 = input_a[1] & input_a[23];
  assign popcount25_h47o_core_059 = input_a[12] | input_a[0];
  assign popcount25_h47o_core_060 = ~input_a[12];
  assign popcount25_h47o_core_062 = input_a[12] | input_a[11];
  assign popcount25_h47o_core_063 = input_a[14] & input_a[10];
  assign popcount25_h47o_core_064 = input_a[18] & input_a[23];
  assign popcount25_h47o_core_065 = input_a[23] ^ input_a[4];
  assign popcount25_h47o_core_066 = ~(input_a[5] & input_a[3]);
  assign popcount25_h47o_core_067 = input_a[8] ^ input_a[12];
  assign popcount25_h47o_core_068 = ~(input_a[5] | input_a[23]);
  assign popcount25_h47o_core_069 = ~(input_a[24] | input_a[6]);
  assign popcount25_h47o_core_072 = ~(input_a[12] ^ input_a[6]);
  assign popcount25_h47o_core_073 = input_a[3] | input_a[21];
  assign popcount25_h47o_core_074 = input_a[11] ^ input_a[15];
  assign popcount25_h47o_core_075 = ~(input_a[20] ^ input_a[1]);
  assign popcount25_h47o_core_076 = input_a[3] & input_a[9];
  assign popcount25_h47o_core_077 = input_a[14] ^ input_a[0];
  assign popcount25_h47o_core_078 = ~(input_a[22] | input_a[2]);
  assign popcount25_h47o_core_079 = input_a[19] ^ input_a[7];
  assign popcount25_h47o_core_080 = input_a[8] | input_a[7];
  assign popcount25_h47o_core_082 = ~input_a[13];
  assign popcount25_h47o_core_084_not = ~input_a[1];
  assign popcount25_h47o_core_086 = input_a[15] ^ input_a[24];
  assign popcount25_h47o_core_087 = input_a[21] ^ input_a[21];
  assign popcount25_h47o_core_089 = input_a[23] ^ input_a[14];
  assign popcount25_h47o_core_090_not = ~input_a[17];
  assign popcount25_h47o_core_092 = ~input_a[12];
  assign popcount25_h47o_core_093 = ~(input_a[9] | input_a[21]);
  assign popcount25_h47o_core_094 = input_a[4] & input_a[4];
  assign popcount25_h47o_core_095_not = ~input_a[15];
  assign popcount25_h47o_core_097 = ~(input_a[22] | input_a[22]);
  assign popcount25_h47o_core_098 = input_a[21] & input_a[14];
  assign popcount25_h47o_core_099 = input_a[15] ^ input_a[11];
  assign popcount25_h47o_core_100 = ~(input_a[10] ^ input_a[24]);
  assign popcount25_h47o_core_103 = ~(input_a[16] ^ input_a[4]);
  assign popcount25_h47o_core_104 = input_a[17] & input_a[20];
  assign popcount25_h47o_core_109 = ~input_a[9];
  assign popcount25_h47o_core_110 = input_a[19] & input_a[5];
  assign popcount25_h47o_core_111_not = ~input_a[13];
  assign popcount25_h47o_core_112 = input_a[15] ^ input_a[4];
  assign popcount25_h47o_core_113 = input_a[0] ^ input_a[4];
  assign popcount25_h47o_core_116 = ~input_a[4];
  assign popcount25_h47o_core_118 = input_a[10] ^ input_a[24];
  assign popcount25_h47o_core_120 = input_a[12] | input_a[6];
  assign popcount25_h47o_core_124 = ~(input_a[10] | input_a[8]);
  assign popcount25_h47o_core_125 = ~(input_a[0] & input_a[2]);
  assign popcount25_h47o_core_127 = input_a[8] | input_a[3];
  assign popcount25_h47o_core_128 = ~(input_a[17] ^ input_a[10]);
  assign popcount25_h47o_core_129 = ~(input_a[2] ^ input_a[14]);
  assign popcount25_h47o_core_130_not = ~input_a[6];
  assign popcount25_h47o_core_134 = ~input_a[13];
  assign popcount25_h47o_core_137 = input_a[10] & input_a[20];
  assign popcount25_h47o_core_138_not = ~input_a[21];
  assign popcount25_h47o_core_139 = input_a[5] | input_a[19];
  assign popcount25_h47o_core_141 = ~(input_a[6] ^ input_a[6]);
  assign popcount25_h47o_core_142 = input_a[17] | input_a[15];
  assign popcount25_h47o_core_143 = ~(input_a[0] & input_a[4]);
  assign popcount25_h47o_core_144 = input_a[12] | input_a[0];
  assign popcount25_h47o_core_146 = ~(input_a[0] ^ input_a[15]);
  assign popcount25_h47o_core_147 = ~(input_a[15] | input_a[21]);
  assign popcount25_h47o_core_148 = input_a[14] ^ input_a[5];
  assign popcount25_h47o_core_149 = input_a[2] & input_a[7];
  assign popcount25_h47o_core_152 = input_a[23] | input_a[16];
  assign popcount25_h47o_core_156 = input_a[13] & input_a[23];
  assign popcount25_h47o_core_157 = input_a[4] ^ input_a[7];
  assign popcount25_h47o_core_158 = input_a[21] & input_a[18];
  assign popcount25_h47o_core_161 = ~(input_a[4] ^ input_a[10]);
  assign popcount25_h47o_core_162 = ~(input_a[3] & input_a[9]);
  assign popcount25_h47o_core_165 = input_a[21] & input_a[4];
  assign popcount25_h47o_core_166 = ~(input_a[8] ^ input_a[22]);
  assign popcount25_h47o_core_170 = ~(input_a[5] & input_a[2]);
  assign popcount25_h47o_core_172 = input_a[4] | input_a[10];
  assign popcount25_h47o_core_173 = input_a[19] ^ input_a[23];
  assign popcount25_h47o_core_176 = ~input_a[21];
  assign popcount25_h47o_core_177 = input_a[19] ^ input_a[11];
  assign popcount25_h47o_core_179 = ~(input_a[17] | input_a[18]);
  assign popcount25_h47o_core_180 = ~(input_a[19] & input_a[20]);
  assign popcount25_h47o_core_181 = input_a[0] ^ input_a[0];
  assign popcount25_h47o_core_182 = ~(input_a[14] | input_a[18]);
  assign popcount25_h47o_core_183_not = ~input_a[20];

  assign popcount25_h47o_out[0] = 1'b1;
  assign popcount25_h47o_out[1] = input_a[21];
  assign popcount25_h47o_out[2] = input_a[7];
  assign popcount25_h47o_out[3] = input_a[0];
  assign popcount25_h47o_out[4] = 1'b1;
endmodule