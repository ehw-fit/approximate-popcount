// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.13137
// WCE=12.0
// EP=0.988012%
// Printed PDK parameters:
//  Area=15388284.0
//  Delay=26605526.0
//  Power=688170.0

module popcount23_6d1u(input [22:0] input_a, output [4:0] popcount23_6d1u_out);
  wire popcount23_6d1u_core_026;
  wire popcount23_6d1u_core_027_not;
  wire popcount23_6d1u_core_029;
  wire popcount23_6d1u_core_030;
  wire popcount23_6d1u_core_033;
  wire popcount23_6d1u_core_034;
  wire popcount23_6d1u_core_035;
  wire popcount23_6d1u_core_036;
  wire popcount23_6d1u_core_037;
  wire popcount23_6d1u_core_038;
  wire popcount23_6d1u_core_039;
  wire popcount23_6d1u_core_043;
  wire popcount23_6d1u_core_045;
  wire popcount23_6d1u_core_046;
  wire popcount23_6d1u_core_047;
  wire popcount23_6d1u_core_048_not;
  wire popcount23_6d1u_core_050;
  wire popcount23_6d1u_core_052;
  wire popcount23_6d1u_core_054;
  wire popcount23_6d1u_core_055_not;
  wire popcount23_6d1u_core_056;
  wire popcount23_6d1u_core_057;
  wire popcount23_6d1u_core_062;
  wire popcount23_6d1u_core_063;
  wire popcount23_6d1u_core_064;
  wire popcount23_6d1u_core_067;
  wire popcount23_6d1u_core_068;
  wire popcount23_6d1u_core_069;
  wire popcount23_6d1u_core_071;
  wire popcount23_6d1u_core_073;
  wire popcount23_6d1u_core_074;
  wire popcount23_6d1u_core_075;
  wire popcount23_6d1u_core_076;
  wire popcount23_6d1u_core_079;
  wire popcount23_6d1u_core_081;
  wire popcount23_6d1u_core_083;
  wire popcount23_6d1u_core_084;
  wire popcount23_6d1u_core_086;
  wire popcount23_6d1u_core_088;
  wire popcount23_6d1u_core_089;
  wire popcount23_6d1u_core_090;
  wire popcount23_6d1u_core_091;
  wire popcount23_6d1u_core_092;
  wire popcount23_6d1u_core_096;
  wire popcount23_6d1u_core_097;
  wire popcount23_6d1u_core_098;
  wire popcount23_6d1u_core_099;
  wire popcount23_6d1u_core_100;
  wire popcount23_6d1u_core_101;
  wire popcount23_6d1u_core_103;
  wire popcount23_6d1u_core_105;
  wire popcount23_6d1u_core_106;
  wire popcount23_6d1u_core_107;
  wire popcount23_6d1u_core_108;
  wire popcount23_6d1u_core_109;
  wire popcount23_6d1u_core_110;
  wire popcount23_6d1u_core_111;
  wire popcount23_6d1u_core_112;
  wire popcount23_6d1u_core_114;
  wire popcount23_6d1u_core_116;
  wire popcount23_6d1u_core_117_not;
  wire popcount23_6d1u_core_118;
  wire popcount23_6d1u_core_119;
  wire popcount23_6d1u_core_120;
  wire popcount23_6d1u_core_121;
  wire popcount23_6d1u_core_122;
  wire popcount23_6d1u_core_124;
  wire popcount23_6d1u_core_125;
  wire popcount23_6d1u_core_127;
  wire popcount23_6d1u_core_128;
  wire popcount23_6d1u_core_129;
  wire popcount23_6d1u_core_131;
  wire popcount23_6d1u_core_133;
  wire popcount23_6d1u_core_138;
  wire popcount23_6d1u_core_140;
  wire popcount23_6d1u_core_141;
  wire popcount23_6d1u_core_143;
  wire popcount23_6d1u_core_144;
  wire popcount23_6d1u_core_145;
  wire popcount23_6d1u_core_146;
  wire popcount23_6d1u_core_149;
  wire popcount23_6d1u_core_150;
  wire popcount23_6d1u_core_151;
  wire popcount23_6d1u_core_152;
  wire popcount23_6d1u_core_153;
  wire popcount23_6d1u_core_154;
  wire popcount23_6d1u_core_155;
  wire popcount23_6d1u_core_157;
  wire popcount23_6d1u_core_159;
  wire popcount23_6d1u_core_160;
  wire popcount23_6d1u_core_162;
  wire popcount23_6d1u_core_163;
  wire popcount23_6d1u_core_164;
  wire popcount23_6d1u_core_165;
  wire popcount23_6d1u_core_166;
  wire popcount23_6d1u_core_167;
  wire popcount23_6d1u_core_168;

  assign popcount23_6d1u_core_026 = input_a[7] & input_a[3];
  assign popcount23_6d1u_core_027_not = ~input_a[8];
  assign popcount23_6d1u_core_029 = ~(input_a[2] & input_a[19]);
  assign popcount23_6d1u_core_030 = input_a[22] & input_a[13];
  assign popcount23_6d1u_core_033 = input_a[4] | input_a[21];
  assign popcount23_6d1u_core_034 = input_a[16] & input_a[20];
  assign popcount23_6d1u_core_035 = popcount23_6d1u_core_026 ^ popcount23_6d1u_core_030;
  assign popcount23_6d1u_core_036 = popcount23_6d1u_core_026 & popcount23_6d1u_core_030;
  assign popcount23_6d1u_core_037 = popcount23_6d1u_core_035 ^ popcount23_6d1u_core_034;
  assign popcount23_6d1u_core_038 = popcount23_6d1u_core_035 & popcount23_6d1u_core_034;
  assign popcount23_6d1u_core_039 = popcount23_6d1u_core_036 | popcount23_6d1u_core_038;
  assign popcount23_6d1u_core_043 = input_a[18] & input_a[1];
  assign popcount23_6d1u_core_045 = input_a[10] & input_a[6];
  assign popcount23_6d1u_core_046 = popcount23_6d1u_core_043 ^ popcount23_6d1u_core_045;
  assign popcount23_6d1u_core_047 = popcount23_6d1u_core_043 & popcount23_6d1u_core_045;
  assign popcount23_6d1u_core_048_not = ~input_a[10];
  assign popcount23_6d1u_core_050 = input_a[7] ^ input_a[11];
  assign popcount23_6d1u_core_052 = ~input_a[5];
  assign popcount23_6d1u_core_054 = ~(input_a[3] | input_a[14]);
  assign popcount23_6d1u_core_055_not = ~input_a[7];
  assign popcount23_6d1u_core_056 = popcount23_6d1u_core_046 ^ input_a[15];
  assign popcount23_6d1u_core_057 = popcount23_6d1u_core_046 & input_a[15];
  assign popcount23_6d1u_core_062 = ~(input_a[1] ^ input_a[15]);
  assign popcount23_6d1u_core_063 = popcount23_6d1u_core_047 | popcount23_6d1u_core_057;
  assign popcount23_6d1u_core_064 = ~(input_a[17] ^ input_a[16]);
  assign popcount23_6d1u_core_067 = ~(input_a[15] | input_a[7]);
  assign popcount23_6d1u_core_068 = ~(input_a[22] ^ input_a[0]);
  assign popcount23_6d1u_core_069 = popcount23_6d1u_core_037 & popcount23_6d1u_core_056;
  assign popcount23_6d1u_core_071 = input_a[21] & input_a[7];
  assign popcount23_6d1u_core_073 = popcount23_6d1u_core_039 ^ popcount23_6d1u_core_063;
  assign popcount23_6d1u_core_074 = popcount23_6d1u_core_039 & popcount23_6d1u_core_063;
  assign popcount23_6d1u_core_075 = popcount23_6d1u_core_073 ^ popcount23_6d1u_core_069;
  assign popcount23_6d1u_core_076 = popcount23_6d1u_core_073 & popcount23_6d1u_core_069;
  assign popcount23_6d1u_core_079 = input_a[6] & input_a[15];
  assign popcount23_6d1u_core_081 = ~(input_a[20] | input_a[19]);
  assign popcount23_6d1u_core_083 = ~(input_a[15] | input_a[13]);
  assign popcount23_6d1u_core_084 = input_a[17] & input_a[19];
  assign popcount23_6d1u_core_086 = input_a[4] | input_a[0];
  assign popcount23_6d1u_core_088 = ~(input_a[21] | input_a[10]);
  assign popcount23_6d1u_core_089 = ~(input_a[11] ^ input_a[10]);
  assign popcount23_6d1u_core_090 = input_a[14] & input_a[9];
  assign popcount23_6d1u_core_091 = input_a[0] & input_a[19];
  assign popcount23_6d1u_core_092 = input_a[20] | input_a[22];
  assign popcount23_6d1u_core_096 = input_a[2] & input_a[0];
  assign popcount23_6d1u_core_097 = ~(popcount23_6d1u_core_084 & popcount23_6d1u_core_090);
  assign popcount23_6d1u_core_098 = popcount23_6d1u_core_084 & popcount23_6d1u_core_090;
  assign popcount23_6d1u_core_099 = popcount23_6d1u_core_097 ^ popcount23_6d1u_core_096;
  assign popcount23_6d1u_core_100 = input_a[2] & input_a[0];
  assign popcount23_6d1u_core_101 = popcount23_6d1u_core_098 | popcount23_6d1u_core_100;
  assign popcount23_6d1u_core_103 = ~(input_a[14] ^ input_a[19]);
  assign popcount23_6d1u_core_105 = ~(input_a[12] ^ input_a[8]);
  assign popcount23_6d1u_core_106 = ~(input_a[15] | input_a[22]);
  assign popcount23_6d1u_core_107 = ~(input_a[21] ^ input_a[6]);
  assign popcount23_6d1u_core_108 = input_a[21] ^ input_a[1];
  assign popcount23_6d1u_core_109 = ~(input_a[21] | input_a[12]);
  assign popcount23_6d1u_core_110 = ~(input_a[10] ^ input_a[9]);
  assign popcount23_6d1u_core_111 = ~(input_a[10] ^ input_a[7]);
  assign popcount23_6d1u_core_112 = ~(input_a[13] | input_a[2]);
  assign popcount23_6d1u_core_114 = input_a[19] & input_a[11];
  assign popcount23_6d1u_core_116 = ~(input_a[20] & input_a[7]);
  assign popcount23_6d1u_core_117_not = ~input_a[12];
  assign popcount23_6d1u_core_118 = input_a[2] | input_a[3];
  assign popcount23_6d1u_core_119 = ~(input_a[4] & input_a[6]);
  assign popcount23_6d1u_core_120 = ~(input_a[9] & input_a[20]);
  assign popcount23_6d1u_core_121 = ~input_a[5];
  assign popcount23_6d1u_core_122 = ~(input_a[6] | input_a[5]);
  assign popcount23_6d1u_core_124 = input_a[3] & input_a[2];
  assign popcount23_6d1u_core_125 = ~(input_a[17] & input_a[19]);
  assign popcount23_6d1u_core_127 = ~(input_a[7] & input_a[16]);
  assign popcount23_6d1u_core_128 = ~(input_a[13] ^ input_a[6]);
  assign popcount23_6d1u_core_129 = ~input_a[3];
  assign popcount23_6d1u_core_131 = ~(input_a[13] ^ input_a[0]);
  assign popcount23_6d1u_core_133 = popcount23_6d1u_core_099 | popcount23_6d1u_core_121;
  assign popcount23_6d1u_core_138 = popcount23_6d1u_core_101 ^ input_a[5];
  assign popcount23_6d1u_core_140 = popcount23_6d1u_core_138 ^ popcount23_6d1u_core_133;
  assign popcount23_6d1u_core_141 = ~(input_a[7] & input_a[5]);
  assign popcount23_6d1u_core_143 = input_a[19] & input_a[6];
  assign popcount23_6d1u_core_144 = ~input_a[21];
  assign popcount23_6d1u_core_145 = input_a[5] | popcount23_6d1u_core_101;
  assign popcount23_6d1u_core_146 = ~(input_a[3] | input_a[10]);
  assign popcount23_6d1u_core_149 = input_a[4] & input_a[22];
  assign popcount23_6d1u_core_150 = ~(input_a[0] & input_a[5]);
  assign popcount23_6d1u_core_151 = ~(input_a[21] | input_a[21]);
  assign popcount23_6d1u_core_152 = input_a[21] | input_a[9];
  assign popcount23_6d1u_core_153 = input_a[7] | input_a[19];
  assign popcount23_6d1u_core_154 = input_a[0] & input_a[10];
  assign popcount23_6d1u_core_155 = popcount23_6d1u_core_075 ^ popcount23_6d1u_core_140;
  assign popcount23_6d1u_core_157 = ~popcount23_6d1u_core_155;
  assign popcount23_6d1u_core_159 = popcount23_6d1u_core_075 | popcount23_6d1u_core_155;
  assign popcount23_6d1u_core_160 = input_a[5] | popcount23_6d1u_core_145;
  assign popcount23_6d1u_core_162 = input_a[19] ^ input_a[10];
  assign popcount23_6d1u_core_163 = popcount23_6d1u_core_160 & popcount23_6d1u_core_159;
  assign popcount23_6d1u_core_164 = popcount23_6d1u_core_074 | popcount23_6d1u_core_163;
  assign popcount23_6d1u_core_165 = input_a[13] ^ input_a[12];
  assign popcount23_6d1u_core_166 = ~(input_a[13] & input_a[11]);
  assign popcount23_6d1u_core_167 = ~(input_a[15] ^ input_a[0]);
  assign popcount23_6d1u_core_168 = ~(input_a[22] ^ input_a[5]);

  assign popcount23_6d1u_out[0] = input_a[4];
  assign popcount23_6d1u_out[1] = popcount23_6d1u_core_140;
  assign popcount23_6d1u_out[2] = popcount23_6d1u_core_157;
  assign popcount23_6d1u_out[3] = popcount23_6d1u_core_076;
  assign popcount23_6d1u_out[4] = popcount23_6d1u_core_164;
endmodule