// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.78923
// WCE=25.0
// EP=0.824561%
// Printed PDK parameters:
//  Area=53341019.0
//  Delay=69420144.0
//  Power=2272200.0

module popcount36_pocl(input [35:0] input_a, output [5:0] popcount36_pocl_out);
  wire popcount36_pocl_core_038;
  wire popcount36_pocl_core_039;
  wire popcount36_pocl_core_040;
  wire popcount36_pocl_core_041;
  wire popcount36_pocl_core_043;
  wire popcount36_pocl_core_044;
  wire popcount36_pocl_core_045;
  wire popcount36_pocl_core_046;
  wire popcount36_pocl_core_049;
  wire popcount36_pocl_core_050;
  wire popcount36_pocl_core_051;
  wire popcount36_pocl_core_054;
  wire popcount36_pocl_core_057;
  wire popcount36_pocl_core_059;
  wire popcount36_pocl_core_060;
  wire popcount36_pocl_core_061;
  wire popcount36_pocl_core_062;
  wire popcount36_pocl_core_063;
  wire popcount36_pocl_core_066;
  wire popcount36_pocl_core_067;
  wire popcount36_pocl_core_068;
  wire popcount36_pocl_core_069;
  wire popcount36_pocl_core_071;
  wire popcount36_pocl_core_073;
  wire popcount36_pocl_core_074;
  wire popcount36_pocl_core_075;
  wire popcount36_pocl_core_076;
  wire popcount36_pocl_core_077;
  wire popcount36_pocl_core_080;
  wire popcount36_pocl_core_081;
  wire popcount36_pocl_core_083;
  wire popcount36_pocl_core_084;
  wire popcount36_pocl_core_085;
  wire popcount36_pocl_core_086;
  wire popcount36_pocl_core_087;
  wire popcount36_pocl_core_090;
  wire popcount36_pocl_core_091;
  wire popcount36_pocl_core_092;
  wire popcount36_pocl_core_093_not;
  wire popcount36_pocl_core_094;
  wire popcount36_pocl_core_095;
  wire popcount36_pocl_core_096;
  wire popcount36_pocl_core_097;
  wire popcount36_pocl_core_099;
  wire popcount36_pocl_core_100;
  wire popcount36_pocl_core_101;
  wire popcount36_pocl_core_103;
  wire popcount36_pocl_core_104;
  wire popcount36_pocl_core_105;
  wire popcount36_pocl_core_109;
  wire popcount36_pocl_core_112;
  wire popcount36_pocl_core_113;
  wire popcount36_pocl_core_115;
  wire popcount36_pocl_core_116;
  wire popcount36_pocl_core_117;
  wire popcount36_pocl_core_118;
  wire popcount36_pocl_core_119;
  wire popcount36_pocl_core_121;
  wire popcount36_pocl_core_124;
  wire popcount36_pocl_core_125;
  wire popcount36_pocl_core_126;
  wire popcount36_pocl_core_127;
  wire popcount36_pocl_core_128;
  wire popcount36_pocl_core_129;
  wire popcount36_pocl_core_130;
  wire popcount36_pocl_core_131;
  wire popcount36_pocl_core_132;
  wire popcount36_pocl_core_133;
  wire popcount36_pocl_core_134;
  wire popcount36_pocl_core_136;
  wire popcount36_pocl_core_137;
  wire popcount36_pocl_core_138;
  wire popcount36_pocl_core_140;
  wire popcount36_pocl_core_142;
  wire popcount36_pocl_core_143;
  wire popcount36_pocl_core_144;
  wire popcount36_pocl_core_147;
  wire popcount36_pocl_core_148;
  wire popcount36_pocl_core_149;
  wire popcount36_pocl_core_151;
  wire popcount36_pocl_core_153;
  wire popcount36_pocl_core_155;
  wire popcount36_pocl_core_157;
  wire popcount36_pocl_core_158;
  wire popcount36_pocl_core_160;
  wire popcount36_pocl_core_161;
  wire popcount36_pocl_core_162;
  wire popcount36_pocl_core_163_not;
  wire popcount36_pocl_core_164;
  wire popcount36_pocl_core_168;
  wire popcount36_pocl_core_169;
  wire popcount36_pocl_core_171;
  wire popcount36_pocl_core_172;
  wire popcount36_pocl_core_174;
  wire popcount36_pocl_core_175;
  wire popcount36_pocl_core_177;
  wire popcount36_pocl_core_180;
  wire popcount36_pocl_core_184;
  wire popcount36_pocl_core_185;
  wire popcount36_pocl_core_188;
  wire popcount36_pocl_core_189;
  wire popcount36_pocl_core_190;
  wire popcount36_pocl_core_191;
  wire popcount36_pocl_core_192;
  wire popcount36_pocl_core_193;
  wire popcount36_pocl_core_195;
  wire popcount36_pocl_core_197;
  wire popcount36_pocl_core_198;
  wire popcount36_pocl_core_199;
  wire popcount36_pocl_core_201;
  wire popcount36_pocl_core_208;
  wire popcount36_pocl_core_210;
  wire popcount36_pocl_core_211;
  wire popcount36_pocl_core_212;
  wire popcount36_pocl_core_213;
  wire popcount36_pocl_core_214;
  wire popcount36_pocl_core_215_not;
  wire popcount36_pocl_core_216;
  wire popcount36_pocl_core_217;
  wire popcount36_pocl_core_219;
  wire popcount36_pocl_core_222;
  wire popcount36_pocl_core_223;
  wire popcount36_pocl_core_224;
  wire popcount36_pocl_core_225;
  wire popcount36_pocl_core_226;
  wire popcount36_pocl_core_227;
  wire popcount36_pocl_core_228;
  wire popcount36_pocl_core_230;
  wire popcount36_pocl_core_231;
  wire popcount36_pocl_core_232;
  wire popcount36_pocl_core_233;
  wire popcount36_pocl_core_234;
  wire popcount36_pocl_core_235;
  wire popcount36_pocl_core_236;
  wire popcount36_pocl_core_237;
  wire popcount36_pocl_core_238;
  wire popcount36_pocl_core_239;
  wire popcount36_pocl_core_241;
  wire popcount36_pocl_core_243;
  wire popcount36_pocl_core_244;
  wire popcount36_pocl_core_245;
  wire popcount36_pocl_core_247;
  wire popcount36_pocl_core_249;
  wire popcount36_pocl_core_252;
  wire popcount36_pocl_core_253;
  wire popcount36_pocl_core_254;
  wire popcount36_pocl_core_255;
  wire popcount36_pocl_core_256;
  wire popcount36_pocl_core_257;
  wire popcount36_pocl_core_258;
  wire popcount36_pocl_core_259;
  wire popcount36_pocl_core_260;
  wire popcount36_pocl_core_261;
  wire popcount36_pocl_core_262;
  wire popcount36_pocl_core_263;
  wire popcount36_pocl_core_264;
  wire popcount36_pocl_core_265;
  wire popcount36_pocl_core_266;
  wire popcount36_pocl_core_268;
  wire popcount36_pocl_core_269;
  wire popcount36_pocl_core_270;
  wire popcount36_pocl_core_271;
  wire popcount36_pocl_core_272;
  wire popcount36_pocl_core_274;
  wire popcount36_pocl_core_275;
  wire popcount36_pocl_core_276;

  assign popcount36_pocl_core_038 = input_a[17] | input_a[0];
  assign popcount36_pocl_core_039 = input_a[6] & input_a[15];
  assign popcount36_pocl_core_040 = input_a[31] ^ input_a[18];
  assign popcount36_pocl_core_041 = input_a[28] & input_a[33];
  assign popcount36_pocl_core_043 = input_a[3] & input_a[23];
  assign popcount36_pocl_core_044 = popcount36_pocl_core_039 ^ popcount36_pocl_core_041;
  assign popcount36_pocl_core_045 = popcount36_pocl_core_039 & popcount36_pocl_core_041;
  assign popcount36_pocl_core_046 = popcount36_pocl_core_044 | popcount36_pocl_core_043;
  assign popcount36_pocl_core_049 = ~(input_a[12] & input_a[22]);
  assign popcount36_pocl_core_050 = input_a[34] & input_a[11];
  assign popcount36_pocl_core_051 = input_a[29] | input_a[7];
  assign popcount36_pocl_core_054 = input_a[1] & popcount36_pocl_core_051;
  assign popcount36_pocl_core_057 = ~input_a[12];
  assign popcount36_pocl_core_059 = popcount36_pocl_core_050 ^ popcount36_pocl_core_054;
  assign popcount36_pocl_core_060 = popcount36_pocl_core_050 & popcount36_pocl_core_054;
  assign popcount36_pocl_core_061 = popcount36_pocl_core_059 ^ popcount36_pocl_core_049;
  assign popcount36_pocl_core_062 = popcount36_pocl_core_059 & popcount36_pocl_core_049;
  assign popcount36_pocl_core_063 = popcount36_pocl_core_060 | popcount36_pocl_core_062;
  assign popcount36_pocl_core_066 = input_a[22] | popcount36_pocl_core_057;
  assign popcount36_pocl_core_067 = ~(input_a[20] | input_a[23]);
  assign popcount36_pocl_core_068 = popcount36_pocl_core_046 ^ popcount36_pocl_core_061;
  assign popcount36_pocl_core_069 = popcount36_pocl_core_046 & popcount36_pocl_core_061;
  assign popcount36_pocl_core_071 = ~(input_a[31] ^ input_a[2]);
  assign popcount36_pocl_core_073 = popcount36_pocl_core_045 ^ popcount36_pocl_core_063;
  assign popcount36_pocl_core_074 = popcount36_pocl_core_045 & popcount36_pocl_core_063;
  assign popcount36_pocl_core_075 = popcount36_pocl_core_073 ^ popcount36_pocl_core_069;
  assign popcount36_pocl_core_076 = popcount36_pocl_core_073 & popcount36_pocl_core_069;
  assign popcount36_pocl_core_077 = popcount36_pocl_core_074 | popcount36_pocl_core_076;
  assign popcount36_pocl_core_080 = input_a[0] & input_a[18];
  assign popcount36_pocl_core_081 = input_a[3] ^ input_a[24];
  assign popcount36_pocl_core_083 = input_a[34] | input_a[19];
  assign popcount36_pocl_core_084 = ~(input_a[18] ^ input_a[5]);
  assign popcount36_pocl_core_085 = input_a[29] ^ input_a[28];
  assign popcount36_pocl_core_086 = input_a[8] | input_a[7];
  assign popcount36_pocl_core_087 = input_a[5] ^ input_a[13];
  assign popcount36_pocl_core_090 = ~input_a[33];
  assign popcount36_pocl_core_091 = input_a[13] ^ input_a[14];
  assign popcount36_pocl_core_092 = input_a[13] & input_a[14];
  assign popcount36_pocl_core_093_not = ~input_a[35];
  assign popcount36_pocl_core_094 = ~input_a[12];
  assign popcount36_pocl_core_095 = input_a[15] ^ input_a[13];
  assign popcount36_pocl_core_096 = ~(input_a[15] & input_a[28]);
  assign popcount36_pocl_core_097 = input_a[24] ^ input_a[18];
  assign popcount36_pocl_core_099 = input_a[22] & input_a[20];
  assign popcount36_pocl_core_100 = popcount36_pocl_core_091 & input_a[0];
  assign popcount36_pocl_core_101 = ~popcount36_pocl_core_092;
  assign popcount36_pocl_core_103 = popcount36_pocl_core_101 ^ popcount36_pocl_core_100;
  assign popcount36_pocl_core_104 = input_a[0] & popcount36_pocl_core_100;
  assign popcount36_pocl_core_105 = popcount36_pocl_core_092 | popcount36_pocl_core_104;
  assign popcount36_pocl_core_109 = input_a[32] & input_a[8];
  assign popcount36_pocl_core_112 = popcount36_pocl_core_103 ^ popcount36_pocl_core_109;
  assign popcount36_pocl_core_113 = popcount36_pocl_core_103 & popcount36_pocl_core_109;
  assign popcount36_pocl_core_115 = input_a[12] ^ popcount36_pocl_core_105;
  assign popcount36_pocl_core_116 = input_a[12] & popcount36_pocl_core_105;
  assign popcount36_pocl_core_117 = popcount36_pocl_core_115 ^ popcount36_pocl_core_113;
  assign popcount36_pocl_core_118 = input_a[12] & popcount36_pocl_core_113;
  assign popcount36_pocl_core_119 = popcount36_pocl_core_116 | popcount36_pocl_core_118;
  assign popcount36_pocl_core_121 = ~(input_a[12] ^ input_a[9]);
  assign popcount36_pocl_core_124 = popcount36_pocl_core_068 ^ popcount36_pocl_core_112;
  assign popcount36_pocl_core_125 = popcount36_pocl_core_068 & popcount36_pocl_core_112;
  assign popcount36_pocl_core_126 = popcount36_pocl_core_124 ^ popcount36_pocl_core_066;
  assign popcount36_pocl_core_127 = popcount36_pocl_core_124 & popcount36_pocl_core_066;
  assign popcount36_pocl_core_128 = popcount36_pocl_core_125 | popcount36_pocl_core_127;
  assign popcount36_pocl_core_129 = popcount36_pocl_core_075 ^ popcount36_pocl_core_117;
  assign popcount36_pocl_core_130 = popcount36_pocl_core_075 & popcount36_pocl_core_117;
  assign popcount36_pocl_core_131 = popcount36_pocl_core_129 ^ popcount36_pocl_core_128;
  assign popcount36_pocl_core_132 = popcount36_pocl_core_129 & popcount36_pocl_core_128;
  assign popcount36_pocl_core_133 = popcount36_pocl_core_130 | popcount36_pocl_core_132;
  assign popcount36_pocl_core_134 = popcount36_pocl_core_077 ^ popcount36_pocl_core_119;
  assign popcount36_pocl_core_136 = popcount36_pocl_core_134 ^ popcount36_pocl_core_133;
  assign popcount36_pocl_core_137 = popcount36_pocl_core_134 & popcount36_pocl_core_133;
  assign popcount36_pocl_core_138 = popcount36_pocl_core_077 | popcount36_pocl_core_137;
  assign popcount36_pocl_core_140 = ~input_a[35];
  assign popcount36_pocl_core_142 = input_a[6] & input_a[34];
  assign popcount36_pocl_core_143 = input_a[16] | input_a[34];
  assign popcount36_pocl_core_144 = input_a[17] | input_a[26];
  assign popcount36_pocl_core_147 = input_a[10] & input_a[20];
  assign popcount36_pocl_core_148 = ~(input_a[31] ^ input_a[23]);
  assign popcount36_pocl_core_149 = ~(input_a[31] | input_a[34]);
  assign popcount36_pocl_core_151 = input_a[0] ^ input_a[17];
  assign popcount36_pocl_core_153 = ~(input_a[2] & input_a[10]);
  assign popcount36_pocl_core_155 = ~(input_a[13] & input_a[30]);
  assign popcount36_pocl_core_157 = ~(input_a[26] | input_a[1]);
  assign popcount36_pocl_core_158 = input_a[31] & input_a[27];
  assign popcount36_pocl_core_160 = input_a[9] & input_a[19];
  assign popcount36_pocl_core_161 = popcount36_pocl_core_158 | popcount36_pocl_core_160;
  assign popcount36_pocl_core_162 = input_a[13] | input_a[14];
  assign popcount36_pocl_core_163_not = ~input_a[2];
  assign popcount36_pocl_core_164 = input_a[8] & input_a[18];
  assign popcount36_pocl_core_168 = input_a[11] & input_a[5];
  assign popcount36_pocl_core_169 = input_a[23] & input_a[35];
  assign popcount36_pocl_core_171 = ~input_a[22];
  assign popcount36_pocl_core_172 = input_a[21] | input_a[18];
  assign popcount36_pocl_core_174 = popcount36_pocl_core_147 ^ popcount36_pocl_core_161;
  assign popcount36_pocl_core_175 = popcount36_pocl_core_147 & popcount36_pocl_core_161;
  assign popcount36_pocl_core_177 = ~(input_a[7] ^ input_a[4]);
  assign popcount36_pocl_core_180 = input_a[32] | input_a[19];
  assign popcount36_pocl_core_184 = input_a[29] | input_a[3];
  assign popcount36_pocl_core_185 = ~(input_a[11] ^ input_a[5]);
  assign popcount36_pocl_core_188 = input_a[27] | input_a[33];
  assign popcount36_pocl_core_189 = input_a[35] & input_a[4];
  assign popcount36_pocl_core_190 = input_a[1] & input_a[20];
  assign popcount36_pocl_core_191 = ~input_a[15];
  assign popcount36_pocl_core_192 = input_a[24] ^ popcount36_pocl_core_189;
  assign popcount36_pocl_core_193 = input_a[24] & popcount36_pocl_core_189;
  assign popcount36_pocl_core_195 = ~input_a[24];
  assign popcount36_pocl_core_197 = ~(input_a[3] | input_a[21]);
  assign popcount36_pocl_core_198 = input_a[16] & input_a[30];
  assign popcount36_pocl_core_199 = ~(input_a[5] | input_a[25]);
  assign popcount36_pocl_core_201 = input_a[28] ^ input_a[29];
  assign popcount36_pocl_core_208 = ~(input_a[11] & input_a[33]);
  assign popcount36_pocl_core_210 = ~input_a[17];
  assign popcount36_pocl_core_211 = ~(input_a[7] | input_a[20]);
  assign popcount36_pocl_core_212 = ~(input_a[16] ^ input_a[33]);
  assign popcount36_pocl_core_213 = ~(input_a[10] ^ input_a[24]);
  assign popcount36_pocl_core_214 = input_a[1] | input_a[10];
  assign popcount36_pocl_core_215_not = ~input_a[35];
  assign popcount36_pocl_core_216 = popcount36_pocl_core_192 ^ popcount36_pocl_core_198;
  assign popcount36_pocl_core_217 = popcount36_pocl_core_192 & popcount36_pocl_core_198;
  assign popcount36_pocl_core_219 = ~(input_a[20] & input_a[23]);
  assign popcount36_pocl_core_222 = ~(input_a[32] | input_a[31]);
  assign popcount36_pocl_core_223 = popcount36_pocl_core_193 | popcount36_pocl_core_217;
  assign popcount36_pocl_core_224 = ~input_a[18];
  assign popcount36_pocl_core_225 = ~input_a[26];
  assign popcount36_pocl_core_226 = ~input_a[35];
  assign popcount36_pocl_core_227 = ~(input_a[28] ^ input_a[5]);
  assign popcount36_pocl_core_228 = ~(input_a[31] | input_a[9]);
  assign popcount36_pocl_core_230 = popcount36_pocl_core_174 ^ popcount36_pocl_core_216;
  assign popcount36_pocl_core_231 = popcount36_pocl_core_174 & popcount36_pocl_core_216;
  assign popcount36_pocl_core_232 = popcount36_pocl_core_230 ^ popcount36_pocl_core_172;
  assign popcount36_pocl_core_233 = popcount36_pocl_core_230 & popcount36_pocl_core_172;
  assign popcount36_pocl_core_234 = popcount36_pocl_core_231 | popcount36_pocl_core_233;
  assign popcount36_pocl_core_235 = popcount36_pocl_core_175 ^ popcount36_pocl_core_223;
  assign popcount36_pocl_core_236 = popcount36_pocl_core_175 & popcount36_pocl_core_223;
  assign popcount36_pocl_core_237 = popcount36_pocl_core_235 ^ popcount36_pocl_core_234;
  assign popcount36_pocl_core_238 = popcount36_pocl_core_235 & popcount36_pocl_core_234;
  assign popcount36_pocl_core_239 = popcount36_pocl_core_236 | popcount36_pocl_core_238;
  assign popcount36_pocl_core_241 = input_a[25] & input_a[8];
  assign popcount36_pocl_core_243 = input_a[15] ^ input_a[20];
  assign popcount36_pocl_core_244 = input_a[16] ^ input_a[5];
  assign popcount36_pocl_core_245 = ~(input_a[5] & input_a[6]);
  assign popcount36_pocl_core_247 = ~(input_a[4] | input_a[1]);
  assign popcount36_pocl_core_249 = input_a[5] | input_a[23];
  assign popcount36_pocl_core_252 = popcount36_pocl_core_126 ^ popcount36_pocl_core_232;
  assign popcount36_pocl_core_253 = popcount36_pocl_core_126 & popcount36_pocl_core_232;
  assign popcount36_pocl_core_254 = ~(popcount36_pocl_core_252 & popcount36_pocl_core_066);
  assign popcount36_pocl_core_255 = popcount36_pocl_core_252 & popcount36_pocl_core_066;
  assign popcount36_pocl_core_256 = popcount36_pocl_core_253 | popcount36_pocl_core_255;
  assign popcount36_pocl_core_257 = popcount36_pocl_core_131 ^ popcount36_pocl_core_237;
  assign popcount36_pocl_core_258 = popcount36_pocl_core_131 & popcount36_pocl_core_237;
  assign popcount36_pocl_core_259 = popcount36_pocl_core_257 ^ popcount36_pocl_core_256;
  assign popcount36_pocl_core_260 = popcount36_pocl_core_257 & popcount36_pocl_core_256;
  assign popcount36_pocl_core_261 = popcount36_pocl_core_258 | popcount36_pocl_core_260;
  assign popcount36_pocl_core_262 = popcount36_pocl_core_136 ^ popcount36_pocl_core_239;
  assign popcount36_pocl_core_263 = popcount36_pocl_core_136 & popcount36_pocl_core_239;
  assign popcount36_pocl_core_264 = popcount36_pocl_core_262 ^ popcount36_pocl_core_261;
  assign popcount36_pocl_core_265 = popcount36_pocl_core_262 & popcount36_pocl_core_261;
  assign popcount36_pocl_core_266 = popcount36_pocl_core_263 | popcount36_pocl_core_265;
  assign popcount36_pocl_core_268 = input_a[32] | input_a[18];
  assign popcount36_pocl_core_269 = popcount36_pocl_core_138 | popcount36_pocl_core_266;
  assign popcount36_pocl_core_270 = ~(input_a[7] & input_a[11]);
  assign popcount36_pocl_core_271 = input_a[8] ^ input_a[5];
  assign popcount36_pocl_core_272 = input_a[19] | input_a[14];
  assign popcount36_pocl_core_274 = ~(input_a[14] ^ input_a[8]);
  assign popcount36_pocl_core_275 = ~(input_a[3] | input_a[2]);
  assign popcount36_pocl_core_276 = input_a[6] | input_a[2];

  assign popcount36_pocl_out[0] = popcount36_pocl_core_264;
  assign popcount36_pocl_out[1] = popcount36_pocl_core_254;
  assign popcount36_pocl_out[2] = popcount36_pocl_core_259;
  assign popcount36_pocl_out[3] = popcount36_pocl_core_264;
  assign popcount36_pocl_out[4] = popcount36_pocl_core_269;
  assign popcount36_pocl_out[5] = 1'b0;
endmodule