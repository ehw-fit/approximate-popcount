// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.66933
// WCE=15.0
// EP=0.938547%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_bwjn(input [21:0] input_a, output [4:0] popcount22_bwjn_out);
  wire popcount22_bwjn_core_027;
  wire popcount22_bwjn_core_028;
  wire popcount22_bwjn_core_030;
  wire popcount22_bwjn_core_031;
  wire popcount22_bwjn_core_033;
  wire popcount22_bwjn_core_034;
  wire popcount22_bwjn_core_038;
  wire popcount22_bwjn_core_039;
  wire popcount22_bwjn_core_040;
  wire popcount22_bwjn_core_042_not;
  wire popcount22_bwjn_core_043;
  wire popcount22_bwjn_core_044;
  wire popcount22_bwjn_core_046;
  wire popcount22_bwjn_core_048;
  wire popcount22_bwjn_core_051_not;
  wire popcount22_bwjn_core_053;
  wire popcount22_bwjn_core_055;
  wire popcount22_bwjn_core_056;
  wire popcount22_bwjn_core_057;
  wire popcount22_bwjn_core_058;
  wire popcount22_bwjn_core_059;
  wire popcount22_bwjn_core_060;
  wire popcount22_bwjn_core_062;
  wire popcount22_bwjn_core_063;
  wire popcount22_bwjn_core_064_not;
  wire popcount22_bwjn_core_065_not;
  wire popcount22_bwjn_core_067;
  wire popcount22_bwjn_core_070;
  wire popcount22_bwjn_core_072;
  wire popcount22_bwjn_core_074;
  wire popcount22_bwjn_core_077;
  wire popcount22_bwjn_core_078;
  wire popcount22_bwjn_core_079;
  wire popcount22_bwjn_core_080;
  wire popcount22_bwjn_core_081_not;
  wire popcount22_bwjn_core_083;
  wire popcount22_bwjn_core_086;
  wire popcount22_bwjn_core_088_not;
  wire popcount22_bwjn_core_090;
  wire popcount22_bwjn_core_091;
  wire popcount22_bwjn_core_093;
  wire popcount22_bwjn_core_094;
  wire popcount22_bwjn_core_099;
  wire popcount22_bwjn_core_102;
  wire popcount22_bwjn_core_103;
  wire popcount22_bwjn_core_105;
  wire popcount22_bwjn_core_106;
  wire popcount22_bwjn_core_107;
  wire popcount22_bwjn_core_112;
  wire popcount22_bwjn_core_113;
  wire popcount22_bwjn_core_116;
  wire popcount22_bwjn_core_117;
  wire popcount22_bwjn_core_121;
  wire popcount22_bwjn_core_122;
  wire popcount22_bwjn_core_124;
  wire popcount22_bwjn_core_125;
  wire popcount22_bwjn_core_127;
  wire popcount22_bwjn_core_129;
  wire popcount22_bwjn_core_133;
  wire popcount22_bwjn_core_134;
  wire popcount22_bwjn_core_136;
  wire popcount22_bwjn_core_137;
  wire popcount22_bwjn_core_139;
  wire popcount22_bwjn_core_141;
  wire popcount22_bwjn_core_143;
  wire popcount22_bwjn_core_144;
  wire popcount22_bwjn_core_145;
  wire popcount22_bwjn_core_146;
  wire popcount22_bwjn_core_149;
  wire popcount22_bwjn_core_150;
  wire popcount22_bwjn_core_155;
  wire popcount22_bwjn_core_158;
  wire popcount22_bwjn_core_160;
  wire popcount22_bwjn_core_161;

  assign popcount22_bwjn_core_027 = ~(input_a[15] | input_a[5]);
  assign popcount22_bwjn_core_028 = input_a[1] ^ input_a[17];
  assign popcount22_bwjn_core_030 = input_a[17] & input_a[2];
  assign popcount22_bwjn_core_031 = ~(input_a[12] & input_a[5]);
  assign popcount22_bwjn_core_033 = input_a[0] | input_a[15];
  assign popcount22_bwjn_core_034 = input_a[13] ^ input_a[1];
  assign popcount22_bwjn_core_038 = ~input_a[6];
  assign popcount22_bwjn_core_039 = input_a[14] | input_a[16];
  assign popcount22_bwjn_core_040 = ~(input_a[7] & input_a[10]);
  assign popcount22_bwjn_core_042_not = ~input_a[15];
  assign popcount22_bwjn_core_043 = ~(input_a[15] | input_a[3]);
  assign popcount22_bwjn_core_044 = input_a[9] ^ input_a[21];
  assign popcount22_bwjn_core_046 = ~input_a[1];
  assign popcount22_bwjn_core_048 = input_a[6] ^ input_a[3];
  assign popcount22_bwjn_core_051_not = ~input_a[7];
  assign popcount22_bwjn_core_053 = input_a[4] | input_a[4];
  assign popcount22_bwjn_core_055 = ~input_a[9];
  assign popcount22_bwjn_core_056 = ~(input_a[6] ^ input_a[5]);
  assign popcount22_bwjn_core_057 = input_a[14] & input_a[19];
  assign popcount22_bwjn_core_058 = input_a[5] & input_a[15];
  assign popcount22_bwjn_core_059 = ~input_a[17];
  assign popcount22_bwjn_core_060 = input_a[12] ^ input_a[17];
  assign popcount22_bwjn_core_062 = input_a[14] ^ input_a[9];
  assign popcount22_bwjn_core_063 = ~(input_a[10] | input_a[13]);
  assign popcount22_bwjn_core_064_not = ~input_a[11];
  assign popcount22_bwjn_core_065_not = ~input_a[12];
  assign popcount22_bwjn_core_067 = ~(input_a[15] | input_a[0]);
  assign popcount22_bwjn_core_070 = ~(input_a[4] & input_a[12]);
  assign popcount22_bwjn_core_072 = input_a[7] & input_a[15];
  assign popcount22_bwjn_core_074 = ~(input_a[13] | input_a[21]);
  assign popcount22_bwjn_core_077 = input_a[9] & input_a[13];
  assign popcount22_bwjn_core_078 = input_a[4] & input_a[11];
  assign popcount22_bwjn_core_079 = input_a[6] & input_a[5];
  assign popcount22_bwjn_core_080 = input_a[4] ^ input_a[13];
  assign popcount22_bwjn_core_081_not = ~input_a[1];
  assign popcount22_bwjn_core_083 = input_a[15] & input_a[4];
  assign popcount22_bwjn_core_086 = input_a[13] & input_a[6];
  assign popcount22_bwjn_core_088_not = ~input_a[15];
  assign popcount22_bwjn_core_090 = input_a[0] ^ input_a[0];
  assign popcount22_bwjn_core_091 = input_a[10] ^ input_a[21];
  assign popcount22_bwjn_core_093 = ~(input_a[7] | input_a[14]);
  assign popcount22_bwjn_core_094 = ~(input_a[8] & input_a[11]);
  assign popcount22_bwjn_core_099 = ~(input_a[21] | input_a[4]);
  assign popcount22_bwjn_core_102 = ~input_a[4];
  assign popcount22_bwjn_core_103 = input_a[19] | input_a[21];
  assign popcount22_bwjn_core_105 = ~(input_a[0] & input_a[15]);
  assign popcount22_bwjn_core_106 = ~input_a[16];
  assign popcount22_bwjn_core_107 = input_a[7] ^ input_a[13];
  assign popcount22_bwjn_core_112 = ~(input_a[1] ^ input_a[8]);
  assign popcount22_bwjn_core_113 = input_a[15] ^ input_a[10];
  assign popcount22_bwjn_core_116 = ~(input_a[5] & input_a[17]);
  assign popcount22_bwjn_core_117 = ~(input_a[6] ^ input_a[8]);
  assign popcount22_bwjn_core_121 = ~(input_a[7] | input_a[4]);
  assign popcount22_bwjn_core_122 = ~input_a[18];
  assign popcount22_bwjn_core_124 = ~(input_a[14] ^ input_a[1]);
  assign popcount22_bwjn_core_125 = ~(input_a[9] & input_a[4]);
  assign popcount22_bwjn_core_127 = input_a[19] ^ input_a[17];
  assign popcount22_bwjn_core_129 = ~(input_a[18] & input_a[20]);
  assign popcount22_bwjn_core_133 = ~(input_a[12] & input_a[20]);
  assign popcount22_bwjn_core_134 = ~input_a[0];
  assign popcount22_bwjn_core_136 = ~(input_a[5] & input_a[5]);
  assign popcount22_bwjn_core_137 = input_a[14] ^ input_a[5];
  assign popcount22_bwjn_core_139 = ~input_a[5];
  assign popcount22_bwjn_core_141 = ~(input_a[9] & input_a[15]);
  assign popcount22_bwjn_core_143 = ~(input_a[10] & input_a[19]);
  assign popcount22_bwjn_core_144 = input_a[11] | input_a[18];
  assign popcount22_bwjn_core_145 = ~(input_a[16] ^ input_a[17]);
  assign popcount22_bwjn_core_146 = input_a[21] | input_a[15];
  assign popcount22_bwjn_core_149 = ~(input_a[9] | input_a[9]);
  assign popcount22_bwjn_core_150 = input_a[7] | input_a[5];
  assign popcount22_bwjn_core_155 = ~(input_a[18] | input_a[9]);
  assign popcount22_bwjn_core_158 = ~(input_a[6] ^ input_a[11]);
  assign popcount22_bwjn_core_160 = ~(input_a[9] ^ input_a[10]);
  assign popcount22_bwjn_core_161 = input_a[20] ^ input_a[1];

  assign popcount22_bwjn_out[0] = 1'b1;
  assign popcount22_bwjn_out[1] = input_a[0];
  assign popcount22_bwjn_out[2] = 1'b1;
  assign popcount22_bwjn_out[3] = input_a[14];
  assign popcount22_bwjn_out[4] = 1'b0;
endmodule