// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.61389
// WCE=14.0
// EP=0.944553%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_n0hk(input [21:0] input_a, output [4:0] popcount22_n0hk_out);
  wire popcount22_n0hk_core_024_not;
  wire popcount22_n0hk_core_026;
  wire popcount22_n0hk_core_027;
  wire popcount22_n0hk_core_028;
  wire popcount22_n0hk_core_031;
  wire popcount22_n0hk_core_032;
  wire popcount22_n0hk_core_033;
  wire popcount22_n0hk_core_034;
  wire popcount22_n0hk_core_035;
  wire popcount22_n0hk_core_036;
  wire popcount22_n0hk_core_037;
  wire popcount22_n0hk_core_038;
  wire popcount22_n0hk_core_042;
  wire popcount22_n0hk_core_044;
  wire popcount22_n0hk_core_045;
  wire popcount22_n0hk_core_046;
  wire popcount22_n0hk_core_051_not;
  wire popcount22_n0hk_core_053;
  wire popcount22_n0hk_core_054;
  wire popcount22_n0hk_core_055;
  wire popcount22_n0hk_core_057;
  wire popcount22_n0hk_core_062;
  wire popcount22_n0hk_core_063;
  wire popcount22_n0hk_core_065;
  wire popcount22_n0hk_core_067;
  wire popcount22_n0hk_core_068;
  wire popcount22_n0hk_core_069;
  wire popcount22_n0hk_core_070;
  wire popcount22_n0hk_core_071;
  wire popcount22_n0hk_core_074;
  wire popcount22_n0hk_core_076;
  wire popcount22_n0hk_core_077;
  wire popcount22_n0hk_core_078;
  wire popcount22_n0hk_core_079;
  wire popcount22_n0hk_core_080;
  wire popcount22_n0hk_core_081;
  wire popcount22_n0hk_core_082;
  wire popcount22_n0hk_core_083;
  wire popcount22_n0hk_core_084;
  wire popcount22_n0hk_core_085;
  wire popcount22_n0hk_core_086;
  wire popcount22_n0hk_core_088;
  wire popcount22_n0hk_core_089;
  wire popcount22_n0hk_core_091;
  wire popcount22_n0hk_core_093;
  wire popcount22_n0hk_core_094;
  wire popcount22_n0hk_core_095;
  wire popcount22_n0hk_core_096;
  wire popcount22_n0hk_core_097;
  wire popcount22_n0hk_core_099_not;
  wire popcount22_n0hk_core_103;
  wire popcount22_n0hk_core_105;
  wire popcount22_n0hk_core_106;
  wire popcount22_n0hk_core_107;
  wire popcount22_n0hk_core_108;
  wire popcount22_n0hk_core_109;
  wire popcount22_n0hk_core_110;
  wire popcount22_n0hk_core_111;
  wire popcount22_n0hk_core_113;
  wire popcount22_n0hk_core_114;
  wire popcount22_n0hk_core_118;
  wire popcount22_n0hk_core_120;
  wire popcount22_n0hk_core_125;
  wire popcount22_n0hk_core_126;
  wire popcount22_n0hk_core_130;
  wire popcount22_n0hk_core_131;
  wire popcount22_n0hk_core_132;
  wire popcount22_n0hk_core_133;
  wire popcount22_n0hk_core_134;
  wire popcount22_n0hk_core_135;
  wire popcount22_n0hk_core_136;
  wire popcount22_n0hk_core_138;
  wire popcount22_n0hk_core_141;
  wire popcount22_n0hk_core_146;
  wire popcount22_n0hk_core_147;
  wire popcount22_n0hk_core_149;
  wire popcount22_n0hk_core_150;
  wire popcount22_n0hk_core_152;
  wire popcount22_n0hk_core_153_not;
  wire popcount22_n0hk_core_156;
  wire popcount22_n0hk_core_158;
  wire popcount22_n0hk_core_159;
  wire popcount22_n0hk_core_160_not;

  assign popcount22_n0hk_core_024_not = ~input_a[17];
  assign popcount22_n0hk_core_026 = input_a[10] & input_a[5];
  assign popcount22_n0hk_core_027 = ~(input_a[18] | input_a[3]);
  assign popcount22_n0hk_core_028 = ~(input_a[21] ^ input_a[16]);
  assign popcount22_n0hk_core_031 = input_a[0] ^ input_a[5];
  assign popcount22_n0hk_core_032 = input_a[17] ^ input_a[13];
  assign popcount22_n0hk_core_033 = ~(input_a[18] ^ input_a[17]);
  assign popcount22_n0hk_core_034 = input_a[11] | input_a[17];
  assign popcount22_n0hk_core_035 = input_a[5] | input_a[1];
  assign popcount22_n0hk_core_036 = input_a[19] & input_a[14];
  assign popcount22_n0hk_core_037 = ~(input_a[13] & input_a[2]);
  assign popcount22_n0hk_core_038 = ~(input_a[14] ^ input_a[20]);
  assign popcount22_n0hk_core_042 = ~(input_a[15] ^ input_a[11]);
  assign popcount22_n0hk_core_044 = input_a[14] ^ input_a[7];
  assign popcount22_n0hk_core_045 = ~input_a[21];
  assign popcount22_n0hk_core_046 = input_a[13] & input_a[21];
  assign popcount22_n0hk_core_051_not = ~input_a[14];
  assign popcount22_n0hk_core_053 = input_a[10] & input_a[17];
  assign popcount22_n0hk_core_054 = input_a[17] | input_a[1];
  assign popcount22_n0hk_core_055 = ~(input_a[10] ^ input_a[17]);
  assign popcount22_n0hk_core_057 = ~(input_a[7] & input_a[13]);
  assign popcount22_n0hk_core_062 = input_a[2] | input_a[12];
  assign popcount22_n0hk_core_063 = ~(input_a[15] & input_a[7]);
  assign popcount22_n0hk_core_065 = ~(input_a[4] & input_a[17]);
  assign popcount22_n0hk_core_067 = input_a[21] & input_a[3];
  assign popcount22_n0hk_core_068 = input_a[20] | input_a[8];
  assign popcount22_n0hk_core_069 = ~(input_a[19] & input_a[7]);
  assign popcount22_n0hk_core_070 = ~(input_a[4] | input_a[16]);
  assign popcount22_n0hk_core_071 = input_a[2] & input_a[17];
  assign popcount22_n0hk_core_074 = input_a[14] | input_a[19];
  assign popcount22_n0hk_core_076 = ~(input_a[19] | input_a[8]);
  assign popcount22_n0hk_core_077 = ~input_a[14];
  assign popcount22_n0hk_core_078 = input_a[1] | input_a[7];
  assign popcount22_n0hk_core_079 = ~(input_a[2] | input_a[7]);
  assign popcount22_n0hk_core_080 = ~(input_a[0] | input_a[8]);
  assign popcount22_n0hk_core_081 = ~(input_a[2] & input_a[21]);
  assign popcount22_n0hk_core_082 = ~input_a[15];
  assign popcount22_n0hk_core_083 = input_a[10] ^ input_a[19];
  assign popcount22_n0hk_core_084 = ~(input_a[13] ^ input_a[19]);
  assign popcount22_n0hk_core_085 = input_a[18] ^ input_a[4];
  assign popcount22_n0hk_core_086 = input_a[4] ^ input_a[8];
  assign popcount22_n0hk_core_088 = input_a[20] | input_a[13];
  assign popcount22_n0hk_core_089 = ~(input_a[7] ^ input_a[6]);
  assign popcount22_n0hk_core_091 = ~(input_a[14] & input_a[6]);
  assign popcount22_n0hk_core_093 = input_a[8] & input_a[0];
  assign popcount22_n0hk_core_094 = input_a[21] & input_a[2];
  assign popcount22_n0hk_core_095 = input_a[21] | input_a[0];
  assign popcount22_n0hk_core_096 = ~(input_a[8] & input_a[9]);
  assign popcount22_n0hk_core_097 = ~input_a[13];
  assign popcount22_n0hk_core_099_not = ~input_a[7];
  assign popcount22_n0hk_core_103 = input_a[21] | input_a[21];
  assign popcount22_n0hk_core_105 = input_a[8] ^ input_a[7];
  assign popcount22_n0hk_core_106 = input_a[16] & input_a[19];
  assign popcount22_n0hk_core_107 = ~(input_a[10] | input_a[18]);
  assign popcount22_n0hk_core_108 = ~(input_a[12] & input_a[15]);
  assign popcount22_n0hk_core_109 = input_a[11] | input_a[17];
  assign popcount22_n0hk_core_110 = ~(input_a[18] & input_a[0]);
  assign popcount22_n0hk_core_111 = input_a[21] ^ input_a[20];
  assign popcount22_n0hk_core_113 = input_a[1] & input_a[20];
  assign popcount22_n0hk_core_114 = ~(input_a[9] | input_a[2]);
  assign popcount22_n0hk_core_118 = input_a[10] | input_a[18];
  assign popcount22_n0hk_core_120 = ~(input_a[18] | input_a[0]);
  assign popcount22_n0hk_core_125 = input_a[17] | input_a[6];
  assign popcount22_n0hk_core_126 = ~(input_a[17] | input_a[18]);
  assign popcount22_n0hk_core_130 = input_a[9] ^ input_a[17];
  assign popcount22_n0hk_core_131 = input_a[1] | input_a[18];
  assign popcount22_n0hk_core_132 = input_a[10] | input_a[16];
  assign popcount22_n0hk_core_133 = ~(input_a[20] & input_a[21]);
  assign popcount22_n0hk_core_134 = input_a[12] ^ input_a[10];
  assign popcount22_n0hk_core_135 = ~(input_a[6] ^ input_a[15]);
  assign popcount22_n0hk_core_136 = ~(input_a[11] | input_a[6]);
  assign popcount22_n0hk_core_138 = ~(input_a[13] & input_a[5]);
  assign popcount22_n0hk_core_141 = input_a[15] & input_a[9];
  assign popcount22_n0hk_core_146 = ~(input_a[10] ^ input_a[19]);
  assign popcount22_n0hk_core_147 = ~(input_a[7] ^ input_a[13]);
  assign popcount22_n0hk_core_149 = ~(input_a[14] | input_a[8]);
  assign popcount22_n0hk_core_150 = ~(input_a[12] | input_a[7]);
  assign popcount22_n0hk_core_152 = input_a[3] ^ input_a[11];
  assign popcount22_n0hk_core_153_not = ~input_a[19];
  assign popcount22_n0hk_core_156 = ~(input_a[21] & input_a[13]);
  assign popcount22_n0hk_core_158 = input_a[10] & input_a[19];
  assign popcount22_n0hk_core_159 = input_a[17] ^ input_a[19];
  assign popcount22_n0hk_core_160_not = ~input_a[18];

  assign popcount22_n0hk_out[0] = input_a[6];
  assign popcount22_n0hk_out[1] = 1'b1;
  assign popcount22_n0hk_out[2] = 1'b1;
  assign popcount22_n0hk_out[3] = input_a[10];
  assign popcount22_n0hk_out[4] = 1'b0;
endmodule