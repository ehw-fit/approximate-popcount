// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.09399
// WCE=19.0
// EP=0.904678%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_zx80(input [33:0] input_a, output [5:0] popcount34_zx80_out);
  wire popcount34_zx80_core_037;
  wire popcount34_zx80_core_038;
  wire popcount34_zx80_core_039;
  wire popcount34_zx80_core_040;
  wire popcount34_zx80_core_043;
  wire popcount34_zx80_core_044;
  wire popcount34_zx80_core_048;
  wire popcount34_zx80_core_049;
  wire popcount34_zx80_core_050;
  wire popcount34_zx80_core_051;
  wire popcount34_zx80_core_054;
  wire popcount34_zx80_core_059;
  wire popcount34_zx80_core_060;
  wire popcount34_zx80_core_061;
  wire popcount34_zx80_core_062;
  wire popcount34_zx80_core_063;
  wire popcount34_zx80_core_065;
  wire popcount34_zx80_core_066;
  wire popcount34_zx80_core_067_not;
  wire popcount34_zx80_core_069;
  wire popcount34_zx80_core_073;
  wire popcount34_zx80_core_075;
  wire popcount34_zx80_core_077;
  wire popcount34_zx80_core_081;
  wire popcount34_zx80_core_082;
  wire popcount34_zx80_core_084;
  wire popcount34_zx80_core_085;
  wire popcount34_zx80_core_086;
  wire popcount34_zx80_core_087;
  wire popcount34_zx80_core_088;
  wire popcount34_zx80_core_091;
  wire popcount34_zx80_core_094;
  wire popcount34_zx80_core_095;
  wire popcount34_zx80_core_097;
  wire popcount34_zx80_core_098;
  wire popcount34_zx80_core_099;
  wire popcount34_zx80_core_100;
  wire popcount34_zx80_core_103;
  wire popcount34_zx80_core_106;
  wire popcount34_zx80_core_107;
  wire popcount34_zx80_core_108;
  wire popcount34_zx80_core_111;
  wire popcount34_zx80_core_112;
  wire popcount34_zx80_core_113;
  wire popcount34_zx80_core_114;
  wire popcount34_zx80_core_115;
  wire popcount34_zx80_core_117;
  wire popcount34_zx80_core_118;
  wire popcount34_zx80_core_120;
  wire popcount34_zx80_core_122;
  wire popcount34_zx80_core_125;
  wire popcount34_zx80_core_126;
  wire popcount34_zx80_core_131;
  wire popcount34_zx80_core_133;
  wire popcount34_zx80_core_136;
  wire popcount34_zx80_core_137;
  wire popcount34_zx80_core_138;
  wire popcount34_zx80_core_140;
  wire popcount34_zx80_core_145;
  wire popcount34_zx80_core_146;
  wire popcount34_zx80_core_147;
  wire popcount34_zx80_core_148;
  wire popcount34_zx80_core_149;
  wire popcount34_zx80_core_150;
  wire popcount34_zx80_core_151;
  wire popcount34_zx80_core_152;
  wire popcount34_zx80_core_154;
  wire popcount34_zx80_core_155;
  wire popcount34_zx80_core_156_not;
  wire popcount34_zx80_core_158;
  wire popcount34_zx80_core_159;
  wire popcount34_zx80_core_160;
  wire popcount34_zx80_core_162;
  wire popcount34_zx80_core_163;
  wire popcount34_zx80_core_164;
  wire popcount34_zx80_core_165;
  wire popcount34_zx80_core_166;
  wire popcount34_zx80_core_167;
  wire popcount34_zx80_core_168;
  wire popcount34_zx80_core_172;
  wire popcount34_zx80_core_174;
  wire popcount34_zx80_core_176;
  wire popcount34_zx80_core_177;
  wire popcount34_zx80_core_178;
  wire popcount34_zx80_core_180;
  wire popcount34_zx80_core_181;
  wire popcount34_zx80_core_182;
  wire popcount34_zx80_core_183;
  wire popcount34_zx80_core_185_not;
  wire popcount34_zx80_core_186;
  wire popcount34_zx80_core_188;
  wire popcount34_zx80_core_189;
  wire popcount34_zx80_core_191;
  wire popcount34_zx80_core_192;
  wire popcount34_zx80_core_193;
  wire popcount34_zx80_core_194;
  wire popcount34_zx80_core_195;
  wire popcount34_zx80_core_196;
  wire popcount34_zx80_core_198;
  wire popcount34_zx80_core_199;
  wire popcount34_zx80_core_200;
  wire popcount34_zx80_core_203;
  wire popcount34_zx80_core_204;
  wire popcount34_zx80_core_206;
  wire popcount34_zx80_core_207;
  wire popcount34_zx80_core_208;
  wire popcount34_zx80_core_209;
  wire popcount34_zx80_core_210;
  wire popcount34_zx80_core_211;
  wire popcount34_zx80_core_212;
  wire popcount34_zx80_core_213;
  wire popcount34_zx80_core_214;
  wire popcount34_zx80_core_216;
  wire popcount34_zx80_core_218;
  wire popcount34_zx80_core_220;
  wire popcount34_zx80_core_221;
  wire popcount34_zx80_core_222;
  wire popcount34_zx80_core_225;
  wire popcount34_zx80_core_226;
  wire popcount34_zx80_core_229;
  wire popcount34_zx80_core_230;
  wire popcount34_zx80_core_233;
  wire popcount34_zx80_core_234;
  wire popcount34_zx80_core_237;
  wire popcount34_zx80_core_239;
  wire popcount34_zx80_core_240;
  wire popcount34_zx80_core_241;
  wire popcount34_zx80_core_242;
  wire popcount34_zx80_core_243;
  wire popcount34_zx80_core_244;
  wire popcount34_zx80_core_245;
  wire popcount34_zx80_core_248;
  wire popcount34_zx80_core_250;
  wire popcount34_zx80_core_251;
  wire popcount34_zx80_core_252;

  assign popcount34_zx80_core_037 = ~(input_a[21] & input_a[9]);
  assign popcount34_zx80_core_038 = input_a[6] ^ input_a[1];
  assign popcount34_zx80_core_039 = input_a[15] | input_a[31];
  assign popcount34_zx80_core_040 = ~(input_a[28] | input_a[23]);
  assign popcount34_zx80_core_043 = input_a[27] | input_a[4];
  assign popcount34_zx80_core_044 = ~(input_a[20] | input_a[2]);
  assign popcount34_zx80_core_048 = input_a[24] & input_a[0];
  assign popcount34_zx80_core_049 = input_a[29] ^ input_a[30];
  assign popcount34_zx80_core_050 = ~(input_a[24] | input_a[9]);
  assign popcount34_zx80_core_051 = ~(input_a[26] ^ input_a[19]);
  assign popcount34_zx80_core_054 = ~(input_a[30] & input_a[19]);
  assign popcount34_zx80_core_059 = ~(input_a[23] & input_a[3]);
  assign popcount34_zx80_core_060 = ~(input_a[21] & input_a[8]);
  assign popcount34_zx80_core_061 = ~(input_a[2] | input_a[5]);
  assign popcount34_zx80_core_062 = ~(input_a[11] ^ input_a[5]);
  assign popcount34_zx80_core_063 = input_a[21] | input_a[16];
  assign popcount34_zx80_core_065 = input_a[8] & input_a[6];
  assign popcount34_zx80_core_066 = input_a[15] ^ input_a[30];
  assign popcount34_zx80_core_067_not = ~input_a[7];
  assign popcount34_zx80_core_069 = ~(input_a[17] & input_a[18]);
  assign popcount34_zx80_core_073 = ~(input_a[15] & input_a[28]);
  assign popcount34_zx80_core_075 = ~input_a[7];
  assign popcount34_zx80_core_077 = input_a[15] ^ input_a[8];
  assign popcount34_zx80_core_081 = ~(input_a[24] & input_a[30]);
  assign popcount34_zx80_core_082 = input_a[3] & input_a[33];
  assign popcount34_zx80_core_084 = input_a[19] | input_a[7];
  assign popcount34_zx80_core_085 = ~(input_a[26] & input_a[2]);
  assign popcount34_zx80_core_086 = ~(input_a[21] ^ input_a[0]);
  assign popcount34_zx80_core_087 = ~(input_a[27] ^ input_a[33]);
  assign popcount34_zx80_core_088 = input_a[16] | input_a[23];
  assign popcount34_zx80_core_091 = input_a[8] ^ input_a[33];
  assign popcount34_zx80_core_094 = input_a[21] ^ input_a[14];
  assign popcount34_zx80_core_095 = ~(input_a[15] & input_a[20]);
  assign popcount34_zx80_core_097 = input_a[11] & input_a[4];
  assign popcount34_zx80_core_098 = ~(input_a[5] ^ input_a[14]);
  assign popcount34_zx80_core_099 = input_a[4] ^ input_a[22];
  assign popcount34_zx80_core_100 = input_a[10] ^ input_a[4];
  assign popcount34_zx80_core_103 = ~input_a[30];
  assign popcount34_zx80_core_106 = input_a[30] ^ input_a[6];
  assign popcount34_zx80_core_107 = ~input_a[1];
  assign popcount34_zx80_core_108 = ~(input_a[31] & input_a[19]);
  assign popcount34_zx80_core_111 = ~(input_a[22] ^ input_a[19]);
  assign popcount34_zx80_core_112 = input_a[10] & input_a[27];
  assign popcount34_zx80_core_113 = ~input_a[10];
  assign popcount34_zx80_core_114 = ~(input_a[2] ^ input_a[17]);
  assign popcount34_zx80_core_115 = ~(input_a[25] ^ input_a[10]);
  assign popcount34_zx80_core_117 = ~input_a[19];
  assign popcount34_zx80_core_118 = input_a[24] & input_a[28];
  assign popcount34_zx80_core_120 = input_a[10] & input_a[27];
  assign popcount34_zx80_core_122 = ~input_a[17];
  assign popcount34_zx80_core_125 = input_a[7] | input_a[14];
  assign popcount34_zx80_core_126 = ~(input_a[2] & input_a[20]);
  assign popcount34_zx80_core_131 = ~input_a[1];
  assign popcount34_zx80_core_133 = ~(input_a[9] ^ input_a[3]);
  assign popcount34_zx80_core_136 = ~(input_a[29] ^ input_a[15]);
  assign popcount34_zx80_core_137 = ~(input_a[28] & input_a[18]);
  assign popcount34_zx80_core_138 = ~(input_a[27] & input_a[5]);
  assign popcount34_zx80_core_140 = input_a[22] & input_a[30];
  assign popcount34_zx80_core_145 = ~(input_a[29] | input_a[25]);
  assign popcount34_zx80_core_146 = ~(input_a[26] & input_a[19]);
  assign popcount34_zx80_core_147 = ~(input_a[8] & input_a[0]);
  assign popcount34_zx80_core_148 = ~(input_a[10] ^ input_a[24]);
  assign popcount34_zx80_core_149 = ~input_a[0];
  assign popcount34_zx80_core_150 = input_a[18] ^ input_a[5];
  assign popcount34_zx80_core_151 = ~(input_a[28] | input_a[29]);
  assign popcount34_zx80_core_152 = input_a[18] | input_a[6];
  assign popcount34_zx80_core_154 = input_a[33] & input_a[3];
  assign popcount34_zx80_core_155 = input_a[1] | input_a[27];
  assign popcount34_zx80_core_156_not = ~input_a[13];
  assign popcount34_zx80_core_158 = input_a[15] | input_a[18];
  assign popcount34_zx80_core_159 = ~(input_a[11] & input_a[20]);
  assign popcount34_zx80_core_160 = ~input_a[32];
  assign popcount34_zx80_core_162 = input_a[29] & input_a[33];
  assign popcount34_zx80_core_163 = ~(input_a[4] | input_a[21]);
  assign popcount34_zx80_core_164 = ~(input_a[3] | input_a[6]);
  assign popcount34_zx80_core_165 = ~(input_a[27] ^ input_a[9]);
  assign popcount34_zx80_core_166 = ~(input_a[22] & input_a[11]);
  assign popcount34_zx80_core_167 = ~input_a[12];
  assign popcount34_zx80_core_168 = ~(input_a[0] | input_a[29]);
  assign popcount34_zx80_core_172 = ~(input_a[25] ^ input_a[9]);
  assign popcount34_zx80_core_174 = ~input_a[14];
  assign popcount34_zx80_core_176 = ~(input_a[22] ^ input_a[10]);
  assign popcount34_zx80_core_177 = input_a[6] ^ input_a[4];
  assign popcount34_zx80_core_178 = ~(input_a[3] | input_a[9]);
  assign popcount34_zx80_core_180 = ~(input_a[29] | input_a[25]);
  assign popcount34_zx80_core_181 = input_a[31] & input_a[3];
  assign popcount34_zx80_core_182 = ~(input_a[12] ^ input_a[23]);
  assign popcount34_zx80_core_183 = ~(input_a[30] | input_a[17]);
  assign popcount34_zx80_core_185_not = ~input_a[30];
  assign popcount34_zx80_core_186 = ~(input_a[33] ^ input_a[33]);
  assign popcount34_zx80_core_188 = ~(input_a[8] | input_a[20]);
  assign popcount34_zx80_core_189 = ~input_a[15];
  assign popcount34_zx80_core_191 = ~(input_a[10] | input_a[29]);
  assign popcount34_zx80_core_192 = input_a[19] ^ input_a[25];
  assign popcount34_zx80_core_193 = input_a[26] | input_a[33];
  assign popcount34_zx80_core_194 = input_a[32] ^ input_a[2];
  assign popcount34_zx80_core_195 = input_a[5] | input_a[8];
  assign popcount34_zx80_core_196 = input_a[20] | input_a[5];
  assign popcount34_zx80_core_198 = ~input_a[10];
  assign popcount34_zx80_core_199 = input_a[9] & input_a[2];
  assign popcount34_zx80_core_200 = ~(input_a[18] ^ input_a[17]);
  assign popcount34_zx80_core_203 = ~(input_a[7] | input_a[12]);
  assign popcount34_zx80_core_204 = ~(input_a[15] | input_a[25]);
  assign popcount34_zx80_core_206 = input_a[25] | input_a[30];
  assign popcount34_zx80_core_207 = ~(input_a[13] ^ input_a[33]);
  assign popcount34_zx80_core_208 = ~input_a[7];
  assign popcount34_zx80_core_209 = input_a[7] & input_a[15];
  assign popcount34_zx80_core_210 = input_a[19] & input_a[27];
  assign popcount34_zx80_core_211 = input_a[30] & input_a[7];
  assign popcount34_zx80_core_212 = ~(input_a[28] & input_a[21]);
  assign popcount34_zx80_core_213 = ~(input_a[5] & input_a[12]);
  assign popcount34_zx80_core_214 = ~(input_a[13] ^ input_a[1]);
  assign popcount34_zx80_core_216 = input_a[30] & input_a[18];
  assign popcount34_zx80_core_218 = input_a[29] & input_a[12];
  assign popcount34_zx80_core_220 = ~input_a[5];
  assign popcount34_zx80_core_221 = ~(input_a[33] | input_a[3]);
  assign popcount34_zx80_core_222 = input_a[16] | input_a[15];
  assign popcount34_zx80_core_225 = ~(input_a[27] | input_a[19]);
  assign popcount34_zx80_core_226 = input_a[23] | input_a[18];
  assign popcount34_zx80_core_229 = input_a[3] ^ input_a[18];
  assign popcount34_zx80_core_230 = input_a[16] | input_a[11];
  assign popcount34_zx80_core_233 = input_a[13] ^ input_a[25];
  assign popcount34_zx80_core_234 = ~(input_a[8] | input_a[32]);
  assign popcount34_zx80_core_237 = ~(input_a[14] & input_a[18]);
  assign popcount34_zx80_core_239 = ~(input_a[26] ^ input_a[11]);
  assign popcount34_zx80_core_240 = ~(input_a[31] | input_a[22]);
  assign popcount34_zx80_core_241 = input_a[29] ^ input_a[28];
  assign popcount34_zx80_core_242 = ~(input_a[1] ^ input_a[13]);
  assign popcount34_zx80_core_243 = input_a[31] & input_a[22];
  assign popcount34_zx80_core_244 = ~input_a[4];
  assign popcount34_zx80_core_245 = ~(input_a[3] & input_a[27]);
  assign popcount34_zx80_core_248 = ~(input_a[19] & input_a[20]);
  assign popcount34_zx80_core_250 = ~(input_a[25] | input_a[1]);
  assign popcount34_zx80_core_251 = input_a[2] ^ input_a[10];
  assign popcount34_zx80_core_252 = input_a[2] & input_a[23];

  assign popcount34_zx80_out[0] = input_a[20];
  assign popcount34_zx80_out[1] = 1'b1;
  assign popcount34_zx80_out[2] = 1'b1;
  assign popcount34_zx80_out[3] = 1'b1;
  assign popcount34_zx80_out[4] = 1'b0;
  assign popcount34_zx80_out[5] = 1'b0;
endmodule