// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.79152
// WCE=17.0
// EP=0.822902%
// Printed PDK parameters:
//  Area=55606870.0
//  Delay=82154984.0
//  Power=2605600.0

module popcount36_qqdr(input [35:0] input_a, output [5:0] popcount36_qqdr_out);
  wire popcount36_qqdr_core_038;
  wire popcount36_qqdr_core_039;
  wire popcount36_qqdr_core_041;
  wire popcount36_qqdr_core_042;
  wire popcount36_qqdr_core_043;
  wire popcount36_qqdr_core_044;
  wire popcount36_qqdr_core_045;
  wire popcount36_qqdr_core_050;
  wire popcount36_qqdr_core_051;
  wire popcount36_qqdr_core_052;
  wire popcount36_qqdr_core_053;
  wire popcount36_qqdr_core_054;
  wire popcount36_qqdr_core_055;
  wire popcount36_qqdr_core_057;
  wire popcount36_qqdr_core_058;
  wire popcount36_qqdr_core_059;
  wire popcount36_qqdr_core_066;
  wire popcount36_qqdr_core_067;
  wire popcount36_qqdr_core_068;
  wire popcount36_qqdr_core_069;
  wire popcount36_qqdr_core_070;
  wire popcount36_qqdr_core_071;
  wire popcount36_qqdr_core_072;
  wire popcount36_qqdr_core_073;
  wire popcount36_qqdr_core_075;
  wire popcount36_qqdr_core_076;
  wire popcount36_qqdr_core_078;
  wire popcount36_qqdr_core_079;
  wire popcount36_qqdr_core_080;
  wire popcount36_qqdr_core_081;
  wire popcount36_qqdr_core_086;
  wire popcount36_qqdr_core_087;
  wire popcount36_qqdr_core_088;
  wire popcount36_qqdr_core_089;
  wire popcount36_qqdr_core_091;
  wire popcount36_qqdr_core_092;
  wire popcount36_qqdr_core_094;
  wire popcount36_qqdr_core_096;
  wire popcount36_qqdr_core_099;
  wire popcount36_qqdr_core_100;
  wire popcount36_qqdr_core_101;
  wire popcount36_qqdr_core_103;
  wire popcount36_qqdr_core_104;
  wire popcount36_qqdr_core_108;
  wire popcount36_qqdr_core_109;
  wire popcount36_qqdr_core_110;
  wire popcount36_qqdr_core_111;
  wire popcount36_qqdr_core_113;
  wire popcount36_qqdr_core_116;
  wire popcount36_qqdr_core_117;
  wire popcount36_qqdr_core_118;
  wire popcount36_qqdr_core_120;
  wire popcount36_qqdr_core_122;
  wire popcount36_qqdr_core_123;
  wire popcount36_qqdr_core_124;
  wire popcount36_qqdr_core_125;
  wire popcount36_qqdr_core_126;
  wire popcount36_qqdr_core_127;
  wire popcount36_qqdr_core_128;
  wire popcount36_qqdr_core_129;
  wire popcount36_qqdr_core_130;
  wire popcount36_qqdr_core_131;
  wire popcount36_qqdr_core_132;
  wire popcount36_qqdr_core_133;
  wire popcount36_qqdr_core_135;
  wire popcount36_qqdr_core_139;
  wire popcount36_qqdr_core_140;
  wire popcount36_qqdr_core_142;
  wire popcount36_qqdr_core_143;
  wire popcount36_qqdr_core_144;
  wire popcount36_qqdr_core_145;
  wire popcount36_qqdr_core_146;
  wire popcount36_qqdr_core_147;
  wire popcount36_qqdr_core_148;
  wire popcount36_qqdr_core_149;
  wire popcount36_qqdr_core_150;
  wire popcount36_qqdr_core_151;
  wire popcount36_qqdr_core_152;
  wire popcount36_qqdr_core_153;
  wire popcount36_qqdr_core_154;
  wire popcount36_qqdr_core_155;
  wire popcount36_qqdr_core_156;
  wire popcount36_qqdr_core_158;
  wire popcount36_qqdr_core_159_not;
  wire popcount36_qqdr_core_160_not;
  wire popcount36_qqdr_core_161;
  wire popcount36_qqdr_core_163;
  wire popcount36_qqdr_core_164;
  wire popcount36_qqdr_core_165;
  wire popcount36_qqdr_core_166;
  wire popcount36_qqdr_core_167;
  wire popcount36_qqdr_core_168;
  wire popcount36_qqdr_core_169;
  wire popcount36_qqdr_core_172;
  wire popcount36_qqdr_core_173;
  wire popcount36_qqdr_core_174;
  wire popcount36_qqdr_core_175;
  wire popcount36_qqdr_core_176;
  wire popcount36_qqdr_core_177;
  wire popcount36_qqdr_core_178;
  wire popcount36_qqdr_core_179;
  wire popcount36_qqdr_core_181;
  wire popcount36_qqdr_core_182;
  wire popcount36_qqdr_core_183;
  wire popcount36_qqdr_core_185;
  wire popcount36_qqdr_core_186;
  wire popcount36_qqdr_core_187;
  wire popcount36_qqdr_core_188;
  wire popcount36_qqdr_core_189;
  wire popcount36_qqdr_core_190;
  wire popcount36_qqdr_core_191;
  wire popcount36_qqdr_core_192;
  wire popcount36_qqdr_core_194;
  wire popcount36_qqdr_core_195;
  wire popcount36_qqdr_core_198;
  wire popcount36_qqdr_core_201;
  wire popcount36_qqdr_core_202;
  wire popcount36_qqdr_core_204;
  wire popcount36_qqdr_core_205;
  wire popcount36_qqdr_core_206;
  wire popcount36_qqdr_core_207;
  wire popcount36_qqdr_core_211;
  wire popcount36_qqdr_core_212;
  wire popcount36_qqdr_core_213;
  wire popcount36_qqdr_core_214;
  wire popcount36_qqdr_core_215;
  wire popcount36_qqdr_core_216;
  wire popcount36_qqdr_core_219;
  wire popcount36_qqdr_core_222;
  wire popcount36_qqdr_core_223;
  wire popcount36_qqdr_core_224;
  wire popcount36_qqdr_core_225;
  wire popcount36_qqdr_core_226;
  wire popcount36_qqdr_core_228;
  wire popcount36_qqdr_core_229;
  wire popcount36_qqdr_core_230;
  wire popcount36_qqdr_core_231;
  wire popcount36_qqdr_core_232;
  wire popcount36_qqdr_core_233;
  wire popcount36_qqdr_core_234;
  wire popcount36_qqdr_core_235;
  wire popcount36_qqdr_core_236;
  wire popcount36_qqdr_core_237;
  wire popcount36_qqdr_core_238;
  wire popcount36_qqdr_core_239;
  wire popcount36_qqdr_core_242;
  wire popcount36_qqdr_core_243;
  wire popcount36_qqdr_core_246;
  wire popcount36_qqdr_core_247;
  wire popcount36_qqdr_core_250;
  wire popcount36_qqdr_core_251;
  wire popcount36_qqdr_core_252;
  wire popcount36_qqdr_core_253;
  wire popcount36_qqdr_core_254;
  wire popcount36_qqdr_core_255;
  wire popcount36_qqdr_core_256;
  wire popcount36_qqdr_core_257;
  wire popcount36_qqdr_core_258;
  wire popcount36_qqdr_core_259;
  wire popcount36_qqdr_core_260;
  wire popcount36_qqdr_core_261;
  wire popcount36_qqdr_core_262;
  wire popcount36_qqdr_core_263;
  wire popcount36_qqdr_core_264;
  wire popcount36_qqdr_core_265;
  wire popcount36_qqdr_core_266;
  wire popcount36_qqdr_core_268;
  wire popcount36_qqdr_core_270;
  wire popcount36_qqdr_core_271;
  wire popcount36_qqdr_core_272;
  wire popcount36_qqdr_core_274;
  wire popcount36_qqdr_core_275;
  wire popcount36_qqdr_core_276;

  assign popcount36_qqdr_core_038 = input_a[9] | input_a[20];
  assign popcount36_qqdr_core_039 = ~(input_a[12] ^ input_a[5]);
  assign popcount36_qqdr_core_041 = ~(input_a[20] & input_a[12]);
  assign popcount36_qqdr_core_042 = input_a[12] ^ input_a[13];
  assign popcount36_qqdr_core_043 = ~(input_a[31] | input_a[13]);
  assign popcount36_qqdr_core_044 = ~(input_a[25] & input_a[24]);
  assign popcount36_qqdr_core_045 = ~(input_a[4] ^ input_a[27]);
  assign popcount36_qqdr_core_050 = input_a[13] & input_a[5];
  assign popcount36_qqdr_core_051 = ~(input_a[20] | input_a[13]);
  assign popcount36_qqdr_core_052 = input_a[7] | input_a[27];
  assign popcount36_qqdr_core_053 = input_a[27] | input_a[10];
  assign popcount36_qqdr_core_054 = ~input_a[35];
  assign popcount36_qqdr_core_055 = ~input_a[26];
  assign popcount36_qqdr_core_057 = ~(input_a[30] & input_a[8]);
  assign popcount36_qqdr_core_058 = ~(input_a[16] | input_a[3]);
  assign popcount36_qqdr_core_059 = ~popcount36_qqdr_core_050;
  assign popcount36_qqdr_core_066 = input_a[24] | input_a[22];
  assign popcount36_qqdr_core_067 = input_a[26] & input_a[17];
  assign popcount36_qqdr_core_068 = input_a[29] ^ popcount36_qqdr_core_059;
  assign popcount36_qqdr_core_069 = ~(input_a[26] | input_a[25]);
  assign popcount36_qqdr_core_070 = popcount36_qqdr_core_068 ^ popcount36_qqdr_core_067;
  assign popcount36_qqdr_core_071 = input_a[26] & input_a[17];
  assign popcount36_qqdr_core_072 = input_a[29] | popcount36_qqdr_core_071;
  assign popcount36_qqdr_core_073 = input_a[29] | popcount36_qqdr_core_050;
  assign popcount36_qqdr_core_075 = popcount36_qqdr_core_073 | popcount36_qqdr_core_072;
  assign popcount36_qqdr_core_076 = input_a[21] | input_a[10];
  assign popcount36_qqdr_core_078 = input_a[6] & input_a[28];
  assign popcount36_qqdr_core_079 = input_a[13] & input_a[9];
  assign popcount36_qqdr_core_080 = ~(input_a[12] ^ input_a[7]);
  assign popcount36_qqdr_core_081 = ~input_a[35];
  assign popcount36_qqdr_core_086 = input_a[25] | input_a[34];
  assign popcount36_qqdr_core_087 = ~(input_a[2] | input_a[10]);
  assign popcount36_qqdr_core_088 = popcount36_qqdr_core_086 | input_a[20];
  assign popcount36_qqdr_core_089 = ~(input_a[29] & input_a[5]);
  assign popcount36_qqdr_core_091 = ~(input_a[9] ^ input_a[23]);
  assign popcount36_qqdr_core_092 = input_a[18] & input_a[24];
  assign popcount36_qqdr_core_094 = input_a[16] & input_a[2];
  assign popcount36_qqdr_core_096 = ~(input_a[21] & input_a[13]);
  assign popcount36_qqdr_core_099 = ~(input_a[14] ^ input_a[23]);
  assign popcount36_qqdr_core_100 = input_a[12] & input_a[28];
  assign popcount36_qqdr_core_101 = popcount36_qqdr_core_092 | popcount36_qqdr_core_094;
  assign popcount36_qqdr_core_103 = popcount36_qqdr_core_101 ^ popcount36_qqdr_core_100;
  assign popcount36_qqdr_core_104 = popcount36_qqdr_core_101 & popcount36_qqdr_core_100;
  assign popcount36_qqdr_core_108 = ~input_a[9];
  assign popcount36_qqdr_core_109 = input_a[34] & input_a[31];
  assign popcount36_qqdr_core_110 = popcount36_qqdr_core_088 ^ popcount36_qqdr_core_103;
  assign popcount36_qqdr_core_111 = popcount36_qqdr_core_088 & popcount36_qqdr_core_103;
  assign popcount36_qqdr_core_113 = input_a[23] | input_a[27];
  assign popcount36_qqdr_core_116 = input_a[28] & input_a[4];
  assign popcount36_qqdr_core_117 = popcount36_qqdr_core_104 | popcount36_qqdr_core_111;
  assign popcount36_qqdr_core_118 = ~(input_a[15] ^ input_a[25]);
  assign popcount36_qqdr_core_120 = input_a[14] ^ input_a[33];
  assign popcount36_qqdr_core_122 = ~(input_a[32] ^ input_a[35]);
  assign popcount36_qqdr_core_123 = input_a[22] & input_a[12];
  assign popcount36_qqdr_core_124 = popcount36_qqdr_core_070 ^ popcount36_qqdr_core_110;
  assign popcount36_qqdr_core_125 = popcount36_qqdr_core_070 & popcount36_qqdr_core_110;
  assign popcount36_qqdr_core_126 = popcount36_qqdr_core_124 ^ input_a[31];
  assign popcount36_qqdr_core_127 = popcount36_qqdr_core_124 & input_a[31];
  assign popcount36_qqdr_core_128 = popcount36_qqdr_core_125 | popcount36_qqdr_core_127;
  assign popcount36_qqdr_core_129 = popcount36_qqdr_core_075 ^ popcount36_qqdr_core_117;
  assign popcount36_qqdr_core_130 = popcount36_qqdr_core_075 & popcount36_qqdr_core_117;
  assign popcount36_qqdr_core_131 = popcount36_qqdr_core_129 ^ popcount36_qqdr_core_128;
  assign popcount36_qqdr_core_132 = popcount36_qqdr_core_129 & popcount36_qqdr_core_128;
  assign popcount36_qqdr_core_133 = popcount36_qqdr_core_130 | popcount36_qqdr_core_132;
  assign popcount36_qqdr_core_135 = input_a[35] | input_a[6];
  assign popcount36_qqdr_core_139 = input_a[15] | input_a[34];
  assign popcount36_qqdr_core_140 = ~(input_a[27] & input_a[0]);
  assign popcount36_qqdr_core_142 = ~(input_a[4] ^ input_a[24]);
  assign popcount36_qqdr_core_143 = input_a[13] & input_a[19];
  assign popcount36_qqdr_core_144 = ~(input_a[9] & input_a[19]);
  assign popcount36_qqdr_core_145 = input_a[0] & input_a[11];
  assign popcount36_qqdr_core_146 = input_a[19] ^ input_a[27];
  assign popcount36_qqdr_core_147 = input_a[6] & input_a[35];
  assign popcount36_qqdr_core_148 = ~(input_a[34] | input_a[8]);
  assign popcount36_qqdr_core_149 = input_a[19] & input_a[14];
  assign popcount36_qqdr_core_150 = popcount36_qqdr_core_145 ^ popcount36_qqdr_core_147;
  assign popcount36_qqdr_core_151 = popcount36_qqdr_core_145 & popcount36_qqdr_core_147;
  assign popcount36_qqdr_core_152 = popcount36_qqdr_core_150 ^ popcount36_qqdr_core_149;
  assign popcount36_qqdr_core_153 = popcount36_qqdr_core_150 & popcount36_qqdr_core_149;
  assign popcount36_qqdr_core_154 = popcount36_qqdr_core_151 | popcount36_qqdr_core_153;
  assign popcount36_qqdr_core_155 = input_a[22] ^ input_a[23];
  assign popcount36_qqdr_core_156 = input_a[22] & input_a[23];
  assign popcount36_qqdr_core_158 = input_a[25] | input_a[14];
  assign popcount36_qqdr_core_159_not = ~input_a[28];
  assign popcount36_qqdr_core_160_not = ~input_a[25];
  assign popcount36_qqdr_core_161 = input_a[1] | input_a[10];
  assign popcount36_qqdr_core_163 = ~input_a[18];
  assign popcount36_qqdr_core_164 = popcount36_qqdr_core_155 & input_a[7];
  assign popcount36_qqdr_core_165 = popcount36_qqdr_core_156 ^ popcount36_qqdr_core_161;
  assign popcount36_qqdr_core_166 = popcount36_qqdr_core_156 & popcount36_qqdr_core_161;
  assign popcount36_qqdr_core_167 = popcount36_qqdr_core_165 ^ popcount36_qqdr_core_164;
  assign popcount36_qqdr_core_168 = popcount36_qqdr_core_165 & popcount36_qqdr_core_164;
  assign popcount36_qqdr_core_169 = popcount36_qqdr_core_166 | popcount36_qqdr_core_168;
  assign popcount36_qqdr_core_172 = input_a[29] | input_a[29];
  assign popcount36_qqdr_core_173 = input_a[20] | input_a[24];
  assign popcount36_qqdr_core_174 = popcount36_qqdr_core_152 ^ popcount36_qqdr_core_167;
  assign popcount36_qqdr_core_175 = popcount36_qqdr_core_152 & popcount36_qqdr_core_167;
  assign popcount36_qqdr_core_176 = popcount36_qqdr_core_174 ^ input_a[9];
  assign popcount36_qqdr_core_177 = popcount36_qqdr_core_174 & input_a[9];
  assign popcount36_qqdr_core_178 = popcount36_qqdr_core_175 | popcount36_qqdr_core_177;
  assign popcount36_qqdr_core_179 = popcount36_qqdr_core_154 ^ popcount36_qqdr_core_169;
  assign popcount36_qqdr_core_181 = popcount36_qqdr_core_179 ^ popcount36_qqdr_core_178;
  assign popcount36_qqdr_core_182 = popcount36_qqdr_core_179 & input_a[9];
  assign popcount36_qqdr_core_183 = popcount36_qqdr_core_154 | popcount36_qqdr_core_182;
  assign popcount36_qqdr_core_185 = ~input_a[29];
  assign popcount36_qqdr_core_186 = input_a[35] ^ input_a[8];
  assign popcount36_qqdr_core_187 = input_a[8] & input_a[21];
  assign popcount36_qqdr_core_188 = ~(input_a[26] | input_a[19]);
  assign popcount36_qqdr_core_189 = input_a[9] & input_a[30];
  assign popcount36_qqdr_core_190 = input_a[35] | input_a[27];
  assign popcount36_qqdr_core_191 = ~(input_a[24] ^ input_a[29]);
  assign popcount36_qqdr_core_192 = popcount36_qqdr_core_187 ^ popcount36_qqdr_core_189;
  assign popcount36_qqdr_core_194 = popcount36_qqdr_core_192 ^ input_a[30];
  assign popcount36_qqdr_core_195 = ~(input_a[23] & input_a[16]);
  assign popcount36_qqdr_core_198 = ~input_a[15];
  assign popcount36_qqdr_core_201 = input_a[28] | input_a[11];
  assign popcount36_qqdr_core_202 = ~(input_a[21] ^ input_a[8]);
  assign popcount36_qqdr_core_204 = input_a[35] ^ input_a[33];
  assign popcount36_qqdr_core_205 = ~(input_a[21] & input_a[30]);
  assign popcount36_qqdr_core_206 = input_a[13] & input_a[19];
  assign popcount36_qqdr_core_207 = input_a[31] | input_a[10];
  assign popcount36_qqdr_core_211 = ~(input_a[16] & input_a[6]);
  assign popcount36_qqdr_core_212 = ~(input_a[3] | input_a[35]);
  assign popcount36_qqdr_core_213 = ~input_a[0];
  assign popcount36_qqdr_core_214 = input_a[11] | input_a[13];
  assign popcount36_qqdr_core_215 = input_a[10] | input_a[14];
  assign popcount36_qqdr_core_216 = ~popcount36_qqdr_core_194;
  assign popcount36_qqdr_core_219 = input_a[23] ^ input_a[14];
  assign popcount36_qqdr_core_222 = ~(input_a[5] ^ input_a[12]);
  assign popcount36_qqdr_core_223 = popcount36_qqdr_core_187 | popcount36_qqdr_core_194;
  assign popcount36_qqdr_core_224 = ~(input_a[17] & input_a[27]);
  assign popcount36_qqdr_core_225 = input_a[20] ^ input_a[8];
  assign popcount36_qqdr_core_226 = ~(input_a[13] ^ input_a[33]);
  assign popcount36_qqdr_core_228 = ~(input_a[6] ^ input_a[28]);
  assign popcount36_qqdr_core_229 = input_a[3] & input_a[15];
  assign popcount36_qqdr_core_230 = popcount36_qqdr_core_176 ^ popcount36_qqdr_core_216;
  assign popcount36_qqdr_core_231 = popcount36_qqdr_core_176 & popcount36_qqdr_core_216;
  assign popcount36_qqdr_core_232 = popcount36_qqdr_core_230 ^ popcount36_qqdr_core_229;
  assign popcount36_qqdr_core_233 = popcount36_qqdr_core_230 & popcount36_qqdr_core_229;
  assign popcount36_qqdr_core_234 = popcount36_qqdr_core_231 | popcount36_qqdr_core_233;
  assign popcount36_qqdr_core_235 = popcount36_qqdr_core_181 ^ popcount36_qqdr_core_223;
  assign popcount36_qqdr_core_236 = popcount36_qqdr_core_181 & popcount36_qqdr_core_223;
  assign popcount36_qqdr_core_237 = popcount36_qqdr_core_235 ^ popcount36_qqdr_core_234;
  assign popcount36_qqdr_core_238 = popcount36_qqdr_core_235 & popcount36_qqdr_core_234;
  assign popcount36_qqdr_core_239 = popcount36_qqdr_core_236 | popcount36_qqdr_core_238;
  assign popcount36_qqdr_core_242 = popcount36_qqdr_core_183 | popcount36_qqdr_core_239;
  assign popcount36_qqdr_core_243 = ~(input_a[34] & input_a[30]);
  assign popcount36_qqdr_core_246 = ~(input_a[34] ^ input_a[27]);
  assign popcount36_qqdr_core_247 = ~(input_a[7] | input_a[3]);
  assign popcount36_qqdr_core_250 = ~(input_a[15] | input_a[5]);
  assign popcount36_qqdr_core_251 = input_a[33] & input_a[1];
  assign popcount36_qqdr_core_252 = popcount36_qqdr_core_126 ^ popcount36_qqdr_core_232;
  assign popcount36_qqdr_core_253 = popcount36_qqdr_core_126 & popcount36_qqdr_core_232;
  assign popcount36_qqdr_core_254 = popcount36_qqdr_core_252 ^ input_a[33];
  assign popcount36_qqdr_core_255 = popcount36_qqdr_core_252 & input_a[33];
  assign popcount36_qqdr_core_256 = popcount36_qqdr_core_253 | popcount36_qqdr_core_255;
  assign popcount36_qqdr_core_257 = popcount36_qqdr_core_131 ^ popcount36_qqdr_core_237;
  assign popcount36_qqdr_core_258 = popcount36_qqdr_core_131 & popcount36_qqdr_core_237;
  assign popcount36_qqdr_core_259 = popcount36_qqdr_core_257 ^ popcount36_qqdr_core_256;
  assign popcount36_qqdr_core_260 = popcount36_qqdr_core_257 & popcount36_qqdr_core_256;
  assign popcount36_qqdr_core_261 = popcount36_qqdr_core_258 | popcount36_qqdr_core_260;
  assign popcount36_qqdr_core_262 = popcount36_qqdr_core_133 ^ popcount36_qqdr_core_242;
  assign popcount36_qqdr_core_263 = popcount36_qqdr_core_133 & popcount36_qqdr_core_242;
  assign popcount36_qqdr_core_264 = popcount36_qqdr_core_262 ^ popcount36_qqdr_core_261;
  assign popcount36_qqdr_core_265 = popcount36_qqdr_core_262 & popcount36_qqdr_core_261;
  assign popcount36_qqdr_core_266 = popcount36_qqdr_core_263 | popcount36_qqdr_core_265;
  assign popcount36_qqdr_core_268 = input_a[14] | input_a[1];
  assign popcount36_qqdr_core_270 = input_a[5] ^ input_a[7];
  assign popcount36_qqdr_core_271 = ~(input_a[35] | input_a[9]);
  assign popcount36_qqdr_core_272 = input_a[12] | input_a[9];
  assign popcount36_qqdr_core_274 = ~(input_a[5] ^ input_a[12]);
  assign popcount36_qqdr_core_275 = input_a[17] | input_a[30];
  assign popcount36_qqdr_core_276 = input_a[35] | input_a[14];

  assign popcount36_qqdr_out[0] = popcount36_qqdr_core_264;
  assign popcount36_qqdr_out[1] = popcount36_qqdr_core_254;
  assign popcount36_qqdr_out[2] = popcount36_qqdr_core_259;
  assign popcount36_qqdr_out[3] = popcount36_qqdr_core_264;
  assign popcount36_qqdr_out[4] = popcount36_qqdr_core_266;
  assign popcount36_qqdr_out[5] = 1'b0;
endmodule