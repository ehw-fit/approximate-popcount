// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.34411
// WCE=31.0
// EP=0.86233%
// Printed PDK parameters:
//  Area=100565385.0
//  Delay=90704800.0
//  Power=5205100.0

module popcount47_hpsm(input [46:0] input_a, output [5:0] popcount47_hpsm_out);
  wire popcount47_hpsm_core_050;
  wire popcount47_hpsm_core_051;
  wire popcount47_hpsm_core_052;
  wire popcount47_hpsm_core_053;
  wire popcount47_hpsm_core_055;
  wire popcount47_hpsm_core_056;
  wire popcount47_hpsm_core_059;
  wire popcount47_hpsm_core_060;
  wire popcount47_hpsm_core_064;
  wire popcount47_hpsm_core_065;
  wire popcount47_hpsm_core_066;
  wire popcount47_hpsm_core_067;
  wire popcount47_hpsm_core_068;
  wire popcount47_hpsm_core_069;
  wire popcount47_hpsm_core_070;
  wire popcount47_hpsm_core_071;
  wire popcount47_hpsm_core_072;
  wire popcount47_hpsm_core_073;
  wire popcount47_hpsm_core_074;
  wire popcount47_hpsm_core_077;
  wire popcount47_hpsm_core_078;
  wire popcount47_hpsm_core_079;
  wire popcount47_hpsm_core_080;
  wire popcount47_hpsm_core_081;
  wire popcount47_hpsm_core_082;
  wire popcount47_hpsm_core_083;
  wire popcount47_hpsm_core_084;
  wire popcount47_hpsm_core_086;
  wire popcount47_hpsm_core_087;
  wire popcount47_hpsm_core_088;
  wire popcount47_hpsm_core_089;
  wire popcount47_hpsm_core_090_not;
  wire popcount47_hpsm_core_092;
  wire popcount47_hpsm_core_093;
  wire popcount47_hpsm_core_097;
  wire popcount47_hpsm_core_098;
  wire popcount47_hpsm_core_099;
  wire popcount47_hpsm_core_100;
  wire popcount47_hpsm_core_101;
  wire popcount47_hpsm_core_103;
  wire popcount47_hpsm_core_104;
  wire popcount47_hpsm_core_107;
  wire popcount47_hpsm_core_108;
  wire popcount47_hpsm_core_110;
  wire popcount47_hpsm_core_111;
  wire popcount47_hpsm_core_114;
  wire popcount47_hpsm_core_115;
  wire popcount47_hpsm_core_121;
  wire popcount47_hpsm_core_122;
  wire popcount47_hpsm_core_131;
  wire popcount47_hpsm_core_132;
  wire popcount47_hpsm_core_133;
  wire popcount47_hpsm_core_134;
  wire popcount47_hpsm_core_135;
  wire popcount47_hpsm_core_136;
  wire popcount47_hpsm_core_137;
  wire popcount47_hpsm_core_138;
  wire popcount47_hpsm_core_140;
  wire popcount47_hpsm_core_142;
  wire popcount47_hpsm_core_145;
  wire popcount47_hpsm_core_146;
  wire popcount47_hpsm_core_150;
  wire popcount47_hpsm_core_151;
  wire popcount47_hpsm_core_152;
  wire popcount47_hpsm_core_153;
  wire popcount47_hpsm_core_157;
  wire popcount47_hpsm_core_158;
  wire popcount47_hpsm_core_159;
  wire popcount47_hpsm_core_160;
  wire popcount47_hpsm_core_161;
  wire popcount47_hpsm_core_162;
  wire popcount47_hpsm_core_163;
  wire popcount47_hpsm_core_164;
  wire popcount47_hpsm_core_165;
  wire popcount47_hpsm_core_166;
  wire popcount47_hpsm_core_168_not;
  wire popcount47_hpsm_core_170;
  wire popcount47_hpsm_core_171;
  wire popcount47_hpsm_core_173;
  wire popcount47_hpsm_core_174;
  wire popcount47_hpsm_core_175;
  wire popcount47_hpsm_core_176;
  wire popcount47_hpsm_core_177;
  wire popcount47_hpsm_core_178;
  wire popcount47_hpsm_core_179;
  wire popcount47_hpsm_core_180;
  wire popcount47_hpsm_core_181;
  wire popcount47_hpsm_core_182;
  wire popcount47_hpsm_core_183;
  wire popcount47_hpsm_core_184;
  wire popcount47_hpsm_core_186;
  wire popcount47_hpsm_core_187;
  wire popcount47_hpsm_core_189;
  wire popcount47_hpsm_core_190;
  wire popcount47_hpsm_core_191;
  wire popcount47_hpsm_core_192;
  wire popcount47_hpsm_core_193;
  wire popcount47_hpsm_core_194;
  wire popcount47_hpsm_core_195;
  wire popcount47_hpsm_core_196;
  wire popcount47_hpsm_core_197;
  wire popcount47_hpsm_core_198;
  wire popcount47_hpsm_core_199;
  wire popcount47_hpsm_core_200;
  wire popcount47_hpsm_core_201;
  wire popcount47_hpsm_core_202;
  wire popcount47_hpsm_core_203;
  wire popcount47_hpsm_core_205;
  wire popcount47_hpsm_core_207;
  wire popcount47_hpsm_core_208;
  wire popcount47_hpsm_core_209;
  wire popcount47_hpsm_core_210;
  wire popcount47_hpsm_core_211;
  wire popcount47_hpsm_core_212;
  wire popcount47_hpsm_core_213;
  wire popcount47_hpsm_core_214;
  wire popcount47_hpsm_core_215;
  wire popcount47_hpsm_core_216;
  wire popcount47_hpsm_core_217;
  wire popcount47_hpsm_core_220;
  wire popcount47_hpsm_core_221;
  wire popcount47_hpsm_core_222;
  wire popcount47_hpsm_core_225;
  wire popcount47_hpsm_core_227;
  wire popcount47_hpsm_core_231;
  wire popcount47_hpsm_core_234_not;
  wire popcount47_hpsm_core_235;
  wire popcount47_hpsm_core_236;
  wire popcount47_hpsm_core_237;
  wire popcount47_hpsm_core_240;
  wire popcount47_hpsm_core_241;
  wire popcount47_hpsm_core_244;
  wire popcount47_hpsm_core_245;
  wire popcount47_hpsm_core_249_not;
  wire popcount47_hpsm_core_251;
  wire popcount47_hpsm_core_252;
  wire popcount47_hpsm_core_253;
  wire popcount47_hpsm_core_254;
  wire popcount47_hpsm_core_255;
  wire popcount47_hpsm_core_256;
  wire popcount47_hpsm_core_259;
  wire popcount47_hpsm_core_260;
  wire popcount47_hpsm_core_261;
  wire popcount47_hpsm_core_262;
  wire popcount47_hpsm_core_263;
  wire popcount47_hpsm_core_264;
  wire popcount47_hpsm_core_265;
  wire popcount47_hpsm_core_266;
  wire popcount47_hpsm_core_267;
  wire popcount47_hpsm_core_268;
  wire popcount47_hpsm_core_269;
  wire popcount47_hpsm_core_270;
  wire popcount47_hpsm_core_273;
  wire popcount47_hpsm_core_274;
  wire popcount47_hpsm_core_278;
  wire popcount47_hpsm_core_279;
  wire popcount47_hpsm_core_280;
  wire popcount47_hpsm_core_281;
  wire popcount47_hpsm_core_282;
  wire popcount47_hpsm_core_283;
  wire popcount47_hpsm_core_284;
  wire popcount47_hpsm_core_285;
  wire popcount47_hpsm_core_286;
  wire popcount47_hpsm_core_287;
  wire popcount47_hpsm_core_288;
  wire popcount47_hpsm_core_289;
  wire popcount47_hpsm_core_290;
  wire popcount47_hpsm_core_291;
  wire popcount47_hpsm_core_292;
  wire popcount47_hpsm_core_293;
  wire popcount47_hpsm_core_294;
  wire popcount47_hpsm_core_295;
  wire popcount47_hpsm_core_296;
  wire popcount47_hpsm_core_297;
  wire popcount47_hpsm_core_298;
  wire popcount47_hpsm_core_299;
  wire popcount47_hpsm_core_300;
  wire popcount47_hpsm_core_301;
  wire popcount47_hpsm_core_302;
  wire popcount47_hpsm_core_304;
  wire popcount47_hpsm_core_305;
  wire popcount47_hpsm_core_306_not;
  wire popcount47_hpsm_core_307_not;
  wire popcount47_hpsm_core_309;
  wire popcount47_hpsm_core_310;
  wire popcount47_hpsm_core_311;
  wire popcount47_hpsm_core_312;
  wire popcount47_hpsm_core_313;
  wire popcount47_hpsm_core_314;
  wire popcount47_hpsm_core_315;
  wire popcount47_hpsm_core_316;
  wire popcount47_hpsm_core_317;
  wire popcount47_hpsm_core_318;
  wire popcount47_hpsm_core_322_not;
  wire popcount47_hpsm_core_324_not;
  wire popcount47_hpsm_core_326;
  wire popcount47_hpsm_core_327;
  wire popcount47_hpsm_core_328;
  wire popcount47_hpsm_core_329;
  wire popcount47_hpsm_core_330;
  wire popcount47_hpsm_core_331;
  wire popcount47_hpsm_core_332;
  wire popcount47_hpsm_core_333;
  wire popcount47_hpsm_core_334;
  wire popcount47_hpsm_core_335;
  wire popcount47_hpsm_core_336;
  wire popcount47_hpsm_core_337;
  wire popcount47_hpsm_core_338;
  wire popcount47_hpsm_core_339;
  wire popcount47_hpsm_core_340;
  wire popcount47_hpsm_core_344;
  wire popcount47_hpsm_core_345;
  wire popcount47_hpsm_core_347;
  wire popcount47_hpsm_core_348;
  wire popcount47_hpsm_core_349;
  wire popcount47_hpsm_core_350;
  wire popcount47_hpsm_core_351;
  wire popcount47_hpsm_core_352;
  wire popcount47_hpsm_core_353;
  wire popcount47_hpsm_core_354;
  wire popcount47_hpsm_core_355;
  wire popcount47_hpsm_core_356;
  wire popcount47_hpsm_core_357;
  wire popcount47_hpsm_core_358;
  wire popcount47_hpsm_core_359;
  wire popcount47_hpsm_core_360;
  wire popcount47_hpsm_core_361;
  wire popcount47_hpsm_core_362;
  wire popcount47_hpsm_core_363;
  wire popcount47_hpsm_core_364;
  wire popcount47_hpsm_core_365;
  wire popcount47_hpsm_core_366;
  wire popcount47_hpsm_core_367;
  wire popcount47_hpsm_core_369;
  wire popcount47_hpsm_core_370;
  wire popcount47_hpsm_core_371;

  assign popcount47_hpsm_core_050 = input_a[24] & input_a[1];
  assign popcount47_hpsm_core_051 = input_a[46] ^ input_a[39];
  assign popcount47_hpsm_core_052 = input_a[32] & input_a[4];
  assign popcount47_hpsm_core_053 = ~input_a[5];
  assign popcount47_hpsm_core_055 = popcount47_hpsm_core_052 ^ input_a[2];
  assign popcount47_hpsm_core_056 = popcount47_hpsm_core_052 & input_a[2];
  assign popcount47_hpsm_core_059 = popcount47_hpsm_core_050 ^ popcount47_hpsm_core_055;
  assign popcount47_hpsm_core_060 = popcount47_hpsm_core_050 & popcount47_hpsm_core_055;
  assign popcount47_hpsm_core_064 = popcount47_hpsm_core_056 ^ popcount47_hpsm_core_060;
  assign popcount47_hpsm_core_065 = popcount47_hpsm_core_056 & popcount47_hpsm_core_060;
  assign popcount47_hpsm_core_066 = input_a[6] ^ input_a[7];
  assign popcount47_hpsm_core_067 = input_a[6] & input_a[7];
  assign popcount47_hpsm_core_068 = input_a[5] ^ popcount47_hpsm_core_066;
  assign popcount47_hpsm_core_069 = input_a[5] & popcount47_hpsm_core_066;
  assign popcount47_hpsm_core_070 = popcount47_hpsm_core_067 ^ popcount47_hpsm_core_069;
  assign popcount47_hpsm_core_071 = popcount47_hpsm_core_067 & popcount47_hpsm_core_069;
  assign popcount47_hpsm_core_072 = input_a[30] ^ input_a[10];
  assign popcount47_hpsm_core_073 = input_a[9] & input_a[10];
  assign popcount47_hpsm_core_074 = input_a[16] | input_a[45];
  assign popcount47_hpsm_core_077 = ~(input_a[5] & input_a[19]);
  assign popcount47_hpsm_core_078 = popcount47_hpsm_core_068 | popcount47_hpsm_core_074;
  assign popcount47_hpsm_core_079 = popcount47_hpsm_core_068 & input_a[44];
  assign popcount47_hpsm_core_080 = popcount47_hpsm_core_070 ^ popcount47_hpsm_core_073;
  assign popcount47_hpsm_core_081 = popcount47_hpsm_core_070 & popcount47_hpsm_core_073;
  assign popcount47_hpsm_core_082 = popcount47_hpsm_core_080 ^ popcount47_hpsm_core_079;
  assign popcount47_hpsm_core_083 = popcount47_hpsm_core_080 & popcount47_hpsm_core_079;
  assign popcount47_hpsm_core_084 = popcount47_hpsm_core_081 | popcount47_hpsm_core_083;
  assign popcount47_hpsm_core_086 = popcount47_hpsm_core_071 & input_a[37];
  assign popcount47_hpsm_core_087 = popcount47_hpsm_core_071 ^ popcount47_hpsm_core_084;
  assign popcount47_hpsm_core_088 = popcount47_hpsm_core_071 & input_a[23];
  assign popcount47_hpsm_core_089 = popcount47_hpsm_core_086 | popcount47_hpsm_core_088;
  assign popcount47_hpsm_core_090_not = ~input_a[4];
  assign popcount47_hpsm_core_092 = popcount47_hpsm_core_059 ^ popcount47_hpsm_core_082;
  assign popcount47_hpsm_core_093 = popcount47_hpsm_core_059 & popcount47_hpsm_core_082;
  assign popcount47_hpsm_core_097 = popcount47_hpsm_core_064 ^ popcount47_hpsm_core_087;
  assign popcount47_hpsm_core_098 = popcount47_hpsm_core_064 & popcount47_hpsm_core_087;
  assign popcount47_hpsm_core_099 = popcount47_hpsm_core_097 ^ popcount47_hpsm_core_093;
  assign popcount47_hpsm_core_100 = popcount47_hpsm_core_097 & popcount47_hpsm_core_093;
  assign popcount47_hpsm_core_101 = popcount47_hpsm_core_098 | popcount47_hpsm_core_100;
  assign popcount47_hpsm_core_103 = input_a[40] & popcount47_hpsm_core_089;
  assign popcount47_hpsm_core_104 = popcount47_hpsm_core_065 ^ popcount47_hpsm_core_101;
  assign popcount47_hpsm_core_107 = input_a[12] ^ input_a[13];
  assign popcount47_hpsm_core_108 = input_a[12] & input_a[13];
  assign popcount47_hpsm_core_110 = input_a[11] & popcount47_hpsm_core_107;
  assign popcount47_hpsm_core_111 = popcount47_hpsm_core_108 | popcount47_hpsm_core_110;
  assign popcount47_hpsm_core_114 = input_a[15] & input_a[16];
  assign popcount47_hpsm_core_115 = input_a[45] & input_a[37];
  assign popcount47_hpsm_core_121 = popcount47_hpsm_core_111 ^ popcount47_hpsm_core_114;
  assign popcount47_hpsm_core_122 = popcount47_hpsm_core_111 & popcount47_hpsm_core_114;
  assign popcount47_hpsm_core_131 = ~(input_a[18] & input_a[19]);
  assign popcount47_hpsm_core_132 = input_a[18] & input_a[19];
  assign popcount47_hpsm_core_133 = input_a[17] ^ popcount47_hpsm_core_131;
  assign popcount47_hpsm_core_134 = input_a[17] & popcount47_hpsm_core_131;
  assign popcount47_hpsm_core_135 = popcount47_hpsm_core_132 | popcount47_hpsm_core_134;
  assign popcount47_hpsm_core_136 = popcount47_hpsm_core_132 & popcount47_hpsm_core_134;
  assign popcount47_hpsm_core_137 = ~input_a[21];
  assign popcount47_hpsm_core_138 = input_a[21] & input_a[22];
  assign popcount47_hpsm_core_140 = input_a[43] & popcount47_hpsm_core_137;
  assign popcount47_hpsm_core_142 = popcount47_hpsm_core_138 & popcount47_hpsm_core_140;
  assign popcount47_hpsm_core_145 = popcount47_hpsm_core_135 ^ popcount47_hpsm_core_138;
  assign popcount47_hpsm_core_146 = popcount47_hpsm_core_135 & popcount47_hpsm_core_138;
  assign popcount47_hpsm_core_150 = popcount47_hpsm_core_136 ^ popcount47_hpsm_core_142;
  assign popcount47_hpsm_core_151 = popcount47_hpsm_core_136 & input_a[29];
  assign popcount47_hpsm_core_152 = popcount47_hpsm_core_150 ^ popcount47_hpsm_core_146;
  assign popcount47_hpsm_core_153 = ~(popcount47_hpsm_core_150 | input_a[26]);
  assign popcount47_hpsm_core_157 = popcount47_hpsm_core_121 ^ popcount47_hpsm_core_145;
  assign popcount47_hpsm_core_158 = popcount47_hpsm_core_121 & popcount47_hpsm_core_145;
  assign popcount47_hpsm_core_159 = popcount47_hpsm_core_157 ^ popcount47_hpsm_core_133;
  assign popcount47_hpsm_core_160 = popcount47_hpsm_core_157 & popcount47_hpsm_core_133;
  assign popcount47_hpsm_core_161 = popcount47_hpsm_core_158 | popcount47_hpsm_core_160;
  assign popcount47_hpsm_core_162 = popcount47_hpsm_core_122 ^ popcount47_hpsm_core_152;
  assign popcount47_hpsm_core_163 = popcount47_hpsm_core_122 & popcount47_hpsm_core_152;
  assign popcount47_hpsm_core_164 = popcount47_hpsm_core_162 ^ popcount47_hpsm_core_161;
  assign popcount47_hpsm_core_165 = popcount47_hpsm_core_162 & popcount47_hpsm_core_161;
  assign popcount47_hpsm_core_166 = popcount47_hpsm_core_163 | popcount47_hpsm_core_165;
  assign popcount47_hpsm_core_168_not = ~input_a[31];
  assign popcount47_hpsm_core_170 = input_a[29] & input_a[40];
  assign popcount47_hpsm_core_171 = input_a[5] & input_a[10];
  assign popcount47_hpsm_core_173 = popcount47_hpsm_core_090_not & input_a[31];
  assign popcount47_hpsm_core_174 = popcount47_hpsm_core_092 ^ popcount47_hpsm_core_159;
  assign popcount47_hpsm_core_175 = popcount47_hpsm_core_092 & popcount47_hpsm_core_159;
  assign popcount47_hpsm_core_176 = popcount47_hpsm_core_174 ^ popcount47_hpsm_core_173;
  assign popcount47_hpsm_core_177 = popcount47_hpsm_core_174 & popcount47_hpsm_core_173;
  assign popcount47_hpsm_core_178 = popcount47_hpsm_core_175 | popcount47_hpsm_core_177;
  assign popcount47_hpsm_core_179 = popcount47_hpsm_core_099 ^ popcount47_hpsm_core_164;
  assign popcount47_hpsm_core_180 = popcount47_hpsm_core_099 & popcount47_hpsm_core_164;
  assign popcount47_hpsm_core_181 = popcount47_hpsm_core_179 ^ popcount47_hpsm_core_178;
  assign popcount47_hpsm_core_182 = popcount47_hpsm_core_179 & popcount47_hpsm_core_178;
  assign popcount47_hpsm_core_183 = popcount47_hpsm_core_180 | popcount47_hpsm_core_182;
  assign popcount47_hpsm_core_184 = popcount47_hpsm_core_104 ^ popcount47_hpsm_core_166;
  assign popcount47_hpsm_core_186 = popcount47_hpsm_core_184 ^ popcount47_hpsm_core_183;
  assign popcount47_hpsm_core_187 = popcount47_hpsm_core_184 & popcount47_hpsm_core_183;
  assign popcount47_hpsm_core_189 = popcount47_hpsm_core_103 & popcount47_hpsm_core_171;
  assign popcount47_hpsm_core_190 = popcount47_hpsm_core_103 & input_a[33];
  assign popcount47_hpsm_core_191 = popcount47_hpsm_core_189 | popcount47_hpsm_core_187;
  assign popcount47_hpsm_core_192 = popcount47_hpsm_core_189 & input_a[21];
  assign popcount47_hpsm_core_193 = popcount47_hpsm_core_190 | popcount47_hpsm_core_192;
  assign popcount47_hpsm_core_194 = ~input_a[44];
  assign popcount47_hpsm_core_195 = input_a[24] & input_a[25];
  assign popcount47_hpsm_core_196 = input_a[3] & input_a[14];
  assign popcount47_hpsm_core_197 = input_a[0] & popcount47_hpsm_core_194;
  assign popcount47_hpsm_core_198 = popcount47_hpsm_core_195 ^ popcount47_hpsm_core_197;
  assign popcount47_hpsm_core_199 = popcount47_hpsm_core_195 & popcount47_hpsm_core_197;
  assign popcount47_hpsm_core_200 = ~input_a[27];
  assign popcount47_hpsm_core_201 = input_a[34] & input_a[28];
  assign popcount47_hpsm_core_202 = ~input_a[26];
  assign popcount47_hpsm_core_203 = input_a[27] & popcount47_hpsm_core_200;
  assign popcount47_hpsm_core_205 = input_a[42] & popcount47_hpsm_core_203;
  assign popcount47_hpsm_core_207 = popcount47_hpsm_core_196 & input_a[43];
  assign popcount47_hpsm_core_208 = popcount47_hpsm_core_198 ^ popcount47_hpsm_core_201;
  assign popcount47_hpsm_core_209 = popcount47_hpsm_core_198 & popcount47_hpsm_core_201;
  assign popcount47_hpsm_core_210 = popcount47_hpsm_core_208 ^ popcount47_hpsm_core_207;
  assign popcount47_hpsm_core_211 = popcount47_hpsm_core_208 & popcount47_hpsm_core_207;
  assign popcount47_hpsm_core_212 = popcount47_hpsm_core_209 | popcount47_hpsm_core_211;
  assign popcount47_hpsm_core_213 = popcount47_hpsm_core_199 ^ popcount47_hpsm_core_205;
  assign popcount47_hpsm_core_214 = popcount47_hpsm_core_199 & input_a[44];
  assign popcount47_hpsm_core_215 = popcount47_hpsm_core_213 ^ popcount47_hpsm_core_212;
  assign popcount47_hpsm_core_216 = popcount47_hpsm_core_213 & input_a[31];
  assign popcount47_hpsm_core_217 = popcount47_hpsm_core_214 & input_a[30];
  assign popcount47_hpsm_core_220 = input_a[19] | input_a[40];
  assign popcount47_hpsm_core_221 = ~input_a[13];
  assign popcount47_hpsm_core_222 = input_a[4] ^ input_a[3];
  assign popcount47_hpsm_core_225 = ~(input_a[9] ^ input_a[43]);
  assign popcount47_hpsm_core_227 = ~(input_a[10] ^ input_a[5]);
  assign popcount47_hpsm_core_231 = input_a[29] & input_a[36];
  assign popcount47_hpsm_core_234_not = ~input_a[28];
  assign popcount47_hpsm_core_235 = ~(input_a[1] & input_a[25]);
  assign popcount47_hpsm_core_236 = input_a[15] | input_a[39];
  assign popcount47_hpsm_core_237 = input_a[24] ^ input_a[28];
  assign popcount47_hpsm_core_240 = input_a[19] & input_a[31];
  assign popcount47_hpsm_core_241 = input_a[38] | input_a[4];
  assign popcount47_hpsm_core_244 = popcount47_hpsm_core_210 ^ popcount47_hpsm_core_234_not;
  assign popcount47_hpsm_core_245 = popcount47_hpsm_core_210 & popcount47_hpsm_core_234_not;
  assign popcount47_hpsm_core_249_not = ~popcount47_hpsm_core_215;
  assign popcount47_hpsm_core_251 = popcount47_hpsm_core_249_not ^ popcount47_hpsm_core_245;
  assign popcount47_hpsm_core_252 = popcount47_hpsm_core_249_not & popcount47_hpsm_core_245;
  assign popcount47_hpsm_core_253 = popcount47_hpsm_core_215 | popcount47_hpsm_core_252;
  assign popcount47_hpsm_core_254 = popcount47_hpsm_core_217 & input_a[19];
  assign popcount47_hpsm_core_255 = input_a[15] ^ popcount47_hpsm_core_241;
  assign popcount47_hpsm_core_256 = popcount47_hpsm_core_254 ^ popcount47_hpsm_core_253;
  assign popcount47_hpsm_core_259 = ~(input_a[36] & input_a[6]);
  assign popcount47_hpsm_core_260 = input_a[36] & input_a[37];
  assign popcount47_hpsm_core_261 = input_a[36] & input_a[6];
  assign popcount47_hpsm_core_262 = input_a[35] & popcount47_hpsm_core_259;
  assign popcount47_hpsm_core_263 = popcount47_hpsm_core_260 ^ popcount47_hpsm_core_262;
  assign popcount47_hpsm_core_264 = popcount47_hpsm_core_260 & popcount47_hpsm_core_262;
  assign popcount47_hpsm_core_265 = input_a[39] ^ input_a[40];
  assign popcount47_hpsm_core_266 = input_a[39] & input_a[40];
  assign popcount47_hpsm_core_267 = ~(input_a[32] ^ input_a[31]);
  assign popcount47_hpsm_core_268 = input_a[38] & popcount47_hpsm_core_265;
  assign popcount47_hpsm_core_269 = popcount47_hpsm_core_266 ^ popcount47_hpsm_core_268;
  assign popcount47_hpsm_core_270 = popcount47_hpsm_core_266 & popcount47_hpsm_core_268;
  assign popcount47_hpsm_core_273 = popcount47_hpsm_core_263 ^ popcount47_hpsm_core_269;
  assign popcount47_hpsm_core_274 = popcount47_hpsm_core_263 & popcount47_hpsm_core_269;
  assign popcount47_hpsm_core_278 = popcount47_hpsm_core_264 | popcount47_hpsm_core_270;
  assign popcount47_hpsm_core_279 = ~(popcount47_hpsm_core_264 | input_a[1]);
  assign popcount47_hpsm_core_280 = popcount47_hpsm_core_278 ^ popcount47_hpsm_core_274;
  assign popcount47_hpsm_core_281 = input_a[32] & input_a[0];
  assign popcount47_hpsm_core_282 = input_a[12] | input_a[34];
  assign popcount47_hpsm_core_283 = ~(input_a[12] | input_a[43]);
  assign popcount47_hpsm_core_284 = input_a[28] & input_a[43];
  assign popcount47_hpsm_core_285 = input_a[41] ^ popcount47_hpsm_core_283;
  assign popcount47_hpsm_core_286 = input_a[42] & popcount47_hpsm_core_283;
  assign popcount47_hpsm_core_287 = popcount47_hpsm_core_284 | popcount47_hpsm_core_286;
  assign popcount47_hpsm_core_288 = popcount47_hpsm_core_284 & popcount47_hpsm_core_286;
  assign popcount47_hpsm_core_289 = input_a[45] ^ input_a[46];
  assign popcount47_hpsm_core_290 = input_a[45] & input_a[46];
  assign popcount47_hpsm_core_291 = input_a[44] ^ popcount47_hpsm_core_289;
  assign popcount47_hpsm_core_292 = input_a[44] & popcount47_hpsm_core_289;
  assign popcount47_hpsm_core_293 = popcount47_hpsm_core_290 ^ popcount47_hpsm_core_292;
  assign popcount47_hpsm_core_294 = popcount47_hpsm_core_290 & popcount47_hpsm_core_292;
  assign popcount47_hpsm_core_295 = popcount47_hpsm_core_285 ^ popcount47_hpsm_core_291;
  assign popcount47_hpsm_core_296 = popcount47_hpsm_core_285 & popcount47_hpsm_core_291;
  assign popcount47_hpsm_core_297 = popcount47_hpsm_core_287 ^ popcount47_hpsm_core_293;
  assign popcount47_hpsm_core_298 = popcount47_hpsm_core_287 & popcount47_hpsm_core_293;
  assign popcount47_hpsm_core_299 = popcount47_hpsm_core_297 ^ popcount47_hpsm_core_296;
  assign popcount47_hpsm_core_300 = popcount47_hpsm_core_297 & popcount47_hpsm_core_296;
  assign popcount47_hpsm_core_301 = popcount47_hpsm_core_298 | popcount47_hpsm_core_300;
  assign popcount47_hpsm_core_302 = popcount47_hpsm_core_288 ^ popcount47_hpsm_core_294;
  assign popcount47_hpsm_core_304 = popcount47_hpsm_core_302 ^ popcount47_hpsm_core_301;
  assign popcount47_hpsm_core_305 = popcount47_hpsm_core_302 & input_a[16];
  assign popcount47_hpsm_core_306_not = ~input_a[25];
  assign popcount47_hpsm_core_307_not = ~popcount47_hpsm_core_295;
  assign popcount47_hpsm_core_309 = popcount47_hpsm_core_273 ^ popcount47_hpsm_core_299;
  assign popcount47_hpsm_core_310 = popcount47_hpsm_core_273 & popcount47_hpsm_core_299;
  assign popcount47_hpsm_core_311 = popcount47_hpsm_core_309 ^ popcount47_hpsm_core_295;
  assign popcount47_hpsm_core_312 = popcount47_hpsm_core_309 & popcount47_hpsm_core_295;
  assign popcount47_hpsm_core_313 = popcount47_hpsm_core_310 | popcount47_hpsm_core_312;
  assign popcount47_hpsm_core_314 = popcount47_hpsm_core_280 ^ popcount47_hpsm_core_304;
  assign popcount47_hpsm_core_315 = popcount47_hpsm_core_280 & popcount47_hpsm_core_304;
  assign popcount47_hpsm_core_316 = popcount47_hpsm_core_314 ^ popcount47_hpsm_core_313;
  assign popcount47_hpsm_core_317 = popcount47_hpsm_core_314 & popcount47_hpsm_core_313;
  assign popcount47_hpsm_core_318 = popcount47_hpsm_core_315 | popcount47_hpsm_core_317;
  assign popcount47_hpsm_core_322_not = ~input_a[34];
  assign popcount47_hpsm_core_324_not = ~popcount47_hpsm_core_307_not;
  assign popcount47_hpsm_core_326 = popcount47_hpsm_core_244 ^ popcount47_hpsm_core_311;
  assign popcount47_hpsm_core_327 = popcount47_hpsm_core_244 & popcount47_hpsm_core_311;
  assign popcount47_hpsm_core_328 = popcount47_hpsm_core_326 ^ popcount47_hpsm_core_307_not;
  assign popcount47_hpsm_core_329 = popcount47_hpsm_core_326 & popcount47_hpsm_core_307_not;
  assign popcount47_hpsm_core_330 = popcount47_hpsm_core_327 | popcount47_hpsm_core_329;
  assign popcount47_hpsm_core_331 = popcount47_hpsm_core_251 ^ popcount47_hpsm_core_316;
  assign popcount47_hpsm_core_332 = popcount47_hpsm_core_251 & popcount47_hpsm_core_316;
  assign popcount47_hpsm_core_333 = popcount47_hpsm_core_331 ^ popcount47_hpsm_core_330;
  assign popcount47_hpsm_core_334 = popcount47_hpsm_core_331 & popcount47_hpsm_core_330;
  assign popcount47_hpsm_core_335 = popcount47_hpsm_core_332 | popcount47_hpsm_core_334;
  assign popcount47_hpsm_core_336 = popcount47_hpsm_core_256 ^ popcount47_hpsm_core_318;
  assign popcount47_hpsm_core_337 = popcount47_hpsm_core_256 & popcount47_hpsm_core_318;
  assign popcount47_hpsm_core_338 = popcount47_hpsm_core_336 ^ popcount47_hpsm_core_335;
  assign popcount47_hpsm_core_339 = popcount47_hpsm_core_336 & popcount47_hpsm_core_335;
  assign popcount47_hpsm_core_340 = popcount47_hpsm_core_337 | popcount47_hpsm_core_339;
  assign popcount47_hpsm_core_344 = input_a[26] | input_a[35];
  assign popcount47_hpsm_core_345 = ~input_a[20];
  assign popcount47_hpsm_core_347 = input_a[17] & popcount47_hpsm_core_324_not;
  assign popcount47_hpsm_core_348 = popcount47_hpsm_core_176 ^ popcount47_hpsm_core_328;
  assign popcount47_hpsm_core_349 = popcount47_hpsm_core_176 & popcount47_hpsm_core_328;
  assign popcount47_hpsm_core_350 = popcount47_hpsm_core_348 ^ popcount47_hpsm_core_347;
  assign popcount47_hpsm_core_351 = popcount47_hpsm_core_348 & popcount47_hpsm_core_347;
  assign popcount47_hpsm_core_352 = popcount47_hpsm_core_349 | popcount47_hpsm_core_351;
  assign popcount47_hpsm_core_353 = popcount47_hpsm_core_181 ^ popcount47_hpsm_core_333;
  assign popcount47_hpsm_core_354 = popcount47_hpsm_core_181 & popcount47_hpsm_core_333;
  assign popcount47_hpsm_core_355 = popcount47_hpsm_core_353 ^ popcount47_hpsm_core_352;
  assign popcount47_hpsm_core_356 = popcount47_hpsm_core_353 & popcount47_hpsm_core_352;
  assign popcount47_hpsm_core_357 = popcount47_hpsm_core_354 | popcount47_hpsm_core_356;
  assign popcount47_hpsm_core_358 = popcount47_hpsm_core_186 ^ popcount47_hpsm_core_338;
  assign popcount47_hpsm_core_359 = popcount47_hpsm_core_186 & popcount47_hpsm_core_338;
  assign popcount47_hpsm_core_360 = popcount47_hpsm_core_358 ^ popcount47_hpsm_core_357;
  assign popcount47_hpsm_core_361 = popcount47_hpsm_core_358 & popcount47_hpsm_core_357;
  assign popcount47_hpsm_core_362 = popcount47_hpsm_core_359 | popcount47_hpsm_core_361;
  assign popcount47_hpsm_core_363 = popcount47_hpsm_core_191 ^ popcount47_hpsm_core_340;
  assign popcount47_hpsm_core_364 = popcount47_hpsm_core_191 & popcount47_hpsm_core_340;
  assign popcount47_hpsm_core_365 = popcount47_hpsm_core_363 ^ popcount47_hpsm_core_362;
  assign popcount47_hpsm_core_366 = popcount47_hpsm_core_363 & popcount47_hpsm_core_362;
  assign popcount47_hpsm_core_367 = popcount47_hpsm_core_364 | popcount47_hpsm_core_366;
  assign popcount47_hpsm_core_369 = input_a[37] & popcount47_hpsm_core_345;
  assign popcount47_hpsm_core_370 = popcount47_hpsm_core_193 | popcount47_hpsm_core_367;
  assign popcount47_hpsm_core_371 = ~(input_a[25] | popcount47_hpsm_core_367);

  assign popcount47_hpsm_out[0] = popcount47_hpsm_core_362;
  assign popcount47_hpsm_out[1] = popcount47_hpsm_core_350;
  assign popcount47_hpsm_out[2] = popcount47_hpsm_core_355;
  assign popcount47_hpsm_out[3] = popcount47_hpsm_core_360;
  assign popcount47_hpsm_out[4] = popcount47_hpsm_core_365;
  assign popcount47_hpsm_out[5] = popcount47_hpsm_core_370;
endmodule