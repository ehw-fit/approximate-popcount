// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.59866
// WCE=13.0
// EP=0.976329%
// Printed PDK parameters:
//  Area=16730925.0
//  Delay=47947768.0
//  Power=840180.0

module popcount25_4jgj(input [24:0] input_a, output [4:0] popcount25_4jgj_out);
  wire popcount25_4jgj_core_028;
  wire popcount25_4jgj_core_030;
  wire popcount25_4jgj_core_031;
  wire popcount25_4jgj_core_032;
  wire popcount25_4jgj_core_033;
  wire popcount25_4jgj_core_034;
  wire popcount25_4jgj_core_035;
  wire popcount25_4jgj_core_036;
  wire popcount25_4jgj_core_037;
  wire popcount25_4jgj_core_038;
  wire popcount25_4jgj_core_039;
  wire popcount25_4jgj_core_040;
  wire popcount25_4jgj_core_041;
  wire popcount25_4jgj_core_042;
  wire popcount25_4jgj_core_043;
  wire popcount25_4jgj_core_044;
  wire popcount25_4jgj_core_045;
  wire popcount25_4jgj_core_047;
  wire popcount25_4jgj_core_049;
  wire popcount25_4jgj_core_050;
  wire popcount25_4jgj_core_051;
  wire popcount25_4jgj_core_052;
  wire popcount25_4jgj_core_054;
  wire popcount25_4jgj_core_055;
  wire popcount25_4jgj_core_057;
  wire popcount25_4jgj_core_059;
  wire popcount25_4jgj_core_060;
  wire popcount25_4jgj_core_062;
  wire popcount25_4jgj_core_063;
  wire popcount25_4jgj_core_066;
  wire popcount25_4jgj_core_068;
  wire popcount25_4jgj_core_069;
  wire popcount25_4jgj_core_070;
  wire popcount25_4jgj_core_071;
  wire popcount25_4jgj_core_072;
  wire popcount25_4jgj_core_075;
  wire popcount25_4jgj_core_076;
  wire popcount25_4jgj_core_077;
  wire popcount25_4jgj_core_078;
  wire popcount25_4jgj_core_080;
  wire popcount25_4jgj_core_082;
  wire popcount25_4jgj_core_083;
  wire popcount25_4jgj_core_084;
  wire popcount25_4jgj_core_085;
  wire popcount25_4jgj_core_086;
  wire popcount25_4jgj_core_089;
  wire popcount25_4jgj_core_090;
  wire popcount25_4jgj_core_091;
  wire popcount25_4jgj_core_092;
  wire popcount25_4jgj_core_095;
  wire popcount25_4jgj_core_096;
  wire popcount25_4jgj_core_097;
  wire popcount25_4jgj_core_098;
  wire popcount25_4jgj_core_099;
  wire popcount25_4jgj_core_100;
  wire popcount25_4jgj_core_103;
  wire popcount25_4jgj_core_104;
  wire popcount25_4jgj_core_106;
  wire popcount25_4jgj_core_107;
  wire popcount25_4jgj_core_109;
  wire popcount25_4jgj_core_110;
  wire popcount25_4jgj_core_111;
  wire popcount25_4jgj_core_115;
  wire popcount25_4jgj_core_117;
  wire popcount25_4jgj_core_119;
  wire popcount25_4jgj_core_121;
  wire popcount25_4jgj_core_123;
  wire popcount25_4jgj_core_127;
  wire popcount25_4jgj_core_129;
  wire popcount25_4jgj_core_131;
  wire popcount25_4jgj_core_135;
  wire popcount25_4jgj_core_136;
  wire popcount25_4jgj_core_137;
  wire popcount25_4jgj_core_138;
  wire popcount25_4jgj_core_139;
  wire popcount25_4jgj_core_143;
  wire popcount25_4jgj_core_148;
  wire popcount25_4jgj_core_150_not;
  wire popcount25_4jgj_core_151;
  wire popcount25_4jgj_core_152;
  wire popcount25_4jgj_core_153_not;
  wire popcount25_4jgj_core_154;
  wire popcount25_4jgj_core_156;
  wire popcount25_4jgj_core_157;
  wire popcount25_4jgj_core_159;
  wire popcount25_4jgj_core_160;
  wire popcount25_4jgj_core_161;
  wire popcount25_4jgj_core_162;
  wire popcount25_4jgj_core_163;
  wire popcount25_4jgj_core_164;
  wire popcount25_4jgj_core_165;
  wire popcount25_4jgj_core_166;
  wire popcount25_4jgj_core_167;
  wire popcount25_4jgj_core_169;
  wire popcount25_4jgj_core_170;
  wire popcount25_4jgj_core_171;
  wire popcount25_4jgj_core_172;
  wire popcount25_4jgj_core_173;
  wire popcount25_4jgj_core_174;
  wire popcount25_4jgj_core_175;
  wire popcount25_4jgj_core_177;
  wire popcount25_4jgj_core_178;
  wire popcount25_4jgj_core_179;
  wire popcount25_4jgj_core_180;
  wire popcount25_4jgj_core_181;
  wire popcount25_4jgj_core_183;

  assign popcount25_4jgj_core_028 = input_a[3] & input_a[9];
  assign popcount25_4jgj_core_030 = input_a[21] & input_a[0];
  assign popcount25_4jgj_core_031 = popcount25_4jgj_core_028 | popcount25_4jgj_core_030;
  assign popcount25_4jgj_core_032 = input_a[21] & input_a[10];
  assign popcount25_4jgj_core_033 = input_a[21] | input_a[22];
  assign popcount25_4jgj_core_034 = input_a[2] & input_a[24];
  assign popcount25_4jgj_core_035 = ~(input_a[11] ^ input_a[3]);
  assign popcount25_4jgj_core_036 = input_a[12] & input_a[5];
  assign popcount25_4jgj_core_037 = popcount25_4jgj_core_034 | popcount25_4jgj_core_036;
  assign popcount25_4jgj_core_038 = input_a[1] | input_a[12];
  assign popcount25_4jgj_core_039 = input_a[19] & input_a[20];
  assign popcount25_4jgj_core_040 = input_a[9] ^ input_a[10];
  assign popcount25_4jgj_core_041 = popcount25_4jgj_core_031 ^ popcount25_4jgj_core_037;
  assign popcount25_4jgj_core_042 = popcount25_4jgj_core_031 & popcount25_4jgj_core_037;
  assign popcount25_4jgj_core_043 = popcount25_4jgj_core_041 ^ input_a[20];
  assign popcount25_4jgj_core_044 = popcount25_4jgj_core_041 & input_a[20];
  assign popcount25_4jgj_core_045 = popcount25_4jgj_core_042 | popcount25_4jgj_core_044;
  assign popcount25_4jgj_core_047 = ~(input_a[14] | input_a[11]);
  assign popcount25_4jgj_core_049 = ~input_a[19];
  assign popcount25_4jgj_core_050 = ~input_a[13];
  assign popcount25_4jgj_core_051 = input_a[22] & input_a[8];
  assign popcount25_4jgj_core_052 = input_a[16] & input_a[1];
  assign popcount25_4jgj_core_054 = input_a[18] & input_a[19];
  assign popcount25_4jgj_core_055 = popcount25_4jgj_core_052 | popcount25_4jgj_core_054;
  assign popcount25_4jgj_core_057 = input_a[22] ^ input_a[15];
  assign popcount25_4jgj_core_059 = ~(input_a[20] & input_a[20]);
  assign popcount25_4jgj_core_060 = ~(input_a[21] | input_a[0]);
  assign popcount25_4jgj_core_062 = input_a[4] | input_a[21];
  assign popcount25_4jgj_core_063 = input_a[13] & input_a[18];
  assign popcount25_4jgj_core_066 = input_a[14] & input_a[15];
  assign popcount25_4jgj_core_068 = input_a[21] ^ input_a[4];
  assign popcount25_4jgj_core_069 = ~(input_a[17] & input_a[10]);
  assign popcount25_4jgj_core_070 = ~(input_a[5] | input_a[9]);
  assign popcount25_4jgj_core_071 = ~(input_a[0] ^ input_a[16]);
  assign popcount25_4jgj_core_072 = input_a[11] | input_a[14];
  assign popcount25_4jgj_core_075 = ~(input_a[5] & input_a[17]);
  assign popcount25_4jgj_core_076 = input_a[23] & input_a[13];
  assign popcount25_4jgj_core_077 = popcount25_4jgj_core_043 ^ popcount25_4jgj_core_055;
  assign popcount25_4jgj_core_078 = popcount25_4jgj_core_043 & popcount25_4jgj_core_055;
  assign popcount25_4jgj_core_080 = input_a[10] ^ input_a[5];
  assign popcount25_4jgj_core_082 = popcount25_4jgj_core_045 ^ popcount25_4jgj_core_072;
  assign popcount25_4jgj_core_083 = popcount25_4jgj_core_045 & popcount25_4jgj_core_072;
  assign popcount25_4jgj_core_084 = popcount25_4jgj_core_082 ^ popcount25_4jgj_core_078;
  assign popcount25_4jgj_core_085 = popcount25_4jgj_core_082 & popcount25_4jgj_core_078;
  assign popcount25_4jgj_core_086 = popcount25_4jgj_core_083 | popcount25_4jgj_core_085;
  assign popcount25_4jgj_core_089 = ~(input_a[16] ^ input_a[2]);
  assign popcount25_4jgj_core_090 = input_a[19] & input_a[3];
  assign popcount25_4jgj_core_091 = ~input_a[15];
  assign popcount25_4jgj_core_092 = ~(input_a[14] & input_a[21]);
  assign popcount25_4jgj_core_095 = ~(input_a[2] & input_a[22]);
  assign popcount25_4jgj_core_096 = ~input_a[21];
  assign popcount25_4jgj_core_097 = ~input_a[22];
  assign popcount25_4jgj_core_098 = ~input_a[2];
  assign popcount25_4jgj_core_099 = input_a[4] | input_a[17];
  assign popcount25_4jgj_core_100 = input_a[20] ^ input_a[21];
  assign popcount25_4jgj_core_103 = ~(input_a[12] | input_a[0]);
  assign popcount25_4jgj_core_104 = ~(input_a[1] ^ input_a[24]);
  assign popcount25_4jgj_core_106 = ~(input_a[8] | input_a[21]);
  assign popcount25_4jgj_core_107 = input_a[8] ^ input_a[22];
  assign popcount25_4jgj_core_109 = ~input_a[0];
  assign popcount25_4jgj_core_110 = input_a[11] ^ input_a[10];
  assign popcount25_4jgj_core_111 = ~(input_a[0] | input_a[19]);
  assign popcount25_4jgj_core_115 = ~(input_a[0] | input_a[17]);
  assign popcount25_4jgj_core_117 = input_a[4] | input_a[13];
  assign popcount25_4jgj_core_119 = ~(input_a[23] ^ input_a[19]);
  assign popcount25_4jgj_core_121 = ~input_a[15];
  assign popcount25_4jgj_core_123 = input_a[20] | input_a[19];
  assign popcount25_4jgj_core_127 = ~(input_a[10] | input_a[20]);
  assign popcount25_4jgj_core_129 = input_a[20] | input_a[16];
  assign popcount25_4jgj_core_131 = input_a[5] | input_a[7];
  assign popcount25_4jgj_core_135 = ~(input_a[20] ^ input_a[14]);
  assign popcount25_4jgj_core_136 = ~(input_a[1] & input_a[15]);
  assign popcount25_4jgj_core_137 = input_a[18] | input_a[11];
  assign popcount25_4jgj_core_138 = input_a[8] & input_a[23];
  assign popcount25_4jgj_core_139 = input_a[10] & popcount25_4jgj_core_138;
  assign popcount25_4jgj_core_143 = input_a[6] | input_a[14];
  assign popcount25_4jgj_core_148 = input_a[4] | input_a[10];
  assign popcount25_4jgj_core_150_not = ~input_a[0];
  assign popcount25_4jgj_core_151 = input_a[16] & input_a[23];
  assign popcount25_4jgj_core_152 = ~(input_a[6] & popcount25_4jgj_core_139);
  assign popcount25_4jgj_core_153_not = ~input_a[0];
  assign popcount25_4jgj_core_154 = ~popcount25_4jgj_core_152;
  assign popcount25_4jgj_core_156 = ~(input_a[21] & input_a[5]);
  assign popcount25_4jgj_core_157 = input_a[7] & input_a[1];
  assign popcount25_4jgj_core_159 = ~(input_a[8] | input_a[4]);
  assign popcount25_4jgj_core_160 = ~input_a[8];
  assign popcount25_4jgj_core_161 = ~(input_a[22] & input_a[18]);
  assign popcount25_4jgj_core_162 = ~(input_a[5] & input_a[3]);
  assign popcount25_4jgj_core_163 = ~input_a[9];
  assign popcount25_4jgj_core_164 = input_a[13] ^ input_a[19];
  assign popcount25_4jgj_core_165 = popcount25_4jgj_core_077 & input_a[13];
  assign popcount25_4jgj_core_166 = ~(input_a[13] & input_a[9]);
  assign popcount25_4jgj_core_167 = input_a[23] | input_a[3];
  assign popcount25_4jgj_core_169 = popcount25_4jgj_core_084 ^ popcount25_4jgj_core_154;
  assign popcount25_4jgj_core_170 = popcount25_4jgj_core_084 & popcount25_4jgj_core_154;
  assign popcount25_4jgj_core_171 = popcount25_4jgj_core_169 ^ popcount25_4jgj_core_165;
  assign popcount25_4jgj_core_172 = popcount25_4jgj_core_169 & popcount25_4jgj_core_165;
  assign popcount25_4jgj_core_173 = popcount25_4jgj_core_170 | popcount25_4jgj_core_172;
  assign popcount25_4jgj_core_174 = ~(input_a[4] | input_a[0]);
  assign popcount25_4jgj_core_175 = ~(input_a[6] | input_a[20]);
  assign popcount25_4jgj_core_177 = ~(input_a[7] & input_a[3]);
  assign popcount25_4jgj_core_178 = ~(input_a[1] | input_a[4]);
  assign popcount25_4jgj_core_179 = ~input_a[7];
  assign popcount25_4jgj_core_180 = ~(input_a[6] & input_a[7]);
  assign popcount25_4jgj_core_181 = input_a[9] | input_a[23];
  assign popcount25_4jgj_core_183 = ~(input_a[13] & input_a[23]);

  assign popcount25_4jgj_out[0] = input_a[4];
  assign popcount25_4jgj_out[1] = popcount25_4jgj_core_047;
  assign popcount25_4jgj_out[2] = popcount25_4jgj_core_171;
  assign popcount25_4jgj_out[3] = popcount25_4jgj_core_173;
  assign popcount25_4jgj_out[4] = popcount25_4jgj_core_086;
endmodule