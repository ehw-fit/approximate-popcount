// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.53154
// WCE=23.0
// EP=0.983879%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_6er0(input [26:0] input_a, output [4:0] popcount27_6er0_out);
  wire popcount27_6er0_core_029;
  wire popcount27_6er0_core_031;
  wire popcount27_6er0_core_033;
  wire popcount27_6er0_core_035;
  wire popcount27_6er0_core_038;
  wire popcount27_6er0_core_039;
  wire popcount27_6er0_core_040;
  wire popcount27_6er0_core_041;
  wire popcount27_6er0_core_043;
  wire popcount27_6er0_core_046;
  wire popcount27_6er0_core_052;
  wire popcount27_6er0_core_054;
  wire popcount27_6er0_core_056;
  wire popcount27_6er0_core_057;
  wire popcount27_6er0_core_058;
  wire popcount27_6er0_core_059;
  wire popcount27_6er0_core_061;
  wire popcount27_6er0_core_065;
  wire popcount27_6er0_core_067;
  wire popcount27_6er0_core_068;
  wire popcount27_6er0_core_069;
  wire popcount27_6er0_core_070;
  wire popcount27_6er0_core_072;
  wire popcount27_6er0_core_073;
  wire popcount27_6er0_core_075_not;
  wire popcount27_6er0_core_077;
  wire popcount27_6er0_core_079;
  wire popcount27_6er0_core_080;
  wire popcount27_6er0_core_081;
  wire popcount27_6er0_core_082;
  wire popcount27_6er0_core_083;
  wire popcount27_6er0_core_086;
  wire popcount27_6er0_core_092;
  wire popcount27_6er0_core_093;
  wire popcount27_6er0_core_094;
  wire popcount27_6er0_core_095;
  wire popcount27_6er0_core_097;
  wire popcount27_6er0_core_098;
  wire popcount27_6er0_core_099;
  wire popcount27_6er0_core_100;
  wire popcount27_6er0_core_101;
  wire popcount27_6er0_core_103;
  wire popcount27_6er0_core_104;
  wire popcount27_6er0_core_106;
  wire popcount27_6er0_core_107;
  wire popcount27_6er0_core_110;
  wire popcount27_6er0_core_113;
  wire popcount27_6er0_core_114;
  wire popcount27_6er0_core_117;
  wire popcount27_6er0_core_118;
  wire popcount27_6er0_core_119;
  wire popcount27_6er0_core_122;
  wire popcount27_6er0_core_123;
  wire popcount27_6er0_core_124;
  wire popcount27_6er0_core_127_not;
  wire popcount27_6er0_core_128;
  wire popcount27_6er0_core_131;
  wire popcount27_6er0_core_132;
  wire popcount27_6er0_core_133;
  wire popcount27_6er0_core_135;
  wire popcount27_6er0_core_136;
  wire popcount27_6er0_core_137;
  wire popcount27_6er0_core_138;
  wire popcount27_6er0_core_139;
  wire popcount27_6er0_core_140;
  wire popcount27_6er0_core_142;
  wire popcount27_6er0_core_145;
  wire popcount27_6er0_core_146;
  wire popcount27_6er0_core_149;
  wire popcount27_6er0_core_152;
  wire popcount27_6er0_core_153;
  wire popcount27_6er0_core_156;
  wire popcount27_6er0_core_157;
  wire popcount27_6er0_core_160;
  wire popcount27_6er0_core_163;
  wire popcount27_6er0_core_164;
  wire popcount27_6er0_core_168;
  wire popcount27_6er0_core_171;
  wire popcount27_6er0_core_172;
  wire popcount27_6er0_core_173;
  wire popcount27_6er0_core_174;
  wire popcount27_6er0_core_175;
  wire popcount27_6er0_core_177;
  wire popcount27_6er0_core_178;
  wire popcount27_6er0_core_179;
  wire popcount27_6er0_core_180;
  wire popcount27_6er0_core_182;
  wire popcount27_6er0_core_183;
  wire popcount27_6er0_core_185;
  wire popcount27_6er0_core_186;
  wire popcount27_6er0_core_191;

  assign popcount27_6er0_core_029 = input_a[25] & input_a[22];
  assign popcount27_6er0_core_031 = input_a[25] ^ input_a[20];
  assign popcount27_6er0_core_033 = ~(input_a[19] & input_a[6]);
  assign popcount27_6er0_core_035 = input_a[5] | input_a[6];
  assign popcount27_6er0_core_038 = input_a[17] & input_a[21];
  assign popcount27_6er0_core_039 = ~(input_a[26] & input_a[13]);
  assign popcount27_6er0_core_040 = ~(input_a[9] & input_a[21]);
  assign popcount27_6er0_core_041 = ~(input_a[11] ^ input_a[1]);
  assign popcount27_6er0_core_043 = input_a[23] & input_a[26];
  assign popcount27_6er0_core_046 = ~(input_a[1] ^ input_a[20]);
  assign popcount27_6er0_core_052 = ~(input_a[26] ^ input_a[1]);
  assign popcount27_6er0_core_054 = input_a[25] ^ input_a[21];
  assign popcount27_6er0_core_056 = input_a[23] | input_a[2];
  assign popcount27_6er0_core_057 = ~input_a[9];
  assign popcount27_6er0_core_058 = input_a[5] | input_a[20];
  assign popcount27_6er0_core_059 = input_a[10] | input_a[3];
  assign popcount27_6er0_core_061 = ~input_a[3];
  assign popcount27_6er0_core_065 = ~input_a[20];
  assign popcount27_6er0_core_067 = ~(input_a[26] & input_a[12]);
  assign popcount27_6er0_core_068 = ~(input_a[6] ^ input_a[13]);
  assign popcount27_6er0_core_069 = ~(input_a[11] & input_a[5]);
  assign popcount27_6er0_core_070 = input_a[13] ^ input_a[16];
  assign popcount27_6er0_core_072 = ~(input_a[21] & input_a[10]);
  assign popcount27_6er0_core_073 = input_a[22] & input_a[15];
  assign popcount27_6er0_core_075_not = ~input_a[14];
  assign popcount27_6er0_core_077 = ~input_a[22];
  assign popcount27_6er0_core_079 = ~input_a[21];
  assign popcount27_6er0_core_080 = ~input_a[20];
  assign popcount27_6er0_core_081 = ~input_a[23];
  assign popcount27_6er0_core_082 = ~(input_a[16] | input_a[7]);
  assign popcount27_6er0_core_083 = input_a[4] | input_a[19];
  assign popcount27_6er0_core_086 = ~input_a[5];
  assign popcount27_6er0_core_092 = ~(input_a[4] & input_a[12]);
  assign popcount27_6er0_core_093 = ~(input_a[18] | input_a[16]);
  assign popcount27_6er0_core_094 = ~(input_a[23] | input_a[21]);
  assign popcount27_6er0_core_095 = ~(input_a[19] | input_a[10]);
  assign popcount27_6er0_core_097 = ~(input_a[22] | input_a[6]);
  assign popcount27_6er0_core_098 = input_a[4] ^ input_a[25];
  assign popcount27_6er0_core_099 = ~(input_a[1] ^ input_a[3]);
  assign popcount27_6er0_core_100 = input_a[2] ^ input_a[26];
  assign popcount27_6er0_core_101 = ~(input_a[22] | input_a[18]);
  assign popcount27_6er0_core_103 = ~input_a[20];
  assign popcount27_6er0_core_104 = input_a[1] & input_a[18];
  assign popcount27_6er0_core_106 = ~input_a[20];
  assign popcount27_6er0_core_107 = input_a[18] | input_a[26];
  assign popcount27_6er0_core_110 = input_a[11] & input_a[14];
  assign popcount27_6er0_core_113 = input_a[22] & input_a[24];
  assign popcount27_6er0_core_114 = ~input_a[4];
  assign popcount27_6er0_core_117 = input_a[26] ^ input_a[22];
  assign popcount27_6er0_core_118 = ~(input_a[8] | input_a[11]);
  assign popcount27_6er0_core_119 = ~input_a[26];
  assign popcount27_6er0_core_122 = ~(input_a[14] | input_a[12]);
  assign popcount27_6er0_core_123 = ~(input_a[23] & input_a[22]);
  assign popcount27_6er0_core_124 = input_a[16] ^ input_a[12];
  assign popcount27_6er0_core_127_not = ~input_a[15];
  assign popcount27_6er0_core_128 = input_a[24] | input_a[1];
  assign popcount27_6er0_core_131 = ~input_a[24];
  assign popcount27_6er0_core_132 = input_a[3] ^ input_a[25];
  assign popcount27_6er0_core_133 = ~(input_a[24] & input_a[7]);
  assign popcount27_6er0_core_135 = input_a[16] ^ input_a[24];
  assign popcount27_6er0_core_136 = input_a[0] | input_a[7];
  assign popcount27_6er0_core_137 = input_a[11] & input_a[16];
  assign popcount27_6er0_core_138 = input_a[12] | input_a[13];
  assign popcount27_6er0_core_139 = ~(input_a[24] ^ input_a[11]);
  assign popcount27_6er0_core_140 = ~(input_a[3] | input_a[12]);
  assign popcount27_6er0_core_142 = input_a[5] ^ input_a[1];
  assign popcount27_6er0_core_145 = ~(input_a[19] & input_a[1]);
  assign popcount27_6er0_core_146 = ~(input_a[5] ^ input_a[21]);
  assign popcount27_6er0_core_149 = ~input_a[16];
  assign popcount27_6er0_core_152 = ~(input_a[17] & input_a[18]);
  assign popcount27_6er0_core_153 = ~(input_a[3] | input_a[25]);
  assign popcount27_6er0_core_156 = ~(input_a[15] & input_a[11]);
  assign popcount27_6er0_core_157 = ~input_a[18];
  assign popcount27_6er0_core_160 = input_a[21] ^ input_a[20];
  assign popcount27_6er0_core_163 = input_a[5] | input_a[9];
  assign popcount27_6er0_core_164 = ~(input_a[24] ^ input_a[15]);
  assign popcount27_6er0_core_168 = input_a[7] ^ input_a[9];
  assign popcount27_6er0_core_171 = input_a[21] & input_a[2];
  assign popcount27_6er0_core_172 = ~input_a[18];
  assign popcount27_6er0_core_173 = input_a[23] & input_a[22];
  assign popcount27_6er0_core_174 = ~(input_a[18] ^ input_a[15]);
  assign popcount27_6er0_core_175 = ~(input_a[0] ^ input_a[26]);
  assign popcount27_6er0_core_177 = ~(input_a[14] | input_a[6]);
  assign popcount27_6er0_core_178 = ~(input_a[17] | input_a[8]);
  assign popcount27_6er0_core_179 = ~(input_a[13] | input_a[4]);
  assign popcount27_6er0_core_180 = input_a[8] ^ input_a[23];
  assign popcount27_6er0_core_182 = ~(input_a[16] ^ input_a[3]);
  assign popcount27_6er0_core_183 = input_a[11] | input_a[10];
  assign popcount27_6er0_core_185 = ~(input_a[26] | input_a[7]);
  assign popcount27_6er0_core_186 = ~(input_a[1] & input_a[23]);
  assign popcount27_6er0_core_191 = ~input_a[23];

  assign popcount27_6er0_out[0] = input_a[1];
  assign popcount27_6er0_out[1] = 1'b0;
  assign popcount27_6er0_out[2] = 1'b0;
  assign popcount27_6er0_out[3] = 1'b1;
  assign popcount27_6er0_out[4] = input_a[6];
endmodule