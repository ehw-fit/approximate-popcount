// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.37596
// WCE=23.0
// EP=0.932675%
// Printed PDK parameters:
//  Area=57556947.0
//  Delay=67009888.0
//  Power=2993400.0

module popcount45_xey9(input [44:0] input_a, output [5:0] popcount45_xey9_out);
  wire popcount45_xey9_core_047;
  wire popcount45_xey9_core_048;
  wire popcount45_xey9_core_049;
  wire popcount45_xey9_core_050;
  wire popcount45_xey9_core_051;
  wire popcount45_xey9_core_052;
  wire popcount45_xey9_core_053;
  wire popcount45_xey9_core_055;
  wire popcount45_xey9_core_056;
  wire popcount45_xey9_core_057;
  wire popcount45_xey9_core_058;
  wire popcount45_xey9_core_060;
  wire popcount45_xey9_core_061;
  wire popcount45_xey9_core_064;
  wire popcount45_xey9_core_065;
  wire popcount45_xey9_core_066;
  wire popcount45_xey9_core_067;
  wire popcount45_xey9_core_068;
  wire popcount45_xey9_core_070;
  wire popcount45_xey9_core_071;
  wire popcount45_xey9_core_072;
  wire popcount45_xey9_core_073;
  wire popcount45_xey9_core_074;
  wire popcount45_xey9_core_075;
  wire popcount45_xey9_core_077;
  wire popcount45_xey9_core_079;
  wire popcount45_xey9_core_084;
  wire popcount45_xey9_core_087;
  wire popcount45_xey9_core_088;
  wire popcount45_xey9_core_089;
  wire popcount45_xey9_core_090;
  wire popcount45_xey9_core_091;
  wire popcount45_xey9_core_093;
  wire popcount45_xey9_core_094;
  wire popcount45_xey9_core_095;
  wire popcount45_xey9_core_096;
  wire popcount45_xey9_core_098;
  wire popcount45_xey9_core_099;
  wire popcount45_xey9_core_101;
  wire popcount45_xey9_core_103;
  wire popcount45_xey9_core_104;
  wire popcount45_xey9_core_106;
  wire popcount45_xey9_core_107;
  wire popcount45_xey9_core_108;
  wire popcount45_xey9_core_109;
  wire popcount45_xey9_core_110;
  wire popcount45_xey9_core_111;
  wire popcount45_xey9_core_115;
  wire popcount45_xey9_core_116;
  wire popcount45_xey9_core_121;
  wire popcount45_xey9_core_122;
  wire popcount45_xey9_core_123;
  wire popcount45_xey9_core_124;
  wire popcount45_xey9_core_125;
  wire popcount45_xey9_core_126;
  wire popcount45_xey9_core_127;
  wire popcount45_xey9_core_129;
  wire popcount45_xey9_core_133_not;
  wire popcount45_xey9_core_135;
  wire popcount45_xey9_core_136;
  wire popcount45_xey9_core_137;
  wire popcount45_xey9_core_138;
  wire popcount45_xey9_core_139;
  wire popcount45_xey9_core_140;
  wire popcount45_xey9_core_144;
  wire popcount45_xey9_core_147;
  wire popcount45_xey9_core_148;
  wire popcount45_xey9_core_149;
  wire popcount45_xey9_core_150;
  wire popcount45_xey9_core_151;
  wire popcount45_xey9_core_152;
  wire popcount45_xey9_core_153;
  wire popcount45_xey9_core_154;
  wire popcount45_xey9_core_155;
  wire popcount45_xey9_core_156;
  wire popcount45_xey9_core_157;
  wire popcount45_xey9_core_161;
  wire popcount45_xey9_core_162;
  wire popcount45_xey9_core_165_not;
  wire popcount45_xey9_core_172;
  wire popcount45_xey9_core_173;
  wire popcount45_xey9_core_175;
  wire popcount45_xey9_core_176;
  wire popcount45_xey9_core_183;
  wire popcount45_xey9_core_185;
  wire popcount45_xey9_core_186;
  wire popcount45_xey9_core_187;
  wire popcount45_xey9_core_188;
  wire popcount45_xey9_core_190;
  wire popcount45_xey9_core_191;
  wire popcount45_xey9_core_192;
  wire popcount45_xey9_core_195;
  wire popcount45_xey9_core_196;
  wire popcount45_xey9_core_200;
  wire popcount45_xey9_core_202;
  wire popcount45_xey9_core_203;
  wire popcount45_xey9_core_204;
  wire popcount45_xey9_core_205;
  wire popcount45_xey9_core_206;
  wire popcount45_xey9_core_207;
  wire popcount45_xey9_core_208;
  wire popcount45_xey9_core_209;
  wire popcount45_xey9_core_210;
  wire popcount45_xey9_core_211;
  wire popcount45_xey9_core_212;
  wire popcount45_xey9_core_213;
  wire popcount45_xey9_core_215;
  wire popcount45_xey9_core_217;
  wire popcount45_xey9_core_221;
  wire popcount45_xey9_core_223;
  wire popcount45_xey9_core_224;
  wire popcount45_xey9_core_226;
  wire popcount45_xey9_core_227;
  wire popcount45_xey9_core_228;
  wire popcount45_xey9_core_230;
  wire popcount45_xey9_core_231;
  wire popcount45_xey9_core_233;
  wire popcount45_xey9_core_234;
  wire popcount45_xey9_core_235;
  wire popcount45_xey9_core_236;
  wire popcount45_xey9_core_237;
  wire popcount45_xey9_core_239;
  wire popcount45_xey9_core_240_not;
  wire popcount45_xey9_core_242;
  wire popcount45_xey9_core_245;
  wire popcount45_xey9_core_247;
  wire popcount45_xey9_core_248_not;
  wire popcount45_xey9_core_249;
  wire popcount45_xey9_core_250;
  wire popcount45_xey9_core_251;
  wire popcount45_xey9_core_252;
  wire popcount45_xey9_core_253;
  wire popcount45_xey9_core_254;
  wire popcount45_xey9_core_258;
  wire popcount45_xey9_core_259_not;
  wire popcount45_xey9_core_260;
  wire popcount45_xey9_core_262;
  wire popcount45_xey9_core_263;
  wire popcount45_xey9_core_264;
  wire popcount45_xey9_core_267;
  wire popcount45_xey9_core_268;
  wire popcount45_xey9_core_269;
  wire popcount45_xey9_core_270;
  wire popcount45_xey9_core_272;
  wire popcount45_xey9_core_274;
  wire popcount45_xey9_core_275;
  wire popcount45_xey9_core_279;
  wire popcount45_xey9_core_280;
  wire popcount45_xey9_core_281;
  wire popcount45_xey9_core_282;
  wire popcount45_xey9_core_285;
  wire popcount45_xey9_core_286;
  wire popcount45_xey9_core_287;
  wire popcount45_xey9_core_288;
  wire popcount45_xey9_core_290;
  wire popcount45_xey9_core_293;
  wire popcount45_xey9_core_296;
  wire popcount45_xey9_core_297;
  wire popcount45_xey9_core_298;
  wire popcount45_xey9_core_299;
  wire popcount45_xey9_core_300;
  wire popcount45_xey9_core_301;
  wire popcount45_xey9_core_302;
  wire popcount45_xey9_core_303;
  wire popcount45_xey9_core_304;
  wire popcount45_xey9_core_306;
  wire popcount45_xey9_core_308;
  wire popcount45_xey9_core_309;
  wire popcount45_xey9_core_310;
  wire popcount45_xey9_core_311;
  wire popcount45_xey9_core_312;
  wire popcount45_xey9_core_313;
  wire popcount45_xey9_core_314;
  wire popcount45_xey9_core_315;
  wire popcount45_xey9_core_316;
  wire popcount45_xey9_core_317;
  wire popcount45_xey9_core_318;
  wire popcount45_xey9_core_319;
  wire popcount45_xey9_core_322;
  wire popcount45_xey9_core_323;
  wire popcount45_xey9_core_327;
  wire popcount45_xey9_core_330;
  wire popcount45_xey9_core_331;
  wire popcount45_xey9_core_333;
  wire popcount45_xey9_core_335;
  wire popcount45_xey9_core_338;
  wire popcount45_xey9_core_342;
  wire popcount45_xey9_core_343;
  wire popcount45_xey9_core_344;
  wire popcount45_xey9_core_345;
  wire popcount45_xey9_core_346;
  wire popcount45_xey9_core_347;
  wire popcount45_xey9_core_348;
  wire popcount45_xey9_core_349;
  wire popcount45_xey9_core_350;
  wire popcount45_xey9_core_351;
  wire popcount45_xey9_core_353;
  wire popcount45_xey9_core_355;

  assign popcount45_xey9_core_047 = input_a[0] ^ input_a[1];
  assign popcount45_xey9_core_048 = input_a[0] & input_a[1];
  assign popcount45_xey9_core_049 = input_a[40] ^ input_a[4];
  assign popcount45_xey9_core_050 = input_a[3] & input_a[4];
  assign popcount45_xey9_core_051 = ~(input_a[2] & input_a[14]);
  assign popcount45_xey9_core_052 = input_a[2] & popcount45_xey9_core_049;
  assign popcount45_xey9_core_053 = popcount45_xey9_core_050 ^ popcount45_xey9_core_052;
  assign popcount45_xey9_core_055 = ~(input_a[25] ^ input_a[7]);
  assign popcount45_xey9_core_056 = popcount45_xey9_core_047 & input_a[38];
  assign popcount45_xey9_core_057 = popcount45_xey9_core_048 ^ popcount45_xey9_core_053;
  assign popcount45_xey9_core_058 = popcount45_xey9_core_048 & popcount45_xey9_core_053;
  assign popcount45_xey9_core_060 = popcount45_xey9_core_057 & popcount45_xey9_core_056;
  assign popcount45_xey9_core_061 = popcount45_xey9_core_058 | popcount45_xey9_core_060;
  assign popcount45_xey9_core_064 = input_a[6] ^ input_a[7];
  assign popcount45_xey9_core_065 = input_a[6] & input_a[7];
  assign popcount45_xey9_core_066 = ~(input_a[22] & popcount45_xey9_core_064);
  assign popcount45_xey9_core_067 = input_a[5] & popcount45_xey9_core_064;
  assign popcount45_xey9_core_068 = popcount45_xey9_core_065 ^ popcount45_xey9_core_067;
  assign popcount45_xey9_core_070 = input_a[9] ^ input_a[10];
  assign popcount45_xey9_core_071 = input_a[9] & input_a[10];
  assign popcount45_xey9_core_072 = ~input_a[14];
  assign popcount45_xey9_core_073 = input_a[43] & popcount45_xey9_core_070;
  assign popcount45_xey9_core_074 = popcount45_xey9_core_071 ^ popcount45_xey9_core_073;
  assign popcount45_xey9_core_075 = ~(input_a[6] | popcount45_xey9_core_073);
  assign popcount45_xey9_core_077 = input_a[8] & input_a[37];
  assign popcount45_xey9_core_079 = popcount45_xey9_core_068 & popcount45_xey9_core_074;
  assign popcount45_xey9_core_084 = ~(input_a[37] & popcount45_xey9_core_075);
  assign popcount45_xey9_core_087 = input_a[43] & input_a[4];
  assign popcount45_xey9_core_088 = input_a[12] ^ input_a[19];
  assign popcount45_xey9_core_089 = input_a[32] & input_a[22];
  assign popcount45_xey9_core_090 = ~(input_a[24] | popcount45_xey9_core_077);
  assign popcount45_xey9_core_091 = input_a[1] & popcount45_xey9_core_077;
  assign popcount45_xey9_core_093 = input_a[35] & input_a[33];
  assign popcount45_xey9_core_094 = popcount45_xey9_core_091 | popcount45_xey9_core_093;
  assign popcount45_xey9_core_095 = popcount45_xey9_core_061 ^ popcount45_xey9_core_079;
  assign popcount45_xey9_core_096 = popcount45_xey9_core_061 & popcount45_xey9_core_079;
  assign popcount45_xey9_core_098 = popcount45_xey9_core_095 & popcount45_xey9_core_094;
  assign popcount45_xey9_core_099 = popcount45_xey9_core_096 | popcount45_xey9_core_098;
  assign popcount45_xey9_core_101 = input_a[24] & input_a[8];
  assign popcount45_xey9_core_103 = ~(input_a[9] ^ input_a[30]);
  assign popcount45_xey9_core_104 = input_a[25] | input_a[13];
  assign popcount45_xey9_core_106 = input_a[11] & input_a[12];
  assign popcount45_xey9_core_107 = input_a[14] ^ input_a[15];
  assign popcount45_xey9_core_108 = input_a[14] & input_a[15];
  assign popcount45_xey9_core_109 = input_a[13] ^ popcount45_xey9_core_107;
  assign popcount45_xey9_core_110 = input_a[13] & popcount45_xey9_core_107;
  assign popcount45_xey9_core_111 = popcount45_xey9_core_108 ^ popcount45_xey9_core_110;
  assign popcount45_xey9_core_115 = popcount45_xey9_core_106 ^ popcount45_xey9_core_111;
  assign popcount45_xey9_core_116 = popcount45_xey9_core_106 & popcount45_xey9_core_111;
  assign popcount45_xey9_core_121 = ~(input_a[35] & input_a[25]);
  assign popcount45_xey9_core_122 = input_a[17] ^ input_a[17];
  assign popcount45_xey9_core_123 = input_a[17] & input_a[18];
  assign popcount45_xey9_core_124 = input_a[16] ^ popcount45_xey9_core_122;
  assign popcount45_xey9_core_125 = input_a[16] & popcount45_xey9_core_122;
  assign popcount45_xey9_core_126 = popcount45_xey9_core_123 ^ popcount45_xey9_core_125;
  assign popcount45_xey9_core_127 = ~(input_a[32] | input_a[11]);
  assign popcount45_xey9_core_129 = input_a[20] & input_a[21];
  assign popcount45_xey9_core_133_not = ~input_a[39];
  assign popcount45_xey9_core_135 = popcount45_xey9_core_124 & input_a[23];
  assign popcount45_xey9_core_136 = popcount45_xey9_core_126 ^ popcount45_xey9_core_129;
  assign popcount45_xey9_core_137 = popcount45_xey9_core_126 & popcount45_xey9_core_129;
  assign popcount45_xey9_core_138 = popcount45_xey9_core_136 ^ popcount45_xey9_core_135;
  assign popcount45_xey9_core_139 = popcount45_xey9_core_136 & popcount45_xey9_core_135;
  assign popcount45_xey9_core_140 = popcount45_xey9_core_137 | popcount45_xey9_core_139;
  assign popcount45_xey9_core_144 = ~input_a[26];
  assign popcount45_xey9_core_147 = popcount45_xey9_core_109 & input_a[36];
  assign popcount45_xey9_core_148 = popcount45_xey9_core_115 ^ popcount45_xey9_core_138;
  assign popcount45_xey9_core_149 = popcount45_xey9_core_115 & popcount45_xey9_core_138;
  assign popcount45_xey9_core_150 = ~(input_a[39] & popcount45_xey9_core_147);
  assign popcount45_xey9_core_151 = popcount45_xey9_core_148 & popcount45_xey9_core_147;
  assign popcount45_xey9_core_152 = popcount45_xey9_core_149 | popcount45_xey9_core_151;
  assign popcount45_xey9_core_153 = popcount45_xey9_core_116 ^ popcount45_xey9_core_140;
  assign popcount45_xey9_core_154 = popcount45_xey9_core_116 & popcount45_xey9_core_140;
  assign popcount45_xey9_core_155 = ~(popcount45_xey9_core_153 | popcount45_xey9_core_152);
  assign popcount45_xey9_core_156 = popcount45_xey9_core_153 & popcount45_xey9_core_152;
  assign popcount45_xey9_core_157 = popcount45_xey9_core_154 | popcount45_xey9_core_156;
  assign popcount45_xey9_core_161 = ~(input_a[43] & input_a[26]);
  assign popcount45_xey9_core_162 = input_a[30] & input_a[40];
  assign popcount45_xey9_core_165_not = ~popcount45_xey9_core_150;
  assign popcount45_xey9_core_172 = popcount45_xey9_core_155 | popcount45_xey9_core_150;
  assign popcount45_xey9_core_173 = ~(input_a[32] & input_a[9]);
  assign popcount45_xey9_core_175 = popcount45_xey9_core_099 ^ popcount45_xey9_core_157;
  assign popcount45_xey9_core_176 = popcount45_xey9_core_099 & popcount45_xey9_core_157;
  assign popcount45_xey9_core_183 = input_a[38] | input_a[14];
  assign popcount45_xey9_core_185 = ~(input_a[43] ^ input_a[23]);
  assign popcount45_xey9_core_186 = input_a[9] ^ input_a[23];
  assign popcount45_xey9_core_187 = input_a[25] ^ input_a[26];
  assign popcount45_xey9_core_188 = input_a[25] & input_a[26];
  assign popcount45_xey9_core_190 = input_a[24] & popcount45_xey9_core_187;
  assign popcount45_xey9_core_191 = popcount45_xey9_core_188 | popcount45_xey9_core_190;
  assign popcount45_xey9_core_192 = popcount45_xey9_core_188 & popcount45_xey9_core_190;
  assign popcount45_xey9_core_195 = ~(input_a[2] | popcount45_xey9_core_191);
  assign popcount45_xey9_core_196 = input_a[39] & popcount45_xey9_core_191;
  assign popcount45_xey9_core_200 = popcount45_xey9_core_192 | popcount45_xey9_core_196;
  assign popcount45_xey9_core_202 = input_a[28] ^ input_a[29];
  assign popcount45_xey9_core_203 = input_a[28] & input_a[29];
  assign popcount45_xey9_core_204 = input_a[27] ^ popcount45_xey9_core_202;
  assign popcount45_xey9_core_205 = input_a[27] & popcount45_xey9_core_202;
  assign popcount45_xey9_core_206 = popcount45_xey9_core_203 ^ popcount45_xey9_core_205;
  assign popcount45_xey9_core_207 = popcount45_xey9_core_203 & popcount45_xey9_core_205;
  assign popcount45_xey9_core_208 = input_a[11] ^ input_a[17];
  assign popcount45_xey9_core_209 = input_a[31] & input_a[32];
  assign popcount45_xey9_core_210 = ~(input_a[13] | input_a[38]);
  assign popcount45_xey9_core_211 = input_a[30] & input_a[44];
  assign popcount45_xey9_core_212 = popcount45_xey9_core_209 | popcount45_xey9_core_211;
  assign popcount45_xey9_core_213 = popcount45_xey9_core_209 & popcount45_xey9_core_211;
  assign popcount45_xey9_core_215 = input_a[29] & input_a[9];
  assign popcount45_xey9_core_217 = popcount45_xey9_core_206 & popcount45_xey9_core_212;
  assign popcount45_xey9_core_221 = popcount45_xey9_core_207 | popcount45_xey9_core_213;
  assign popcount45_xey9_core_223 = popcount45_xey9_core_221 | popcount45_xey9_core_217;
  assign popcount45_xey9_core_224 = ~input_a[23];
  assign popcount45_xey9_core_226 = input_a[22] ^ popcount45_xey9_core_204;
  assign popcount45_xey9_core_227 = input_a[22] & popcount45_xey9_core_204;
  assign popcount45_xey9_core_228 = ~popcount45_xey9_core_195;
  assign popcount45_xey9_core_230 = popcount45_xey9_core_228 ^ popcount45_xey9_core_227;
  assign popcount45_xey9_core_231 = popcount45_xey9_core_228 & popcount45_xey9_core_227;
  assign popcount45_xey9_core_233 = popcount45_xey9_core_200 ^ popcount45_xey9_core_223;
  assign popcount45_xey9_core_234 = popcount45_xey9_core_200 & popcount45_xey9_core_223;
  assign popcount45_xey9_core_235 = popcount45_xey9_core_233 ^ popcount45_xey9_core_231;
  assign popcount45_xey9_core_236 = popcount45_xey9_core_233 & popcount45_xey9_core_231;
  assign popcount45_xey9_core_237 = popcount45_xey9_core_234 | popcount45_xey9_core_236;
  assign popcount45_xey9_core_239 = popcount45_xey9_core_192 & input_a[26];
  assign popcount45_xey9_core_240_not = ~popcount45_xey9_core_237;
  assign popcount45_xey9_core_242 = popcount45_xey9_core_239 | popcount45_xey9_core_237;
  assign popcount45_xey9_core_245 = input_a[42] & input_a[11];
  assign popcount45_xey9_core_247 = ~(input_a[30] & input_a[34]);
  assign popcount45_xey9_core_248_not = ~input_a[26];
  assign popcount45_xey9_core_249 = input_a[10] ^ input_a[22];
  assign popcount45_xey9_core_250 = ~input_a[37];
  assign popcount45_xey9_core_251 = ~(input_a[21] | input_a[44]);
  assign popcount45_xey9_core_252 = ~(input_a[18] ^ input_a[33]);
  assign popcount45_xey9_core_253 = input_a[34] & input_a[21];
  assign popcount45_xey9_core_254 = input_a[17] | input_a[31];
  assign popcount45_xey9_core_258 = input_a[17] & input_a[12];
  assign popcount45_xey9_core_259_not = ~input_a[8];
  assign popcount45_xey9_core_260 = ~(input_a[43] & input_a[30]);
  assign popcount45_xey9_core_262 = input_a[15] ^ input_a[36];
  assign popcount45_xey9_core_263 = ~(input_a[4] & input_a[12]);
  assign popcount45_xey9_core_264 = input_a[28] & input_a[42];
  assign popcount45_xey9_core_267 = input_a[41] & input_a[33];
  assign popcount45_xey9_core_268 = input_a[32] | input_a[18];
  assign popcount45_xey9_core_269 = ~(input_a[39] | input_a[32]);
  assign popcount45_xey9_core_270 = input_a[29] ^ input_a[37];
  assign popcount45_xey9_core_272 = input_a[14] & input_a[13];
  assign popcount45_xey9_core_274 = ~(input_a[2] | input_a[30]);
  assign popcount45_xey9_core_275 = input_a[30] & input_a[31];
  assign popcount45_xey9_core_279 = input_a[43] ^ input_a[25];
  assign popcount45_xey9_core_280 = ~(input_a[3] | input_a[19]);
  assign popcount45_xey9_core_281 = input_a[27] ^ input_a[0];
  assign popcount45_xey9_core_282 = input_a[19] ^ input_a[44];
  assign popcount45_xey9_core_285 = ~(input_a[3] ^ input_a[18]);
  assign popcount45_xey9_core_286 = input_a[29] & input_a[30];
  assign popcount45_xey9_core_287 = ~(input_a[26] ^ input_a[0]);
  assign popcount45_xey9_core_288 = input_a[26] ^ input_a[12];
  assign popcount45_xey9_core_290 = ~(input_a[5] & input_a[44]);
  assign popcount45_xey9_core_293 = input_a[16] | input_a[8];
  assign popcount45_xey9_core_296 = ~(input_a[32] | input_a[26]);
  assign popcount45_xey9_core_297 = input_a[25] | input_a[44];
  assign popcount45_xey9_core_298 = input_a[35] | input_a[4];
  assign popcount45_xey9_core_299 = input_a[39] ^ input_a[41];
  assign popcount45_xey9_core_300 = input_a[41] ^ input_a[36];
  assign popcount45_xey9_core_301 = ~(input_a[9] ^ input_a[9]);
  assign popcount45_xey9_core_302 = ~input_a[11];
  assign popcount45_xey9_core_303 = input_a[32] & input_a[20];
  assign popcount45_xey9_core_304 = input_a[40] ^ input_a[36];
  assign popcount45_xey9_core_306 = ~(input_a[22] & input_a[13]);
  assign popcount45_xey9_core_308 = input_a[12] & input_a[12];
  assign popcount45_xey9_core_309 = popcount45_xey9_core_226 & input_a[36];
  assign popcount45_xey9_core_310 = popcount45_xey9_core_230 ^ input_a[42];
  assign popcount45_xey9_core_311 = popcount45_xey9_core_230 & input_a[42];
  assign popcount45_xey9_core_312 = popcount45_xey9_core_310 ^ popcount45_xey9_core_309;
  assign popcount45_xey9_core_313 = popcount45_xey9_core_310 & popcount45_xey9_core_309;
  assign popcount45_xey9_core_314 = popcount45_xey9_core_311 | popcount45_xey9_core_313;
  assign popcount45_xey9_core_315 = popcount45_xey9_core_235 ^ popcount45_xey9_core_300;
  assign popcount45_xey9_core_316 = popcount45_xey9_core_235 & popcount45_xey9_core_300;
  assign popcount45_xey9_core_317 = popcount45_xey9_core_315 ^ popcount45_xey9_core_314;
  assign popcount45_xey9_core_318 = popcount45_xey9_core_315 & popcount45_xey9_core_314;
  assign popcount45_xey9_core_319 = popcount45_xey9_core_316 | popcount45_xey9_core_318;
  assign popcount45_xey9_core_322 = popcount45_xey9_core_240_not ^ popcount45_xey9_core_319;
  assign popcount45_xey9_core_323 = popcount45_xey9_core_240_not & popcount45_xey9_core_319;
  assign popcount45_xey9_core_327 = popcount45_xey9_core_242 | popcount45_xey9_core_323;
  assign popcount45_xey9_core_330 = input_a[6] ^ input_a[6];
  assign popcount45_xey9_core_331 = ~input_a[13];
  assign popcount45_xey9_core_333 = popcount45_xey9_core_165_not & input_a[41];
  assign popcount45_xey9_core_335 = ~(input_a[27] & input_a[13]);
  assign popcount45_xey9_core_338 = popcount45_xey9_core_172 & popcount45_xey9_core_317;
  assign popcount45_xey9_core_342 = popcount45_xey9_core_175 ^ popcount45_xey9_core_322;
  assign popcount45_xey9_core_343 = popcount45_xey9_core_175 & popcount45_xey9_core_322;
  assign popcount45_xey9_core_344 = popcount45_xey9_core_342 ^ popcount45_xey9_core_338;
  assign popcount45_xey9_core_345 = popcount45_xey9_core_342 & popcount45_xey9_core_338;
  assign popcount45_xey9_core_346 = popcount45_xey9_core_343 | popcount45_xey9_core_345;
  assign popcount45_xey9_core_347 = popcount45_xey9_core_176 ^ popcount45_xey9_core_327;
  assign popcount45_xey9_core_348 = popcount45_xey9_core_176 & popcount45_xey9_core_327;
  assign popcount45_xey9_core_349 = popcount45_xey9_core_347 ^ popcount45_xey9_core_346;
  assign popcount45_xey9_core_350 = popcount45_xey9_core_347 & popcount45_xey9_core_346;
  assign popcount45_xey9_core_351 = popcount45_xey9_core_348 | popcount45_xey9_core_350;
  assign popcount45_xey9_core_353 = ~(input_a[17] ^ input_a[40]);
  assign popcount45_xey9_core_355 = ~(input_a[33] | popcount45_xey9_core_351);

  assign popcount45_xey9_out[0] = 1'b0;
  assign popcount45_xey9_out[1] = 1'b1;
  assign popcount45_xey9_out[2] = popcount45_xey9_core_333;
  assign popcount45_xey9_out[3] = popcount45_xey9_core_344;
  assign popcount45_xey9_out[4] = popcount45_xey9_core_349;
  assign popcount45_xey9_out[5] = popcount45_xey9_core_351;
endmodule