// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.87902
// WCE=28.0
// EP=0.965807%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_jlfi(input [20:0] input_a, output [4:0] popcount21_jlfi_out);
  wire popcount21_jlfi_core_023_not;
  wire popcount21_jlfi_core_024_not;
  wire popcount21_jlfi_core_025;
  wire popcount21_jlfi_core_026;
  wire popcount21_jlfi_core_027;
  wire popcount21_jlfi_core_029;
  wire popcount21_jlfi_core_036;
  wire popcount21_jlfi_core_037;
  wire popcount21_jlfi_core_038;
  wire popcount21_jlfi_core_039;
  wire popcount21_jlfi_core_041;
  wire popcount21_jlfi_core_043;
  wire popcount21_jlfi_core_046;
  wire popcount21_jlfi_core_048;
  wire popcount21_jlfi_core_050;
  wire popcount21_jlfi_core_052;
  wire popcount21_jlfi_core_053;
  wire popcount21_jlfi_core_054;
  wire popcount21_jlfi_core_055;
  wire popcount21_jlfi_core_056;
  wire popcount21_jlfi_core_057;
  wire popcount21_jlfi_core_058;
  wire popcount21_jlfi_core_059;
  wire popcount21_jlfi_core_060;
  wire popcount21_jlfi_core_061;
  wire popcount21_jlfi_core_062;
  wire popcount21_jlfi_core_063;
  wire popcount21_jlfi_core_064;
  wire popcount21_jlfi_core_065;
  wire popcount21_jlfi_core_066;
  wire popcount21_jlfi_core_067;
  wire popcount21_jlfi_core_068;
  wire popcount21_jlfi_core_069;
  wire popcount21_jlfi_core_070;
  wire popcount21_jlfi_core_072;
  wire popcount21_jlfi_core_074;
  wire popcount21_jlfi_core_077;
  wire popcount21_jlfi_core_078;
  wire popcount21_jlfi_core_079;
  wire popcount21_jlfi_core_081;
  wire popcount21_jlfi_core_082;
  wire popcount21_jlfi_core_083;
  wire popcount21_jlfi_core_085;
  wire popcount21_jlfi_core_087;
  wire popcount21_jlfi_core_090;
  wire popcount21_jlfi_core_092;
  wire popcount21_jlfi_core_093;
  wire popcount21_jlfi_core_096;
  wire popcount21_jlfi_core_097;
  wire popcount21_jlfi_core_100;
  wire popcount21_jlfi_core_102;
  wire popcount21_jlfi_core_103;
  wire popcount21_jlfi_core_105;
  wire popcount21_jlfi_core_106;
  wire popcount21_jlfi_core_108;
  wire popcount21_jlfi_core_109;
  wire popcount21_jlfi_core_111;
  wire popcount21_jlfi_core_112;
  wire popcount21_jlfi_core_114;
  wire popcount21_jlfi_core_116;
  wire popcount21_jlfi_core_118;
  wire popcount21_jlfi_core_120;
  wire popcount21_jlfi_core_121;
  wire popcount21_jlfi_core_124;
  wire popcount21_jlfi_core_125;
  wire popcount21_jlfi_core_127;
  wire popcount21_jlfi_core_131;
  wire popcount21_jlfi_core_132;
  wire popcount21_jlfi_core_135;
  wire popcount21_jlfi_core_136;
  wire popcount21_jlfi_core_137;
  wire popcount21_jlfi_core_138;
  wire popcount21_jlfi_core_139;
  wire popcount21_jlfi_core_141;
  wire popcount21_jlfi_core_142;
  wire popcount21_jlfi_core_143;
  wire popcount21_jlfi_core_146;
  wire popcount21_jlfi_core_147;
  wire popcount21_jlfi_core_148;
  wire popcount21_jlfi_core_149;
  wire popcount21_jlfi_core_150;
  wire popcount21_jlfi_core_152;
  wire popcount21_jlfi_core_153;

  assign popcount21_jlfi_core_023_not = ~input_a[16];
  assign popcount21_jlfi_core_024_not = ~input_a[7];
  assign popcount21_jlfi_core_025 = ~(input_a[13] | input_a[6]);
  assign popcount21_jlfi_core_026 = input_a[14] ^ input_a[2];
  assign popcount21_jlfi_core_027 = ~input_a[8];
  assign popcount21_jlfi_core_029 = input_a[1] ^ input_a[12];
  assign popcount21_jlfi_core_036 = ~(input_a[19] ^ input_a[13]);
  assign popcount21_jlfi_core_037 = ~(input_a[10] ^ input_a[1]);
  assign popcount21_jlfi_core_038 = input_a[4] ^ input_a[14];
  assign popcount21_jlfi_core_039 = input_a[5] | input_a[5];
  assign popcount21_jlfi_core_041 = ~(input_a[9] | input_a[10]);
  assign popcount21_jlfi_core_043 = ~input_a[14];
  assign popcount21_jlfi_core_046 = ~(input_a[18] ^ input_a[6]);
  assign popcount21_jlfi_core_048 = ~(input_a[9] | input_a[13]);
  assign popcount21_jlfi_core_050 = ~(input_a[12] & input_a[5]);
  assign popcount21_jlfi_core_052 = input_a[9] ^ input_a[19];
  assign popcount21_jlfi_core_053 = input_a[8] & input_a[20];
  assign popcount21_jlfi_core_054 = ~(input_a[6] | input_a[3]);
  assign popcount21_jlfi_core_055 = ~input_a[11];
  assign popcount21_jlfi_core_056 = input_a[1] & input_a[5];
  assign popcount21_jlfi_core_057 = ~(input_a[6] & input_a[9]);
  assign popcount21_jlfi_core_058 = ~(input_a[3] | input_a[13]);
  assign popcount21_jlfi_core_059 = ~(input_a[19] | input_a[4]);
  assign popcount21_jlfi_core_060 = input_a[3] ^ input_a[17];
  assign popcount21_jlfi_core_061 = ~input_a[13];
  assign popcount21_jlfi_core_062 = ~(input_a[20] & input_a[3]);
  assign popcount21_jlfi_core_063 = input_a[0] & input_a[10];
  assign popcount21_jlfi_core_064 = ~input_a[4];
  assign popcount21_jlfi_core_065 = ~(input_a[1] ^ input_a[18]);
  assign popcount21_jlfi_core_066 = ~(input_a[7] ^ input_a[6]);
  assign popcount21_jlfi_core_067 = ~(input_a[14] & input_a[0]);
  assign popcount21_jlfi_core_068 = input_a[19] ^ input_a[5];
  assign popcount21_jlfi_core_069 = ~(input_a[8] | input_a[8]);
  assign popcount21_jlfi_core_070 = ~input_a[12];
  assign popcount21_jlfi_core_072 = ~(input_a[7] | input_a[12]);
  assign popcount21_jlfi_core_074 = ~(input_a[1] & input_a[2]);
  assign popcount21_jlfi_core_077 = ~(input_a[20] & input_a[14]);
  assign popcount21_jlfi_core_078 = input_a[20] & input_a[11];
  assign popcount21_jlfi_core_079 = ~(input_a[9] ^ input_a[10]);
  assign popcount21_jlfi_core_081 = ~input_a[3];
  assign popcount21_jlfi_core_082 = input_a[11] ^ input_a[14];
  assign popcount21_jlfi_core_083 = input_a[20] | input_a[16];
  assign popcount21_jlfi_core_085 = ~input_a[4];
  assign popcount21_jlfi_core_087 = ~input_a[18];
  assign popcount21_jlfi_core_090 = input_a[8] | input_a[14];
  assign popcount21_jlfi_core_092 = ~(input_a[2] & input_a[9]);
  assign popcount21_jlfi_core_093 = ~(input_a[16] ^ input_a[20]);
  assign popcount21_jlfi_core_096 = ~(input_a[2] & input_a[0]);
  assign popcount21_jlfi_core_097 = ~(input_a[15] ^ input_a[17]);
  assign popcount21_jlfi_core_100 = ~(input_a[0] | input_a[14]);
  assign popcount21_jlfi_core_102 = ~(input_a[12] | input_a[3]);
  assign popcount21_jlfi_core_103 = ~(input_a[7] ^ input_a[20]);
  assign popcount21_jlfi_core_105 = ~(input_a[15] | input_a[14]);
  assign popcount21_jlfi_core_106 = input_a[14] ^ input_a[0];
  assign popcount21_jlfi_core_108 = ~(input_a[3] & input_a[15]);
  assign popcount21_jlfi_core_109 = ~input_a[11];
  assign popcount21_jlfi_core_111 = ~(input_a[5] & input_a[20]);
  assign popcount21_jlfi_core_112 = ~(input_a[20] | input_a[16]);
  assign popcount21_jlfi_core_114 = ~input_a[13];
  assign popcount21_jlfi_core_116 = input_a[13] & input_a[4];
  assign popcount21_jlfi_core_118 = ~input_a[5];
  assign popcount21_jlfi_core_120 = ~input_a[4];
  assign popcount21_jlfi_core_121 = input_a[8] ^ input_a[2];
  assign popcount21_jlfi_core_124 = ~(input_a[5] | input_a[13]);
  assign popcount21_jlfi_core_125 = ~input_a[18];
  assign popcount21_jlfi_core_127 = ~(input_a[17] ^ input_a[19]);
  assign popcount21_jlfi_core_131 = ~(input_a[17] & input_a[13]);
  assign popcount21_jlfi_core_132 = input_a[10] | input_a[2];
  assign popcount21_jlfi_core_135 = input_a[16] | input_a[0];
  assign popcount21_jlfi_core_136 = input_a[4] | input_a[3];
  assign popcount21_jlfi_core_137 = ~(input_a[18] & input_a[6]);
  assign popcount21_jlfi_core_138 = ~(input_a[13] & input_a[3]);
  assign popcount21_jlfi_core_139 = ~(input_a[17] | input_a[4]);
  assign popcount21_jlfi_core_141 = input_a[4] | input_a[20];
  assign popcount21_jlfi_core_142 = ~input_a[18];
  assign popcount21_jlfi_core_143 = ~(input_a[11] & input_a[15]);
  assign popcount21_jlfi_core_146 = ~input_a[11];
  assign popcount21_jlfi_core_147 = ~(input_a[4] & input_a[15]);
  assign popcount21_jlfi_core_148 = input_a[0] ^ input_a[14];
  assign popcount21_jlfi_core_149 = ~(input_a[7] & input_a[16]);
  assign popcount21_jlfi_core_150 = ~(input_a[19] & input_a[3]);
  assign popcount21_jlfi_core_152 = ~(input_a[20] ^ input_a[6]);
  assign popcount21_jlfi_core_153 = input_a[9] ^ input_a[12];

  assign popcount21_jlfi_out[0] = 1'b1;
  assign popcount21_jlfi_out[1] = 1'b1;
  assign popcount21_jlfi_out[2] = input_a[5];
  assign popcount21_jlfi_out[3] = input_a[0];
  assign popcount21_jlfi_out[4] = input_a[19];
endmodule