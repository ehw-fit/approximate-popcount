// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.00693
// WCE=20.0
// EP=0.993878%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_0c31(input [23:0] input_a, output [4:0] popcount24_0c31_out);
  wire popcount24_0c31_core_027_not;
  wire popcount24_0c31_core_028;
  wire popcount24_0c31_core_030;
  wire popcount24_0c31_core_034;
  wire popcount24_0c31_core_035;
  wire popcount24_0c31_core_037;
  wire popcount24_0c31_core_038;
  wire popcount24_0c31_core_039;
  wire popcount24_0c31_core_040;
  wire popcount24_0c31_core_041;
  wire popcount24_0c31_core_042;
  wire popcount24_0c31_core_043_not;
  wire popcount24_0c31_core_044;
  wire popcount24_0c31_core_045;
  wire popcount24_0c31_core_046;
  wire popcount24_0c31_core_047;
  wire popcount24_0c31_core_048;
  wire popcount24_0c31_core_053;
  wire popcount24_0c31_core_055_not;
  wire popcount24_0c31_core_056;
  wire popcount24_0c31_core_058;
  wire popcount24_0c31_core_059_not;
  wire popcount24_0c31_core_061;
  wire popcount24_0c31_core_062;
  wire popcount24_0c31_core_065;
  wire popcount24_0c31_core_066_not;
  wire popcount24_0c31_core_068;
  wire popcount24_0c31_core_069;
  wire popcount24_0c31_core_072;
  wire popcount24_0c31_core_074;
  wire popcount24_0c31_core_076;
  wire popcount24_0c31_core_077;
  wire popcount24_0c31_core_078;
  wire popcount24_0c31_core_080;
  wire popcount24_0c31_core_081;
  wire popcount24_0c31_core_083;
  wire popcount24_0c31_core_084;
  wire popcount24_0c31_core_086;
  wire popcount24_0c31_core_087;
  wire popcount24_0c31_core_089;
  wire popcount24_0c31_core_090;
  wire popcount24_0c31_core_092;
  wire popcount24_0c31_core_093;
  wire popcount24_0c31_core_094;
  wire popcount24_0c31_core_096;
  wire popcount24_0c31_core_097;
  wire popcount24_0c31_core_099;
  wire popcount24_0c31_core_100;
  wire popcount24_0c31_core_101;
  wire popcount24_0c31_core_102;
  wire popcount24_0c31_core_106;
  wire popcount24_0c31_core_112;
  wire popcount24_0c31_core_114;
  wire popcount24_0c31_core_115;
  wire popcount24_0c31_core_116;
  wire popcount24_0c31_core_117;
  wire popcount24_0c31_core_119;
  wire popcount24_0c31_core_120;
  wire popcount24_0c31_core_121;
  wire popcount24_0c31_core_122;
  wire popcount24_0c31_core_124;
  wire popcount24_0c31_core_125;
  wire popcount24_0c31_core_126;
  wire popcount24_0c31_core_127;
  wire popcount24_0c31_core_128;
  wire popcount24_0c31_core_129_not;
  wire popcount24_0c31_core_130;
  wire popcount24_0c31_core_133;
  wire popcount24_0c31_core_134;
  wire popcount24_0c31_core_135;
  wire popcount24_0c31_core_137;
  wire popcount24_0c31_core_139;
  wire popcount24_0c31_core_140;
  wire popcount24_0c31_core_142;
  wire popcount24_0c31_core_143;
  wire popcount24_0c31_core_145;
  wire popcount24_0c31_core_146;
  wire popcount24_0c31_core_147;
  wire popcount24_0c31_core_148;
  wire popcount24_0c31_core_150;
  wire popcount24_0c31_core_151;
  wire popcount24_0c31_core_152;
  wire popcount24_0c31_core_154;
  wire popcount24_0c31_core_155;
  wire popcount24_0c31_core_158;
  wire popcount24_0c31_core_160;
  wire popcount24_0c31_core_161;
  wire popcount24_0c31_core_163;
  wire popcount24_0c31_core_166;
  wire popcount24_0c31_core_168;
  wire popcount24_0c31_core_169;
  wire popcount24_0c31_core_173;
  wire popcount24_0c31_core_175;
  wire popcount24_0c31_core_176;
  wire popcount24_0c31_core_177;

  assign popcount24_0c31_core_027_not = ~input_a[2];
  assign popcount24_0c31_core_028 = ~input_a[9];
  assign popcount24_0c31_core_030 = ~(input_a[11] & input_a[1]);
  assign popcount24_0c31_core_034 = input_a[8] ^ input_a[9];
  assign popcount24_0c31_core_035 = ~(input_a[20] ^ input_a[4]);
  assign popcount24_0c31_core_037 = ~(input_a[3] | input_a[20]);
  assign popcount24_0c31_core_038 = ~input_a[14];
  assign popcount24_0c31_core_039 = ~(input_a[4] ^ input_a[3]);
  assign popcount24_0c31_core_040 = input_a[16] ^ input_a[3];
  assign popcount24_0c31_core_041 = ~input_a[20];
  assign popcount24_0c31_core_042 = input_a[9] & input_a[7];
  assign popcount24_0c31_core_043_not = ~input_a[2];
  assign popcount24_0c31_core_044 = ~input_a[10];
  assign popcount24_0c31_core_045 = input_a[16] & input_a[15];
  assign popcount24_0c31_core_046 = input_a[0] | input_a[21];
  assign popcount24_0c31_core_047 = input_a[3] & input_a[11];
  assign popcount24_0c31_core_048 = ~(input_a[2] & input_a[16]);
  assign popcount24_0c31_core_053 = ~(input_a[14] & input_a[5]);
  assign popcount24_0c31_core_055_not = ~input_a[16];
  assign popcount24_0c31_core_056 = ~(input_a[7] ^ input_a[11]);
  assign popcount24_0c31_core_058 = ~(input_a[8] & input_a[2]);
  assign popcount24_0c31_core_059_not = ~input_a[5];
  assign popcount24_0c31_core_061 = input_a[14] ^ input_a[3];
  assign popcount24_0c31_core_062 = ~(input_a[8] ^ input_a[2]);
  assign popcount24_0c31_core_065 = ~(input_a[15] & input_a[0]);
  assign popcount24_0c31_core_066_not = ~input_a[17];
  assign popcount24_0c31_core_068 = ~(input_a[16] ^ input_a[13]);
  assign popcount24_0c31_core_069 = input_a[0] ^ input_a[7];
  assign popcount24_0c31_core_072 = ~(input_a[21] ^ input_a[14]);
  assign popcount24_0c31_core_074 = ~input_a[2];
  assign popcount24_0c31_core_076 = ~(input_a[21] | input_a[13]);
  assign popcount24_0c31_core_077 = ~(input_a[0] | input_a[5]);
  assign popcount24_0c31_core_078 = ~(input_a[15] ^ input_a[13]);
  assign popcount24_0c31_core_080 = ~(input_a[23] & input_a[12]);
  assign popcount24_0c31_core_081 = input_a[9] & input_a[3];
  assign popcount24_0c31_core_083 = ~(input_a[0] ^ input_a[20]);
  assign popcount24_0c31_core_084 = input_a[4] | input_a[13];
  assign popcount24_0c31_core_086 = input_a[11] | input_a[19];
  assign popcount24_0c31_core_087 = ~(input_a[3] | input_a[2]);
  assign popcount24_0c31_core_089 = ~(input_a[18] & input_a[7]);
  assign popcount24_0c31_core_090 = input_a[6] & input_a[7];
  assign popcount24_0c31_core_092 = ~(input_a[1] ^ input_a[19]);
  assign popcount24_0c31_core_093 = input_a[9] | input_a[21];
  assign popcount24_0c31_core_094 = ~(input_a[5] | input_a[5]);
  assign popcount24_0c31_core_096 = ~input_a[14];
  assign popcount24_0c31_core_097 = input_a[0] & input_a[1];
  assign popcount24_0c31_core_099 = input_a[11] ^ input_a[19];
  assign popcount24_0c31_core_100 = ~(input_a[17] | input_a[23]);
  assign popcount24_0c31_core_101 = input_a[6] ^ input_a[13];
  assign popcount24_0c31_core_102 = input_a[11] | input_a[23];
  assign popcount24_0c31_core_106 = ~(input_a[17] ^ input_a[13]);
  assign popcount24_0c31_core_112 = input_a[20] & input_a[9];
  assign popcount24_0c31_core_114 = ~input_a[8];
  assign popcount24_0c31_core_115 = ~input_a[7];
  assign popcount24_0c31_core_116 = ~(input_a[23] ^ input_a[8]);
  assign popcount24_0c31_core_117 = ~(input_a[7] | input_a[13]);
  assign popcount24_0c31_core_119 = input_a[8] ^ input_a[0];
  assign popcount24_0c31_core_120 = ~(input_a[15] ^ input_a[14]);
  assign popcount24_0c31_core_121 = ~input_a[1];
  assign popcount24_0c31_core_122 = ~input_a[5];
  assign popcount24_0c31_core_124 = ~(input_a[9] ^ input_a[17]);
  assign popcount24_0c31_core_125 = input_a[20] | input_a[0];
  assign popcount24_0c31_core_126 = ~(input_a[15] | input_a[4]);
  assign popcount24_0c31_core_127 = ~input_a[22];
  assign popcount24_0c31_core_128 = input_a[7] ^ input_a[0];
  assign popcount24_0c31_core_129_not = ~input_a[15];
  assign popcount24_0c31_core_130 = ~(input_a[12] | input_a[23]);
  assign popcount24_0c31_core_133 = ~(input_a[22] & input_a[7]);
  assign popcount24_0c31_core_134 = ~input_a[6];
  assign popcount24_0c31_core_135 = input_a[11] | input_a[8];
  assign popcount24_0c31_core_137 = input_a[9] ^ input_a[2];
  assign popcount24_0c31_core_139 = ~(input_a[23] & input_a[5]);
  assign popcount24_0c31_core_140 = ~(input_a[23] & input_a[3]);
  assign popcount24_0c31_core_142 = ~(input_a[19] | input_a[21]);
  assign popcount24_0c31_core_143 = ~(input_a[0] & input_a[22]);
  assign popcount24_0c31_core_145 = input_a[0] | input_a[19];
  assign popcount24_0c31_core_146 = ~(input_a[6] ^ input_a[1]);
  assign popcount24_0c31_core_147 = ~(input_a[16] & input_a[7]);
  assign popcount24_0c31_core_148 = input_a[8] & input_a[7];
  assign popcount24_0c31_core_150 = input_a[12] & input_a[7];
  assign popcount24_0c31_core_151 = input_a[11] | input_a[22];
  assign popcount24_0c31_core_152 = ~(input_a[8] | input_a[15]);
  assign popcount24_0c31_core_154 = ~(input_a[7] | input_a[3]);
  assign popcount24_0c31_core_155 = input_a[6] & input_a[14];
  assign popcount24_0c31_core_158 = ~input_a[17];
  assign popcount24_0c31_core_160 = input_a[10] & input_a[7];
  assign popcount24_0c31_core_161 = ~(input_a[6] | input_a[18]);
  assign popcount24_0c31_core_163 = input_a[17] & input_a[9];
  assign popcount24_0c31_core_166 = input_a[16] & input_a[7];
  assign popcount24_0c31_core_168 = ~(input_a[16] ^ input_a[8]);
  assign popcount24_0c31_core_169 = input_a[1] ^ input_a[21];
  assign popcount24_0c31_core_173 = input_a[21] & input_a[18];
  assign popcount24_0c31_core_175 = ~(input_a[20] ^ input_a[1]);
  assign popcount24_0c31_core_176 = ~(input_a[15] ^ input_a[1]);
  assign popcount24_0c31_core_177 = ~(input_a[13] | input_a[18]);

  assign popcount24_0c31_out[0] = 1'b0;
  assign popcount24_0c31_out[1] = input_a[20];
  assign popcount24_0c31_out[2] = input_a[5];
  assign popcount24_0c31_out[3] = 1'b0;
  assign popcount24_0c31_out[4] = 1'b1;
endmodule