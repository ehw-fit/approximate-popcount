// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.39114
// WCE=15.0
// EP=0.87048%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_90nk(input [26:0] input_a, output [4:0] popcount27_90nk_out);
  wire popcount27_90nk_core_029;
  wire popcount27_90nk_core_030;
  wire popcount27_90nk_core_032;
  wire popcount27_90nk_core_033;
  wire popcount27_90nk_core_034;
  wire popcount27_90nk_core_035;
  wire popcount27_90nk_core_036;
  wire popcount27_90nk_core_037;
  wire popcount27_90nk_core_039;
  wire popcount27_90nk_core_041_not;
  wire popcount27_90nk_core_043;
  wire popcount27_90nk_core_045_not;
  wire popcount27_90nk_core_049;
  wire popcount27_90nk_core_051;
  wire popcount27_90nk_core_053;
  wire popcount27_90nk_core_054;
  wire popcount27_90nk_core_057;
  wire popcount27_90nk_core_059;
  wire popcount27_90nk_core_060;
  wire popcount27_90nk_core_062;
  wire popcount27_90nk_core_063;
  wire popcount27_90nk_core_065;
  wire popcount27_90nk_core_066;
  wire popcount27_90nk_core_067;
  wire popcount27_90nk_core_069;
  wire popcount27_90nk_core_070;
  wire popcount27_90nk_core_071;
  wire popcount27_90nk_core_074;
  wire popcount27_90nk_core_075;
  wire popcount27_90nk_core_076;
  wire popcount27_90nk_core_077;
  wire popcount27_90nk_core_078;
  wire popcount27_90nk_core_079;
  wire popcount27_90nk_core_080;
  wire popcount27_90nk_core_081;
  wire popcount27_90nk_core_084;
  wire popcount27_90nk_core_085;
  wire popcount27_90nk_core_086;
  wire popcount27_90nk_core_087;
  wire popcount27_90nk_core_088;
  wire popcount27_90nk_core_089;
  wire popcount27_90nk_core_091;
  wire popcount27_90nk_core_093;
  wire popcount27_90nk_core_095;
  wire popcount27_90nk_core_096_not;
  wire popcount27_90nk_core_097;
  wire popcount27_90nk_core_098;
  wire popcount27_90nk_core_099_not;
  wire popcount27_90nk_core_100;
  wire popcount27_90nk_core_101;
  wire popcount27_90nk_core_106;
  wire popcount27_90nk_core_107;
  wire popcount27_90nk_core_108;
  wire popcount27_90nk_core_110;
  wire popcount27_90nk_core_111;
  wire popcount27_90nk_core_112;
  wire popcount27_90nk_core_113;
  wire popcount27_90nk_core_116;
  wire popcount27_90nk_core_117;
  wire popcount27_90nk_core_120;
  wire popcount27_90nk_core_121;
  wire popcount27_90nk_core_122;
  wire popcount27_90nk_core_123;
  wire popcount27_90nk_core_127;
  wire popcount27_90nk_core_130;
  wire popcount27_90nk_core_132;
  wire popcount27_90nk_core_133;
  wire popcount27_90nk_core_134;
  wire popcount27_90nk_core_136;
  wire popcount27_90nk_core_137;
  wire popcount27_90nk_core_139;
  wire popcount27_90nk_core_141;
  wire popcount27_90nk_core_142;
  wire popcount27_90nk_core_143;
  wire popcount27_90nk_core_146;
  wire popcount27_90nk_core_148;
  wire popcount27_90nk_core_149;
  wire popcount27_90nk_core_152;
  wire popcount27_90nk_core_153;
  wire popcount27_90nk_core_155;
  wire popcount27_90nk_core_156;
  wire popcount27_90nk_core_157;
  wire popcount27_90nk_core_158;
  wire popcount27_90nk_core_159;
  wire popcount27_90nk_core_160;
  wire popcount27_90nk_core_161;
  wire popcount27_90nk_core_163;
  wire popcount27_90nk_core_165;
  wire popcount27_90nk_core_166;
  wire popcount27_90nk_core_167;
  wire popcount27_90nk_core_169;
  wire popcount27_90nk_core_171;
  wire popcount27_90nk_core_172;
  wire popcount27_90nk_core_173;
  wire popcount27_90nk_core_174;
  wire popcount27_90nk_core_175_not;
  wire popcount27_90nk_core_177;
  wire popcount27_90nk_core_181;
  wire popcount27_90nk_core_184;
  wire popcount27_90nk_core_187;
  wire popcount27_90nk_core_189;
  wire popcount27_90nk_core_190;
  wire popcount27_90nk_core_192;
  wire popcount27_90nk_core_193;
  wire popcount27_90nk_core_194;
  wire popcount27_90nk_core_195;

  assign popcount27_90nk_core_029 = input_a[18] & input_a[24];
  assign popcount27_90nk_core_030 = input_a[24] | input_a[25];
  assign popcount27_90nk_core_032 = ~(input_a[9] | input_a[8]);
  assign popcount27_90nk_core_033 = ~(input_a[14] ^ input_a[3]);
  assign popcount27_90nk_core_034 = ~(input_a[12] & input_a[10]);
  assign popcount27_90nk_core_035 = input_a[5] | input_a[12];
  assign popcount27_90nk_core_036 = ~(input_a[12] & input_a[5]);
  assign popcount27_90nk_core_037 = input_a[14] | input_a[16];
  assign popcount27_90nk_core_039 = ~input_a[23];
  assign popcount27_90nk_core_041_not = ~input_a[0];
  assign popcount27_90nk_core_043 = ~(input_a[0] ^ input_a[16]);
  assign popcount27_90nk_core_045_not = ~input_a[7];
  assign popcount27_90nk_core_049 = ~(input_a[15] | input_a[25]);
  assign popcount27_90nk_core_051 = ~(input_a[18] | input_a[12]);
  assign popcount27_90nk_core_053 = ~(input_a[20] & input_a[14]);
  assign popcount27_90nk_core_054 = ~(input_a[13] ^ input_a[21]);
  assign popcount27_90nk_core_057 = ~(input_a[26] & input_a[25]);
  assign popcount27_90nk_core_059 = input_a[3] & input_a[9];
  assign popcount27_90nk_core_060 = ~input_a[19];
  assign popcount27_90nk_core_062 = input_a[8] | input_a[6];
  assign popcount27_90nk_core_063 = ~(input_a[10] | input_a[24]);
  assign popcount27_90nk_core_065 = ~(input_a[10] & input_a[25]);
  assign popcount27_90nk_core_066 = ~(input_a[15] ^ input_a[4]);
  assign popcount27_90nk_core_067 = ~(input_a[19] ^ input_a[26]);
  assign popcount27_90nk_core_069 = input_a[19] & input_a[5];
  assign popcount27_90nk_core_070 = input_a[7] ^ input_a[24];
  assign popcount27_90nk_core_071 = ~(input_a[4] & input_a[18]);
  assign popcount27_90nk_core_074 = ~(input_a[20] | input_a[23]);
  assign popcount27_90nk_core_075 = ~input_a[15];
  assign popcount27_90nk_core_076 = ~(input_a[20] & input_a[5]);
  assign popcount27_90nk_core_077 = ~input_a[6];
  assign popcount27_90nk_core_078 = input_a[15] & input_a[21];
  assign popcount27_90nk_core_079 = ~(input_a[11] | input_a[16]);
  assign popcount27_90nk_core_080 = ~(input_a[9] & input_a[20]);
  assign popcount27_90nk_core_081 = input_a[16] & input_a[24];
  assign popcount27_90nk_core_084 = input_a[24] | input_a[5];
  assign popcount27_90nk_core_085 = input_a[10] ^ input_a[4];
  assign popcount27_90nk_core_086 = ~(input_a[10] ^ input_a[10]);
  assign popcount27_90nk_core_087 = input_a[24] | input_a[19];
  assign popcount27_90nk_core_088 = ~input_a[5];
  assign popcount27_90nk_core_089 = ~(input_a[11] ^ input_a[25]);
  assign popcount27_90nk_core_091 = ~input_a[23];
  assign popcount27_90nk_core_093 = ~(input_a[22] ^ input_a[4]);
  assign popcount27_90nk_core_095 = ~(input_a[21] ^ input_a[12]);
  assign popcount27_90nk_core_096_not = ~input_a[14];
  assign popcount27_90nk_core_097 = ~(input_a[3] & input_a[21]);
  assign popcount27_90nk_core_098 = input_a[14] & input_a[14];
  assign popcount27_90nk_core_099_not = ~input_a[23];
  assign popcount27_90nk_core_100 = input_a[4] ^ input_a[0];
  assign popcount27_90nk_core_101 = ~(input_a[7] ^ input_a[6]);
  assign popcount27_90nk_core_106 = ~input_a[2];
  assign popcount27_90nk_core_107 = ~input_a[10];
  assign popcount27_90nk_core_108 = input_a[11] & input_a[24];
  assign popcount27_90nk_core_110 = input_a[5] & input_a[19];
  assign popcount27_90nk_core_111 = ~input_a[14];
  assign popcount27_90nk_core_112 = ~(input_a[7] | input_a[11]);
  assign popcount27_90nk_core_113 = ~(input_a[16] & input_a[20]);
  assign popcount27_90nk_core_116 = input_a[26] | input_a[18];
  assign popcount27_90nk_core_117 = input_a[13] & input_a[20];
  assign popcount27_90nk_core_120 = input_a[8] & input_a[5];
  assign popcount27_90nk_core_121 = input_a[13] ^ input_a[23];
  assign popcount27_90nk_core_122 = ~(input_a[10] ^ input_a[2]);
  assign popcount27_90nk_core_123 = ~input_a[12];
  assign popcount27_90nk_core_127 = input_a[1] & input_a[26];
  assign popcount27_90nk_core_130 = input_a[14] | input_a[20];
  assign popcount27_90nk_core_132 = input_a[23] ^ input_a[0];
  assign popcount27_90nk_core_133 = input_a[12] & input_a[8];
  assign popcount27_90nk_core_134 = input_a[5] & input_a[16];
  assign popcount27_90nk_core_136 = ~(input_a[11] | input_a[25]);
  assign popcount27_90nk_core_137 = input_a[13] & input_a[8];
  assign popcount27_90nk_core_139 = ~input_a[0];
  assign popcount27_90nk_core_141 = ~input_a[14];
  assign popcount27_90nk_core_142 = input_a[20] | input_a[16];
  assign popcount27_90nk_core_143 = input_a[14] & input_a[18];
  assign popcount27_90nk_core_146 = input_a[18] | input_a[2];
  assign popcount27_90nk_core_148 = ~(input_a[10] ^ input_a[5]);
  assign popcount27_90nk_core_149 = input_a[25] & input_a[18];
  assign popcount27_90nk_core_152 = ~(input_a[25] ^ input_a[18]);
  assign popcount27_90nk_core_153 = ~(input_a[8] & input_a[13]);
  assign popcount27_90nk_core_155 = input_a[14] & input_a[8];
  assign popcount27_90nk_core_156 = ~(input_a[8] & input_a[20]);
  assign popcount27_90nk_core_157 = input_a[21] | input_a[19];
  assign popcount27_90nk_core_158 = ~(input_a[24] | input_a[0]);
  assign popcount27_90nk_core_159 = input_a[5] ^ input_a[2];
  assign popcount27_90nk_core_160 = ~(input_a[13] | input_a[3]);
  assign popcount27_90nk_core_161 = input_a[2] & input_a[20];
  assign popcount27_90nk_core_163 = ~(input_a[2] & input_a[22]);
  assign popcount27_90nk_core_165 = ~input_a[22];
  assign popcount27_90nk_core_166 = ~(input_a[23] ^ input_a[3]);
  assign popcount27_90nk_core_167 = ~(input_a[26] ^ input_a[3]);
  assign popcount27_90nk_core_169 = ~(input_a[1] ^ input_a[21]);
  assign popcount27_90nk_core_171 = ~(input_a[25] ^ input_a[14]);
  assign popcount27_90nk_core_172 = ~(input_a[25] ^ input_a[13]);
  assign popcount27_90nk_core_173 = input_a[3] & input_a[22];
  assign popcount27_90nk_core_174 = ~(input_a[12] | input_a[4]);
  assign popcount27_90nk_core_175_not = ~input_a[2];
  assign popcount27_90nk_core_177 = ~(input_a[20] ^ input_a[14]);
  assign popcount27_90nk_core_181 = input_a[12] & input_a[24];
  assign popcount27_90nk_core_184 = ~(input_a[16] | input_a[22]);
  assign popcount27_90nk_core_187 = ~(input_a[18] & input_a[18]);
  assign popcount27_90nk_core_189 = input_a[1] ^ input_a[15];
  assign popcount27_90nk_core_190 = input_a[7] | input_a[24];
  assign popcount27_90nk_core_192 = input_a[17] ^ input_a[23];
  assign popcount27_90nk_core_193 = input_a[18] & input_a[15];
  assign popcount27_90nk_core_194 = input_a[11] & input_a[12];
  assign popcount27_90nk_core_195 = ~(input_a[0] & input_a[25]);

  assign popcount27_90nk_out[0] = 1'b0;
  assign popcount27_90nk_out[1] = 1'b0;
  assign popcount27_90nk_out[2] = 1'b1;
  assign popcount27_90nk_out[3] = 1'b1;
  assign popcount27_90nk_out[4] = 1'b0;
endmodule