// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.6047
// WCE=24.0
// EP=0.971946%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_n50r(input [22:0] input_a, output [4:0] popcount23_n50r_out);
  wire popcount23_n50r_core_025;
  wire popcount23_n50r_core_026;
  wire popcount23_n50r_core_027;
  wire popcount23_n50r_core_028;
  wire popcount23_n50r_core_030;
  wire popcount23_n50r_core_031;
  wire popcount23_n50r_core_034;
  wire popcount23_n50r_core_037;
  wire popcount23_n50r_core_038;
  wire popcount23_n50r_core_040;
  wire popcount23_n50r_core_043;
  wire popcount23_n50r_core_045;
  wire popcount23_n50r_core_046;
  wire popcount23_n50r_core_047;
  wire popcount23_n50r_core_048;
  wire popcount23_n50r_core_049;
  wire popcount23_n50r_core_051;
  wire popcount23_n50r_core_052;
  wire popcount23_n50r_core_053;
  wire popcount23_n50r_core_054;
  wire popcount23_n50r_core_055;
  wire popcount23_n50r_core_057_not;
  wire popcount23_n50r_core_059;
  wire popcount23_n50r_core_060_not;
  wire popcount23_n50r_core_061;
  wire popcount23_n50r_core_067;
  wire popcount23_n50r_core_068;
  wire popcount23_n50r_core_069;
  wire popcount23_n50r_core_070;
  wire popcount23_n50r_core_071_not;
  wire popcount23_n50r_core_072;
  wire popcount23_n50r_core_073;
  wire popcount23_n50r_core_074;
  wire popcount23_n50r_core_077;
  wire popcount23_n50r_core_078;
  wire popcount23_n50r_core_079;
  wire popcount23_n50r_core_080;
  wire popcount23_n50r_core_082_not;
  wire popcount23_n50r_core_083;
  wire popcount23_n50r_core_084;
  wire popcount23_n50r_core_085;
  wire popcount23_n50r_core_088;
  wire popcount23_n50r_core_089;
  wire popcount23_n50r_core_091;
  wire popcount23_n50r_core_092_not;
  wire popcount23_n50r_core_093;
  wire popcount23_n50r_core_094;
  wire popcount23_n50r_core_095;
  wire popcount23_n50r_core_099;
  wire popcount23_n50r_core_101;
  wire popcount23_n50r_core_102;
  wire popcount23_n50r_core_103;
  wire popcount23_n50r_core_104;
  wire popcount23_n50r_core_105;
  wire popcount23_n50r_core_107;
  wire popcount23_n50r_core_110;
  wire popcount23_n50r_core_113;
  wire popcount23_n50r_core_114;
  wire popcount23_n50r_core_115;
  wire popcount23_n50r_core_118;
  wire popcount23_n50r_core_119;
  wire popcount23_n50r_core_122;
  wire popcount23_n50r_core_123;
  wire popcount23_n50r_core_124;
  wire popcount23_n50r_core_125;
  wire popcount23_n50r_core_126;
  wire popcount23_n50r_core_129;
  wire popcount23_n50r_core_130;
  wire popcount23_n50r_core_132;
  wire popcount23_n50r_core_133;
  wire popcount23_n50r_core_134;
  wire popcount23_n50r_core_135;
  wire popcount23_n50r_core_136;
  wire popcount23_n50r_core_137;
  wire popcount23_n50r_core_140;
  wire popcount23_n50r_core_141;
  wire popcount23_n50r_core_143;
  wire popcount23_n50r_core_144;
  wire popcount23_n50r_core_147;
  wire popcount23_n50r_core_153;
  wire popcount23_n50r_core_155;
  wire popcount23_n50r_core_157;
  wire popcount23_n50r_core_160;
  wire popcount23_n50r_core_162;
  wire popcount23_n50r_core_163;
  wire popcount23_n50r_core_165;
  wire popcount23_n50r_core_166;
  wire popcount23_n50r_core_168;

  assign popcount23_n50r_core_025 = ~(input_a[15] ^ input_a[20]);
  assign popcount23_n50r_core_026 = input_a[19] & input_a[16];
  assign popcount23_n50r_core_027 = input_a[19] ^ input_a[15];
  assign popcount23_n50r_core_028 = ~(input_a[10] | input_a[4]);
  assign popcount23_n50r_core_030 = ~(input_a[4] | input_a[6]);
  assign popcount23_n50r_core_031 = ~(input_a[13] | input_a[20]);
  assign popcount23_n50r_core_034 = input_a[19] ^ input_a[2];
  assign popcount23_n50r_core_037 = ~(input_a[7] ^ input_a[10]);
  assign popcount23_n50r_core_038 = ~input_a[16];
  assign popcount23_n50r_core_040 = ~input_a[19];
  assign popcount23_n50r_core_043 = input_a[7] ^ input_a[15];
  assign popcount23_n50r_core_045 = ~input_a[18];
  assign popcount23_n50r_core_046 = ~(input_a[3] ^ input_a[21]);
  assign popcount23_n50r_core_047 = input_a[8] | input_a[14];
  assign popcount23_n50r_core_048 = ~(input_a[20] ^ input_a[12]);
  assign popcount23_n50r_core_049 = ~input_a[14];
  assign popcount23_n50r_core_051 = ~(input_a[9] & input_a[19]);
  assign popcount23_n50r_core_052 = input_a[11] ^ input_a[14];
  assign popcount23_n50r_core_053 = ~(input_a[5] ^ input_a[19]);
  assign popcount23_n50r_core_054 = ~(input_a[7] ^ input_a[19]);
  assign popcount23_n50r_core_055 = ~(input_a[18] | input_a[20]);
  assign popcount23_n50r_core_057_not = ~input_a[5];
  assign popcount23_n50r_core_059 = ~input_a[9];
  assign popcount23_n50r_core_060_not = ~input_a[16];
  assign popcount23_n50r_core_061 = input_a[2] & input_a[13];
  assign popcount23_n50r_core_067 = input_a[8] | input_a[13];
  assign popcount23_n50r_core_068 = ~input_a[18];
  assign popcount23_n50r_core_069 = ~(input_a[10] ^ input_a[4]);
  assign popcount23_n50r_core_070 = input_a[11] | input_a[7];
  assign popcount23_n50r_core_071_not = ~input_a[17];
  assign popcount23_n50r_core_072 = ~(input_a[13] | input_a[1]);
  assign popcount23_n50r_core_073 = input_a[19] | input_a[6];
  assign popcount23_n50r_core_074 = input_a[21] ^ input_a[22];
  assign popcount23_n50r_core_077 = input_a[9] & input_a[16];
  assign popcount23_n50r_core_078 = ~(input_a[5] | input_a[8]);
  assign popcount23_n50r_core_079 = ~input_a[17];
  assign popcount23_n50r_core_080 = input_a[7] & input_a[1];
  assign popcount23_n50r_core_082_not = ~input_a[22];
  assign popcount23_n50r_core_083 = ~input_a[22];
  assign popcount23_n50r_core_084 = ~input_a[15];
  assign popcount23_n50r_core_085 = input_a[8] & input_a[14];
  assign popcount23_n50r_core_088 = input_a[4] & input_a[19];
  assign popcount23_n50r_core_089 = ~input_a[2];
  assign popcount23_n50r_core_091 = ~input_a[18];
  assign popcount23_n50r_core_092_not = ~input_a[9];
  assign popcount23_n50r_core_093 = ~(input_a[17] ^ input_a[10]);
  assign popcount23_n50r_core_094 = input_a[8] & input_a[21];
  assign popcount23_n50r_core_095 = input_a[14] | input_a[20];
  assign popcount23_n50r_core_099 = ~(input_a[19] ^ input_a[2]);
  assign popcount23_n50r_core_101 = input_a[1] | input_a[15];
  assign popcount23_n50r_core_102 = ~(input_a[6] ^ input_a[13]);
  assign popcount23_n50r_core_103 = input_a[0] & input_a[15];
  assign popcount23_n50r_core_104 = input_a[0] & input_a[9];
  assign popcount23_n50r_core_105 = ~input_a[2];
  assign popcount23_n50r_core_107 = ~input_a[3];
  assign popcount23_n50r_core_110 = ~input_a[15];
  assign popcount23_n50r_core_113 = ~(input_a[16] | input_a[8]);
  assign popcount23_n50r_core_114 = ~(input_a[4] & input_a[17]);
  assign popcount23_n50r_core_115 = ~(input_a[5] | input_a[6]);
  assign popcount23_n50r_core_118 = ~input_a[15];
  assign popcount23_n50r_core_119 = input_a[20] ^ input_a[21];
  assign popcount23_n50r_core_122 = ~input_a[17];
  assign popcount23_n50r_core_123 = ~(input_a[11] ^ input_a[19]);
  assign popcount23_n50r_core_124 = input_a[20] ^ input_a[11];
  assign popcount23_n50r_core_125 = ~(input_a[13] & input_a[22]);
  assign popcount23_n50r_core_126 = input_a[14] & input_a[18];
  assign popcount23_n50r_core_129 = input_a[15] & input_a[2];
  assign popcount23_n50r_core_130 = input_a[20] & input_a[9];
  assign popcount23_n50r_core_132 = input_a[22] ^ input_a[13];
  assign popcount23_n50r_core_133 = ~input_a[14];
  assign popcount23_n50r_core_134 = ~input_a[18];
  assign popcount23_n50r_core_135 = ~(input_a[5] & input_a[17]);
  assign popcount23_n50r_core_136 = ~(input_a[9] & input_a[15]);
  assign popcount23_n50r_core_137 = input_a[13] | input_a[1];
  assign popcount23_n50r_core_140 = ~input_a[3];
  assign popcount23_n50r_core_141 = input_a[8] | input_a[18];
  assign popcount23_n50r_core_143 = ~(input_a[13] | input_a[0]);
  assign popcount23_n50r_core_144 = ~(input_a[2] | input_a[0]);
  assign popcount23_n50r_core_147 = ~(input_a[5] ^ input_a[8]);
  assign popcount23_n50r_core_153 = ~(input_a[2] | input_a[9]);
  assign popcount23_n50r_core_155 = input_a[19] ^ input_a[15];
  assign popcount23_n50r_core_157 = ~(input_a[20] ^ input_a[0]);
  assign popcount23_n50r_core_160 = ~(input_a[8] | input_a[13]);
  assign popcount23_n50r_core_162 = input_a[17] | input_a[18];
  assign popcount23_n50r_core_163 = ~input_a[9];
  assign popcount23_n50r_core_165 = ~input_a[1];
  assign popcount23_n50r_core_166 = input_a[5] & input_a[1];
  assign popcount23_n50r_core_168 = input_a[1] ^ input_a[10];

  assign popcount23_n50r_out[0] = 1'b0;
  assign popcount23_n50r_out[1] = 1'b0;
  assign popcount23_n50r_out[2] = 1'b0;
  assign popcount23_n50r_out[3] = input_a[19];
  assign popcount23_n50r_out[4] = input_a[2];
endmodule