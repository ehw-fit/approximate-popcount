// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.59546
// WCE=19.0
// EP=0.927471%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_9ybe(input [22:0] input_a, output [4:0] popcount23_9ybe_out);
  wire popcount23_9ybe_core_026;
  wire popcount23_9ybe_core_031;
  wire popcount23_9ybe_core_032;
  wire popcount23_9ybe_core_033;
  wire popcount23_9ybe_core_034;
  wire popcount23_9ybe_core_040;
  wire popcount23_9ybe_core_041;
  wire popcount23_9ybe_core_042;
  wire popcount23_9ybe_core_044;
  wire popcount23_9ybe_core_045;
  wire popcount23_9ybe_core_047;
  wire popcount23_9ybe_core_050;
  wire popcount23_9ybe_core_051;
  wire popcount23_9ybe_core_053;
  wire popcount23_9ybe_core_054;
  wire popcount23_9ybe_core_058;
  wire popcount23_9ybe_core_062;
  wire popcount23_9ybe_core_064;
  wire popcount23_9ybe_core_065;
  wire popcount23_9ybe_core_066;
  wire popcount23_9ybe_core_067;
  wire popcount23_9ybe_core_068;
  wire popcount23_9ybe_core_069;
  wire popcount23_9ybe_core_070;
  wire popcount23_9ybe_core_072;
  wire popcount23_9ybe_core_074;
  wire popcount23_9ybe_core_075;
  wire popcount23_9ybe_core_076_not;
  wire popcount23_9ybe_core_077;
  wire popcount23_9ybe_core_079;
  wire popcount23_9ybe_core_081;
  wire popcount23_9ybe_core_082_not;
  wire popcount23_9ybe_core_084;
  wire popcount23_9ybe_core_085;
  wire popcount23_9ybe_core_087;
  wire popcount23_9ybe_core_089;
  wire popcount23_9ybe_core_090;
  wire popcount23_9ybe_core_091;
  wire popcount23_9ybe_core_092;
  wire popcount23_9ybe_core_096;
  wire popcount23_9ybe_core_098;
  wire popcount23_9ybe_core_101;
  wire popcount23_9ybe_core_102;
  wire popcount23_9ybe_core_103;
  wire popcount23_9ybe_core_105;
  wire popcount23_9ybe_core_107;
  wire popcount23_9ybe_core_108;
  wire popcount23_9ybe_core_109;
  wire popcount23_9ybe_core_112;
  wire popcount23_9ybe_core_113;
  wire popcount23_9ybe_core_114;
  wire popcount23_9ybe_core_115;
  wire popcount23_9ybe_core_117;
  wire popcount23_9ybe_core_118;
  wire popcount23_9ybe_core_119;
  wire popcount23_9ybe_core_120;
  wire popcount23_9ybe_core_122_not;
  wire popcount23_9ybe_core_124;
  wire popcount23_9ybe_core_127;
  wire popcount23_9ybe_core_128;
  wire popcount23_9ybe_core_130;
  wire popcount23_9ybe_core_132;
  wire popcount23_9ybe_core_133;
  wire popcount23_9ybe_core_134;
  wire popcount23_9ybe_core_135;
  wire popcount23_9ybe_core_136;
  wire popcount23_9ybe_core_137;
  wire popcount23_9ybe_core_138;
  wire popcount23_9ybe_core_139;
  wire popcount23_9ybe_core_140;
  wire popcount23_9ybe_core_143;
  wire popcount23_9ybe_core_144;
  wire popcount23_9ybe_core_145;
  wire popcount23_9ybe_core_146;
  wire popcount23_9ybe_core_148;
  wire popcount23_9ybe_core_149;
  wire popcount23_9ybe_core_150;
  wire popcount23_9ybe_core_151;
  wire popcount23_9ybe_core_152;
  wire popcount23_9ybe_core_153;
  wire popcount23_9ybe_core_155;
  wire popcount23_9ybe_core_160;
  wire popcount23_9ybe_core_161;
  wire popcount23_9ybe_core_163;
  wire popcount23_9ybe_core_165;
  wire popcount23_9ybe_core_168;

  assign popcount23_9ybe_core_026 = input_a[0] & input_a[13];
  assign popcount23_9ybe_core_031 = ~(input_a[22] | input_a[20]);
  assign popcount23_9ybe_core_032 = input_a[8] ^ input_a[4];
  assign popcount23_9ybe_core_033 = ~(input_a[8] & input_a[11]);
  assign popcount23_9ybe_core_034 = ~(input_a[12] ^ input_a[16]);
  assign popcount23_9ybe_core_040 = input_a[18] & input_a[22];
  assign popcount23_9ybe_core_041 = input_a[10] & input_a[10];
  assign popcount23_9ybe_core_042 = input_a[2] ^ input_a[19];
  assign popcount23_9ybe_core_044 = ~(input_a[4] & input_a[13]);
  assign popcount23_9ybe_core_045 = input_a[21] & input_a[2];
  assign popcount23_9ybe_core_047 = ~(input_a[8] | input_a[16]);
  assign popcount23_9ybe_core_050 = ~(input_a[21] | input_a[16]);
  assign popcount23_9ybe_core_051 = ~(input_a[10] & input_a[16]);
  assign popcount23_9ybe_core_053 = ~(input_a[8] ^ input_a[14]);
  assign popcount23_9ybe_core_054 = ~(input_a[13] | input_a[22]);
  assign popcount23_9ybe_core_058 = input_a[5] & input_a[15];
  assign popcount23_9ybe_core_062 = ~(input_a[15] | input_a[17]);
  assign popcount23_9ybe_core_064 = ~input_a[11];
  assign popcount23_9ybe_core_065 = ~input_a[6];
  assign popcount23_9ybe_core_066 = ~(input_a[18] ^ input_a[13]);
  assign popcount23_9ybe_core_067 = ~(input_a[7] ^ input_a[19]);
  assign popcount23_9ybe_core_068 = input_a[21] ^ input_a[2];
  assign popcount23_9ybe_core_069 = ~(input_a[7] | input_a[0]);
  assign popcount23_9ybe_core_070 = ~(input_a[11] | input_a[17]);
  assign popcount23_9ybe_core_072 = input_a[4] & input_a[8];
  assign popcount23_9ybe_core_074 = input_a[7] & input_a[19];
  assign popcount23_9ybe_core_075 = input_a[16] | input_a[14];
  assign popcount23_9ybe_core_076_not = ~input_a[16];
  assign popcount23_9ybe_core_077 = ~(input_a[22] | input_a[3]);
  assign popcount23_9ybe_core_079 = ~input_a[16];
  assign popcount23_9ybe_core_081 = ~(input_a[4] | input_a[9]);
  assign popcount23_9ybe_core_082_not = ~input_a[20];
  assign popcount23_9ybe_core_084 = ~input_a[9];
  assign popcount23_9ybe_core_085 = ~(input_a[22] | input_a[4]);
  assign popcount23_9ybe_core_087 = input_a[22] | input_a[8];
  assign popcount23_9ybe_core_089 = ~(input_a[3] & input_a[12]);
  assign popcount23_9ybe_core_090 = ~(input_a[10] ^ input_a[21]);
  assign popcount23_9ybe_core_091 = input_a[2] & input_a[9];
  assign popcount23_9ybe_core_092 = ~(input_a[5] & input_a[14]);
  assign popcount23_9ybe_core_096 = input_a[5] | input_a[3];
  assign popcount23_9ybe_core_098 = input_a[11] & input_a[19];
  assign popcount23_9ybe_core_101 = input_a[21] & input_a[7];
  assign popcount23_9ybe_core_102 = ~input_a[16];
  assign popcount23_9ybe_core_103 = ~(input_a[7] & input_a[6]);
  assign popcount23_9ybe_core_105 = ~(input_a[7] & input_a[8]);
  assign popcount23_9ybe_core_107 = ~(input_a[19] | input_a[10]);
  assign popcount23_9ybe_core_108 = input_a[3] | input_a[17];
  assign popcount23_9ybe_core_109 = ~(input_a[1] | input_a[15]);
  assign popcount23_9ybe_core_112 = input_a[12] ^ input_a[20];
  assign popcount23_9ybe_core_113 = input_a[6] ^ input_a[17];
  assign popcount23_9ybe_core_114 = input_a[11] ^ input_a[10];
  assign popcount23_9ybe_core_115 = ~(input_a[6] | input_a[9]);
  assign popcount23_9ybe_core_117 = input_a[20] ^ input_a[16];
  assign popcount23_9ybe_core_118 = input_a[20] | input_a[22];
  assign popcount23_9ybe_core_119 = input_a[15] & input_a[17];
  assign popcount23_9ybe_core_120 = input_a[20] ^ input_a[14];
  assign popcount23_9ybe_core_122_not = ~input_a[18];
  assign popcount23_9ybe_core_124 = ~(input_a[21] | input_a[20]);
  assign popcount23_9ybe_core_127 = input_a[6] ^ input_a[8];
  assign popcount23_9ybe_core_128 = input_a[11] | input_a[8];
  assign popcount23_9ybe_core_130 = input_a[15] ^ input_a[5];
  assign popcount23_9ybe_core_132 = input_a[19] | input_a[3];
  assign popcount23_9ybe_core_133 = input_a[7] ^ input_a[21];
  assign popcount23_9ybe_core_134 = ~(input_a[8] | input_a[14]);
  assign popcount23_9ybe_core_135 = input_a[17] ^ input_a[11];
  assign popcount23_9ybe_core_136 = input_a[10] & input_a[6];
  assign popcount23_9ybe_core_137 = ~(input_a[3] ^ input_a[15]);
  assign popcount23_9ybe_core_138 = ~input_a[7];
  assign popcount23_9ybe_core_139 = ~(input_a[17] | input_a[6]);
  assign popcount23_9ybe_core_140 = input_a[14] | input_a[16];
  assign popcount23_9ybe_core_143 = input_a[20] & input_a[4];
  assign popcount23_9ybe_core_144 = ~(input_a[22] & input_a[15]);
  assign popcount23_9ybe_core_145 = input_a[1] ^ input_a[14];
  assign popcount23_9ybe_core_146 = input_a[18] & input_a[20];
  assign popcount23_9ybe_core_148 = ~(input_a[8] | input_a[8]);
  assign popcount23_9ybe_core_149 = input_a[1] ^ input_a[6];
  assign popcount23_9ybe_core_150 = ~input_a[9];
  assign popcount23_9ybe_core_151 = ~(input_a[14] | input_a[19]);
  assign popcount23_9ybe_core_152 = ~(input_a[9] | input_a[7]);
  assign popcount23_9ybe_core_153 = ~(input_a[21] ^ input_a[15]);
  assign popcount23_9ybe_core_155 = input_a[11] | input_a[0];
  assign popcount23_9ybe_core_160 = ~(input_a[2] | input_a[21]);
  assign popcount23_9ybe_core_161 = input_a[19] & input_a[17];
  assign popcount23_9ybe_core_163 = input_a[2] ^ input_a[10];
  assign popcount23_9ybe_core_165 = input_a[1] & input_a[21];
  assign popcount23_9ybe_core_168 = ~input_a[10];

  assign popcount23_9ybe_out[0] = 1'b0;
  assign popcount23_9ybe_out[1] = 1'b1;
  assign popcount23_9ybe_out[2] = input_a[1];
  assign popcount23_9ybe_out[3] = input_a[14];
  assign popcount23_9ybe_out[4] = 1'b0;
endmodule