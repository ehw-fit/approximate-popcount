// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.97148
// WCE=17.0
// EP=0.898831%
// Printed PDK parameters:
//  Area=856340.0
//  Delay=2618200.0
//  Power=31251.0

module popcount30_iw31(input [29:0] input_a, output [4:0] popcount30_iw31_out);
  wire popcount30_iw31_core_032;
  wire popcount30_iw31_core_034;
  wire popcount30_iw31_core_035_not;
  wire popcount30_iw31_core_036;
  wire popcount30_iw31_core_038_not;
  wire popcount30_iw31_core_040;
  wire popcount30_iw31_core_042;
  wire popcount30_iw31_core_043;
  wire popcount30_iw31_core_044_not;
  wire popcount30_iw31_core_046;
  wire popcount30_iw31_core_047;
  wire popcount30_iw31_core_048;
  wire popcount30_iw31_core_049;
  wire popcount30_iw31_core_050;
  wire popcount30_iw31_core_052;
  wire popcount30_iw31_core_053;
  wire popcount30_iw31_core_054;
  wire popcount30_iw31_core_056;
  wire popcount30_iw31_core_059;
  wire popcount30_iw31_core_060;
  wire popcount30_iw31_core_061;
  wire popcount30_iw31_core_062;
  wire popcount30_iw31_core_063;
  wire popcount30_iw31_core_064;
  wire popcount30_iw31_core_066;
  wire popcount30_iw31_core_067;
  wire popcount30_iw31_core_069;
  wire popcount30_iw31_core_070;
  wire popcount30_iw31_core_071_not;
  wire popcount30_iw31_core_072;
  wire popcount30_iw31_core_073;
  wire popcount30_iw31_core_074;
  wire popcount30_iw31_core_075;
  wire popcount30_iw31_core_078;
  wire popcount30_iw31_core_081;
  wire popcount30_iw31_core_082;
  wire popcount30_iw31_core_083;
  wire popcount30_iw31_core_084;
  wire popcount30_iw31_core_085;
  wire popcount30_iw31_core_086;
  wire popcount30_iw31_core_087;
  wire popcount30_iw31_core_088;
  wire popcount30_iw31_core_091;
  wire popcount30_iw31_core_092;
  wire popcount30_iw31_core_096;
  wire popcount30_iw31_core_097;
  wire popcount30_iw31_core_098;
  wire popcount30_iw31_core_099;
  wire popcount30_iw31_core_100;
  wire popcount30_iw31_core_107;
  wire popcount30_iw31_core_108;
  wire popcount30_iw31_core_109;
  wire popcount30_iw31_core_110;
  wire popcount30_iw31_core_112;
  wire popcount30_iw31_core_115;
  wire popcount30_iw31_core_116;
  wire popcount30_iw31_core_118;
  wire popcount30_iw31_core_120;
  wire popcount30_iw31_core_121;
  wire popcount30_iw31_core_122;
  wire popcount30_iw31_core_124;
  wire popcount30_iw31_core_125;
  wire popcount30_iw31_core_126;
  wire popcount30_iw31_core_128;
  wire popcount30_iw31_core_130;
  wire popcount30_iw31_core_131;
  wire popcount30_iw31_core_132;
  wire popcount30_iw31_core_135;
  wire popcount30_iw31_core_136;
  wire popcount30_iw31_core_139;
  wire popcount30_iw31_core_140;
  wire popcount30_iw31_core_142;
  wire popcount30_iw31_core_143;
  wire popcount30_iw31_core_145;
  wire popcount30_iw31_core_146;
  wire popcount30_iw31_core_147;
  wire popcount30_iw31_core_148;
  wire popcount30_iw31_core_149;
  wire popcount30_iw31_core_150;
  wire popcount30_iw31_core_152;
  wire popcount30_iw31_core_153;
  wire popcount30_iw31_core_154;
  wire popcount30_iw31_core_155;
  wire popcount30_iw31_core_157;
  wire popcount30_iw31_core_158;
  wire popcount30_iw31_core_159;
  wire popcount30_iw31_core_160;
  wire popcount30_iw31_core_161;
  wire popcount30_iw31_core_162;
  wire popcount30_iw31_core_164;
  wire popcount30_iw31_core_167;
  wire popcount30_iw31_core_170;
  wire popcount30_iw31_core_171;
  wire popcount30_iw31_core_172;
  wire popcount30_iw31_core_173_not;
  wire popcount30_iw31_core_174;
  wire popcount30_iw31_core_175;
  wire popcount30_iw31_core_176;
  wire popcount30_iw31_core_180;
  wire popcount30_iw31_core_181;
  wire popcount30_iw31_core_182;
  wire popcount30_iw31_core_183;
  wire popcount30_iw31_core_184;
  wire popcount30_iw31_core_186;
  wire popcount30_iw31_core_188;
  wire popcount30_iw31_core_189;
  wire popcount30_iw31_core_193;
  wire popcount30_iw31_core_196;
  wire popcount30_iw31_core_197;
  wire popcount30_iw31_core_201;
  wire popcount30_iw31_core_202;
  wire popcount30_iw31_core_204;
  wire popcount30_iw31_core_205;
  wire popcount30_iw31_core_206;
  wire popcount30_iw31_core_207;
  wire popcount30_iw31_core_208_not;
  wire popcount30_iw31_core_209;
  wire popcount30_iw31_core_210;
  wire popcount30_iw31_core_211;
  wire popcount30_iw31_core_212;
  wire popcount30_iw31_core_213;

  assign popcount30_iw31_core_032 = ~(input_a[19] | input_a[13]);
  assign popcount30_iw31_core_034 = ~input_a[7];
  assign popcount30_iw31_core_035_not = ~input_a[15];
  assign popcount30_iw31_core_036 = ~(input_a[25] | input_a[28]);
  assign popcount30_iw31_core_038_not = ~input_a[0];
  assign popcount30_iw31_core_040 = input_a[17] | input_a[28];
  assign popcount30_iw31_core_042 = input_a[4] | input_a[13];
  assign popcount30_iw31_core_043 = input_a[19] & input_a[20];
  assign popcount30_iw31_core_044_not = ~input_a[15];
  assign popcount30_iw31_core_046 = input_a[19] ^ input_a[26];
  assign popcount30_iw31_core_047 = input_a[16] & input_a[23];
  assign popcount30_iw31_core_048 = ~(input_a[29] & input_a[19]);
  assign popcount30_iw31_core_049 = input_a[27] ^ input_a[10];
  assign popcount30_iw31_core_050 = ~input_a[17];
  assign popcount30_iw31_core_052 = input_a[11] & input_a[18];
  assign popcount30_iw31_core_053 = input_a[14] & input_a[23];
  assign popcount30_iw31_core_054 = ~input_a[9];
  assign popcount30_iw31_core_056 = ~input_a[24];
  assign popcount30_iw31_core_059 = ~(input_a[6] | input_a[23]);
  assign popcount30_iw31_core_060 = input_a[3] | input_a[7];
  assign popcount30_iw31_core_061 = ~(input_a[8] & input_a[17]);
  assign popcount30_iw31_core_062 = input_a[27] & input_a[7];
  assign popcount30_iw31_core_063 = input_a[8] & input_a[27];
  assign popcount30_iw31_core_064 = ~(input_a[18] ^ input_a[15]);
  assign popcount30_iw31_core_066 = input_a[11] & input_a[15];
  assign popcount30_iw31_core_067 = ~(input_a[6] & input_a[24]);
  assign popcount30_iw31_core_069 = input_a[10] | input_a[0];
  assign popcount30_iw31_core_070 = ~(input_a[14] & input_a[20]);
  assign popcount30_iw31_core_071_not = ~input_a[23];
  assign popcount30_iw31_core_072 = ~(input_a[10] ^ input_a[28]);
  assign popcount30_iw31_core_073 = ~input_a[24];
  assign popcount30_iw31_core_074 = ~(input_a[27] ^ input_a[3]);
  assign popcount30_iw31_core_075 = input_a[5] | input_a[16];
  assign popcount30_iw31_core_078 = input_a[10] | input_a[5];
  assign popcount30_iw31_core_081 = ~(input_a[22] ^ input_a[22]);
  assign popcount30_iw31_core_082 = ~(input_a[22] & input_a[9]);
  assign popcount30_iw31_core_083 = ~(input_a[29] | input_a[17]);
  assign popcount30_iw31_core_084 = ~(input_a[15] & input_a[28]);
  assign popcount30_iw31_core_085 = input_a[10] | input_a[3];
  assign popcount30_iw31_core_086 = input_a[6] | input_a[17];
  assign popcount30_iw31_core_087 = ~(input_a[1] | input_a[12]);
  assign popcount30_iw31_core_088 = ~(input_a[17] & input_a[12]);
  assign popcount30_iw31_core_091 = input_a[7] | input_a[15];
  assign popcount30_iw31_core_092 = ~(input_a[5] & input_a[25]);
  assign popcount30_iw31_core_096 = input_a[9] ^ input_a[9];
  assign popcount30_iw31_core_097 = input_a[0] & input_a[2];
  assign popcount30_iw31_core_098 = input_a[6] ^ input_a[7];
  assign popcount30_iw31_core_099 = input_a[28] ^ input_a[1];
  assign popcount30_iw31_core_100 = ~(input_a[29] | input_a[9]);
  assign popcount30_iw31_core_107 = ~(input_a[27] & input_a[26]);
  assign popcount30_iw31_core_108 = ~(input_a[28] & input_a[18]);
  assign popcount30_iw31_core_109 = input_a[0] | input_a[6];
  assign popcount30_iw31_core_110 = input_a[5] & input_a[24];
  assign popcount30_iw31_core_112 = input_a[18] ^ input_a[20];
  assign popcount30_iw31_core_115 = ~(input_a[16] | input_a[2]);
  assign popcount30_iw31_core_116 = ~(input_a[27] | input_a[25]);
  assign popcount30_iw31_core_118 = ~(input_a[5] ^ input_a[12]);
  assign popcount30_iw31_core_120 = ~input_a[7];
  assign popcount30_iw31_core_121 = ~input_a[14];
  assign popcount30_iw31_core_122 = input_a[24] & input_a[29];
  assign popcount30_iw31_core_124 = ~(input_a[22] | input_a[3]);
  assign popcount30_iw31_core_125 = input_a[2] & input_a[1];
  assign popcount30_iw31_core_126 = ~input_a[23];
  assign popcount30_iw31_core_128 = input_a[14] & input_a[20];
  assign popcount30_iw31_core_130 = ~(input_a[0] | input_a[10]);
  assign popcount30_iw31_core_131 = ~(input_a[15] | input_a[8]);
  assign popcount30_iw31_core_132 = ~input_a[11];
  assign popcount30_iw31_core_135 = ~(input_a[25] & input_a[11]);
  assign popcount30_iw31_core_136 = ~(input_a[21] & input_a[14]);
  assign popcount30_iw31_core_139 = input_a[7] & input_a[16];
  assign popcount30_iw31_core_140 = ~(input_a[19] | input_a[27]);
  assign popcount30_iw31_core_142 = ~(input_a[16] & input_a[1]);
  assign popcount30_iw31_core_143 = input_a[24] | input_a[27];
  assign popcount30_iw31_core_145 = ~(input_a[6] | input_a[4]);
  assign popcount30_iw31_core_146 = input_a[13] | input_a[12];
  assign popcount30_iw31_core_147 = ~(input_a[20] ^ input_a[13]);
  assign popcount30_iw31_core_148 = ~(input_a[8] | input_a[29]);
  assign popcount30_iw31_core_149 = input_a[8] | input_a[23];
  assign popcount30_iw31_core_150 = ~(input_a[23] ^ input_a[12]);
  assign popcount30_iw31_core_152 = ~(input_a[26] & input_a[20]);
  assign popcount30_iw31_core_153 = input_a[11] | input_a[4];
  assign popcount30_iw31_core_154 = input_a[21] & input_a[10];
  assign popcount30_iw31_core_155 = ~(input_a[9] | input_a[24]);
  assign popcount30_iw31_core_157 = input_a[12] | input_a[26];
  assign popcount30_iw31_core_158 = ~(input_a[7] & input_a[15]);
  assign popcount30_iw31_core_159 = ~(input_a[28] ^ input_a[24]);
  assign popcount30_iw31_core_160 = ~(input_a[3] ^ input_a[9]);
  assign popcount30_iw31_core_161 = ~(input_a[6] | input_a[3]);
  assign popcount30_iw31_core_162 = ~(input_a[22] ^ input_a[27]);
  assign popcount30_iw31_core_164 = ~(input_a[24] & input_a[21]);
  assign popcount30_iw31_core_167 = ~input_a[13];
  assign popcount30_iw31_core_170 = ~(input_a[19] & input_a[22]);
  assign popcount30_iw31_core_171 = ~input_a[21];
  assign popcount30_iw31_core_172 = ~(input_a[17] & input_a[0]);
  assign popcount30_iw31_core_173_not = ~input_a[4];
  assign popcount30_iw31_core_174 = ~input_a[24];
  assign popcount30_iw31_core_175 = ~(input_a[23] | input_a[17]);
  assign popcount30_iw31_core_176 = ~(input_a[29] & input_a[22]);
  assign popcount30_iw31_core_180 = input_a[11] ^ input_a[19];
  assign popcount30_iw31_core_181 = ~(input_a[10] & input_a[16]);
  assign popcount30_iw31_core_182 = ~(input_a[20] & input_a[7]);
  assign popcount30_iw31_core_183 = input_a[28] & input_a[25];
  assign popcount30_iw31_core_184 = ~input_a[1];
  assign popcount30_iw31_core_186 = ~(input_a[11] & input_a[3]);
  assign popcount30_iw31_core_188 = input_a[11] | input_a[22];
  assign popcount30_iw31_core_189 = input_a[28] & input_a[29];
  assign popcount30_iw31_core_193 = input_a[19] & input_a[22];
  assign popcount30_iw31_core_196 = ~(input_a[23] ^ input_a[28]);
  assign popcount30_iw31_core_197 = ~input_a[16];
  assign popcount30_iw31_core_201 = ~(input_a[11] | input_a[26]);
  assign popcount30_iw31_core_202 = popcount30_iw31_core_056 & input_a[16];
  assign popcount30_iw31_core_204 = ~input_a[24];
  assign popcount30_iw31_core_205 = ~(input_a[16] | input_a[24]);
  assign popcount30_iw31_core_206 = popcount30_iw31_core_204 ^ popcount30_iw31_core_202;
  assign popcount30_iw31_core_207 = ~input_a[24];
  assign popcount30_iw31_core_208_not = ~input_a[29];
  assign popcount30_iw31_core_209 = ~(input_a[22] | input_a[14]);
  assign popcount30_iw31_core_210 = ~input_a[20];
  assign popcount30_iw31_core_211 = input_a[16] | input_a[24];
  assign popcount30_iw31_core_212 = input_a[4] | input_a[0];
  assign popcount30_iw31_core_213 = ~(input_a[27] & input_a[10]);

  assign popcount30_iw31_out[0] = input_a[14];
  assign popcount30_iw31_out[1] = popcount30_iw31_core_204;
  assign popcount30_iw31_out[2] = 1'b0;
  assign popcount30_iw31_out[3] = popcount30_iw31_core_206;
  assign popcount30_iw31_out[4] = popcount30_iw31_core_211;
endmodule