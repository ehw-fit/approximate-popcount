// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=10.0243
// WCE=30.0
// EP=0.99045%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_eqge(input [29:0] input_a, output [4:0] popcount30_eqge_out);
  wire popcount30_eqge_core_032;
  wire popcount30_eqge_core_034;
  wire popcount30_eqge_core_035;
  wire popcount30_eqge_core_036;
  wire popcount30_eqge_core_037;
  wire popcount30_eqge_core_038;
  wire popcount30_eqge_core_040;
  wire popcount30_eqge_core_041;
  wire popcount30_eqge_core_042;
  wire popcount30_eqge_core_045;
  wire popcount30_eqge_core_046;
  wire popcount30_eqge_core_048;
  wire popcount30_eqge_core_049;
  wire popcount30_eqge_core_051;
  wire popcount30_eqge_core_052;
  wire popcount30_eqge_core_053;
  wire popcount30_eqge_core_054;
  wire popcount30_eqge_core_056;
  wire popcount30_eqge_core_057;
  wire popcount30_eqge_core_058;
  wire popcount30_eqge_core_059_not;
  wire popcount30_eqge_core_061;
  wire popcount30_eqge_core_063;
  wire popcount30_eqge_core_064;
  wire popcount30_eqge_core_065;
  wire popcount30_eqge_core_070;
  wire popcount30_eqge_core_073;
  wire popcount30_eqge_core_074;
  wire popcount30_eqge_core_075;
  wire popcount30_eqge_core_076;
  wire popcount30_eqge_core_077;
  wire popcount30_eqge_core_080;
  wire popcount30_eqge_core_084;
  wire popcount30_eqge_core_086;
  wire popcount30_eqge_core_088;
  wire popcount30_eqge_core_090;
  wire popcount30_eqge_core_091;
  wire popcount30_eqge_core_092;
  wire popcount30_eqge_core_093;
  wire popcount30_eqge_core_094;
  wire popcount30_eqge_core_095;
  wire popcount30_eqge_core_097;
  wire popcount30_eqge_core_100;
  wire popcount30_eqge_core_101;
  wire popcount30_eqge_core_102;
  wire popcount30_eqge_core_103_not;
  wire popcount30_eqge_core_104;
  wire popcount30_eqge_core_105;
  wire popcount30_eqge_core_107;
  wire popcount30_eqge_core_108;
  wire popcount30_eqge_core_112;
  wire popcount30_eqge_core_114;
  wire popcount30_eqge_core_115;
  wire popcount30_eqge_core_116;
  wire popcount30_eqge_core_117;
  wire popcount30_eqge_core_118;
  wire popcount30_eqge_core_119;
  wire popcount30_eqge_core_120;
  wire popcount30_eqge_core_122;
  wire popcount30_eqge_core_123;
  wire popcount30_eqge_core_124;
  wire popcount30_eqge_core_126;
  wire popcount30_eqge_core_128;
  wire popcount30_eqge_core_130;
  wire popcount30_eqge_core_131;
  wire popcount30_eqge_core_134;
  wire popcount30_eqge_core_137;
  wire popcount30_eqge_core_140;
  wire popcount30_eqge_core_141;
  wire popcount30_eqge_core_142_not;
  wire popcount30_eqge_core_143;
  wire popcount30_eqge_core_144;
  wire popcount30_eqge_core_146;
  wire popcount30_eqge_core_147_not;
  wire popcount30_eqge_core_150;
  wire popcount30_eqge_core_153;
  wire popcount30_eqge_core_155;
  wire popcount30_eqge_core_156;
  wire popcount30_eqge_core_158;
  wire popcount30_eqge_core_159;
  wire popcount30_eqge_core_161;
  wire popcount30_eqge_core_162;
  wire popcount30_eqge_core_163;
  wire popcount30_eqge_core_164;
  wire popcount30_eqge_core_165;
  wire popcount30_eqge_core_167;
  wire popcount30_eqge_core_168;
  wire popcount30_eqge_core_169;
  wire popcount30_eqge_core_170;
  wire popcount30_eqge_core_171;
  wire popcount30_eqge_core_172;
  wire popcount30_eqge_core_173;
  wire popcount30_eqge_core_174;
  wire popcount30_eqge_core_175;
  wire popcount30_eqge_core_178;
  wire popcount30_eqge_core_180_not;
  wire popcount30_eqge_core_183;
  wire popcount30_eqge_core_185;
  wire popcount30_eqge_core_186;
  wire popcount30_eqge_core_187;
  wire popcount30_eqge_core_188;
  wire popcount30_eqge_core_190;
  wire popcount30_eqge_core_191;
  wire popcount30_eqge_core_194;
  wire popcount30_eqge_core_195;
  wire popcount30_eqge_core_197;
  wire popcount30_eqge_core_198;
  wire popcount30_eqge_core_203_not;
  wire popcount30_eqge_core_204;
  wire popcount30_eqge_core_205;
  wire popcount30_eqge_core_206;
  wire popcount30_eqge_core_208;
  wire popcount30_eqge_core_210;
  wire popcount30_eqge_core_212;
  wire popcount30_eqge_core_213;

  assign popcount30_eqge_core_032 = ~input_a[6];
  assign popcount30_eqge_core_034 = input_a[26] | input_a[9];
  assign popcount30_eqge_core_035 = ~input_a[26];
  assign popcount30_eqge_core_036 = input_a[23] ^ input_a[5];
  assign popcount30_eqge_core_037 = input_a[16] | input_a[20];
  assign popcount30_eqge_core_038 = ~(input_a[11] & input_a[14]);
  assign popcount30_eqge_core_040 = input_a[26] & input_a[9];
  assign popcount30_eqge_core_041 = ~(input_a[21] | input_a[0]);
  assign popcount30_eqge_core_042 = input_a[4] ^ input_a[7];
  assign popcount30_eqge_core_045 = input_a[3] ^ input_a[23];
  assign popcount30_eqge_core_046 = ~(input_a[12] | input_a[11]);
  assign popcount30_eqge_core_048 = input_a[17] & input_a[23];
  assign popcount30_eqge_core_049 = ~(input_a[9] ^ input_a[4]);
  assign popcount30_eqge_core_051 = input_a[6] ^ input_a[2];
  assign popcount30_eqge_core_052 = ~(input_a[25] | input_a[11]);
  assign popcount30_eqge_core_053 = input_a[14] | input_a[26];
  assign popcount30_eqge_core_054 = ~(input_a[27] ^ input_a[28]);
  assign popcount30_eqge_core_056 = ~(input_a[1] | input_a[9]);
  assign popcount30_eqge_core_057 = input_a[12] | input_a[28];
  assign popcount30_eqge_core_058 = ~(input_a[14] ^ input_a[7]);
  assign popcount30_eqge_core_059_not = ~input_a[23];
  assign popcount30_eqge_core_061 = ~input_a[6];
  assign popcount30_eqge_core_063 = input_a[19] & input_a[19];
  assign popcount30_eqge_core_064 = ~(input_a[22] & input_a[12]);
  assign popcount30_eqge_core_065 = input_a[5] ^ input_a[5];
  assign popcount30_eqge_core_070 = ~(input_a[17] | input_a[15]);
  assign popcount30_eqge_core_073 = input_a[11] & input_a[29];
  assign popcount30_eqge_core_074 = ~(input_a[18] ^ input_a[18]);
  assign popcount30_eqge_core_075 = ~input_a[18];
  assign popcount30_eqge_core_076 = input_a[5] | input_a[16];
  assign popcount30_eqge_core_077 = ~(input_a[2] ^ input_a[23]);
  assign popcount30_eqge_core_080 = ~(input_a[20] & input_a[14]);
  assign popcount30_eqge_core_084 = ~(input_a[9] | input_a[12]);
  assign popcount30_eqge_core_086 = ~(input_a[19] | input_a[24]);
  assign popcount30_eqge_core_088 = ~input_a[7];
  assign popcount30_eqge_core_090 = input_a[20] & input_a[19];
  assign popcount30_eqge_core_091 = input_a[1] | input_a[7];
  assign popcount30_eqge_core_092 = ~(input_a[20] & input_a[21]);
  assign popcount30_eqge_core_093 = input_a[16] ^ input_a[9];
  assign popcount30_eqge_core_094 = input_a[16] & input_a[14];
  assign popcount30_eqge_core_095 = ~(input_a[3] & input_a[16]);
  assign popcount30_eqge_core_097 = input_a[18] | input_a[4];
  assign popcount30_eqge_core_100 = input_a[28] & input_a[11];
  assign popcount30_eqge_core_101 = input_a[18] ^ input_a[16];
  assign popcount30_eqge_core_102 = ~(input_a[29] | input_a[4]);
  assign popcount30_eqge_core_103_not = ~input_a[2];
  assign popcount30_eqge_core_104 = ~(input_a[15] ^ input_a[24]);
  assign popcount30_eqge_core_105 = ~(input_a[11] ^ input_a[1]);
  assign popcount30_eqge_core_107 = ~(input_a[15] & input_a[28]);
  assign popcount30_eqge_core_108 = ~(input_a[24] | input_a[29]);
  assign popcount30_eqge_core_112 = ~input_a[11];
  assign popcount30_eqge_core_114 = input_a[12] ^ input_a[14];
  assign popcount30_eqge_core_115 = input_a[15] ^ input_a[29];
  assign popcount30_eqge_core_116 = input_a[15] & input_a[14];
  assign popcount30_eqge_core_117 = ~(input_a[18] & input_a[8]);
  assign popcount30_eqge_core_118 = input_a[19] ^ input_a[12];
  assign popcount30_eqge_core_119 = input_a[1] | input_a[21];
  assign popcount30_eqge_core_120 = input_a[2] ^ input_a[12];
  assign popcount30_eqge_core_122 = input_a[13] & input_a[8];
  assign popcount30_eqge_core_123 = input_a[8] | input_a[5];
  assign popcount30_eqge_core_124 = ~(input_a[6] ^ input_a[23]);
  assign popcount30_eqge_core_126 = ~(input_a[26] & input_a[6]);
  assign popcount30_eqge_core_128 = ~(input_a[28] & input_a[5]);
  assign popcount30_eqge_core_130 = ~(input_a[24] | input_a[5]);
  assign popcount30_eqge_core_131 = input_a[21] ^ input_a[23];
  assign popcount30_eqge_core_134 = ~(input_a[4] & input_a[11]);
  assign popcount30_eqge_core_137 = ~(input_a[13] ^ input_a[1]);
  assign popcount30_eqge_core_140 = ~(input_a[16] | input_a[26]);
  assign popcount30_eqge_core_141 = ~(input_a[11] ^ input_a[25]);
  assign popcount30_eqge_core_142_not = ~input_a[9];
  assign popcount30_eqge_core_143 = input_a[4] & input_a[16];
  assign popcount30_eqge_core_144 = ~(input_a[25] & input_a[4]);
  assign popcount30_eqge_core_146 = input_a[2] ^ input_a[1];
  assign popcount30_eqge_core_147_not = ~input_a[13];
  assign popcount30_eqge_core_150 = input_a[25] & input_a[2];
  assign popcount30_eqge_core_153 = input_a[26] & input_a[9];
  assign popcount30_eqge_core_155 = ~(input_a[28] ^ input_a[25]);
  assign popcount30_eqge_core_156 = input_a[1] ^ input_a[26];
  assign popcount30_eqge_core_158 = ~(input_a[19] | input_a[1]);
  assign popcount30_eqge_core_159 = input_a[22] | input_a[1];
  assign popcount30_eqge_core_161 = input_a[24] | input_a[26];
  assign popcount30_eqge_core_162 = ~input_a[24];
  assign popcount30_eqge_core_163 = ~(input_a[28] & input_a[21]);
  assign popcount30_eqge_core_164 = input_a[12] & input_a[13];
  assign popcount30_eqge_core_165 = input_a[29] & input_a[6];
  assign popcount30_eqge_core_167 = ~(input_a[19] & input_a[10]);
  assign popcount30_eqge_core_168 = ~(input_a[21] & input_a[22]);
  assign popcount30_eqge_core_169 = ~(input_a[3] | input_a[16]);
  assign popcount30_eqge_core_170 = input_a[24] | input_a[15];
  assign popcount30_eqge_core_171 = ~input_a[17];
  assign popcount30_eqge_core_172 = ~(input_a[19] | input_a[25]);
  assign popcount30_eqge_core_173 = ~input_a[17];
  assign popcount30_eqge_core_174 = input_a[27] & input_a[29];
  assign popcount30_eqge_core_175 = ~(input_a[26] | input_a[18]);
  assign popcount30_eqge_core_178 = ~(input_a[2] | input_a[19]);
  assign popcount30_eqge_core_180_not = ~input_a[7];
  assign popcount30_eqge_core_183 = ~input_a[13];
  assign popcount30_eqge_core_185 = ~input_a[21];
  assign popcount30_eqge_core_186 = ~(input_a[20] | input_a[29]);
  assign popcount30_eqge_core_187 = ~(input_a[17] & input_a[10]);
  assign popcount30_eqge_core_188 = input_a[23] | input_a[24];
  assign popcount30_eqge_core_190 = ~(input_a[29] & input_a[8]);
  assign popcount30_eqge_core_191 = input_a[7] | input_a[28];
  assign popcount30_eqge_core_194 = ~(input_a[0] | input_a[10]);
  assign popcount30_eqge_core_195 = ~(input_a[4] | input_a[21]);
  assign popcount30_eqge_core_197 = input_a[23] ^ input_a[6];
  assign popcount30_eqge_core_198 = ~input_a[14];
  assign popcount30_eqge_core_203_not = ~input_a[13];
  assign popcount30_eqge_core_204 = ~input_a[15];
  assign popcount30_eqge_core_205 = input_a[17] | input_a[11];
  assign popcount30_eqge_core_206 = input_a[13] ^ input_a[11];
  assign popcount30_eqge_core_208 = input_a[8] ^ input_a[18];
  assign popcount30_eqge_core_210 = ~(input_a[20] & input_a[19]);
  assign popcount30_eqge_core_212 = input_a[28] | input_a[13];
  assign popcount30_eqge_core_213 = ~(input_a[6] | input_a[24]);

  assign popcount30_eqge_out[0] = 1'b1;
  assign popcount30_eqge_out[1] = 1'b1;
  assign popcount30_eqge_out[2] = 1'b1;
  assign popcount30_eqge_out[3] = input_a[5];
  assign popcount30_eqge_out[4] = 1'b1;
endmodule