// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.37493
// WCE=18.0
// EP=0.937464%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_2p23(input [21:0] input_a, output [4:0] popcount22_2p23_out);
  wire popcount22_2p23_core_027;
  wire popcount22_2p23_core_028;
  wire popcount22_2p23_core_031;
  wire popcount22_2p23_core_032;
  wire popcount22_2p23_core_033;
  wire popcount22_2p23_core_035_not;
  wire popcount22_2p23_core_036;
  wire popcount22_2p23_core_037;
  wire popcount22_2p23_core_038;
  wire popcount22_2p23_core_039;
  wire popcount22_2p23_core_041;
  wire popcount22_2p23_core_042;
  wire popcount22_2p23_core_047;
  wire popcount22_2p23_core_048;
  wire popcount22_2p23_core_050_not;
  wire popcount22_2p23_core_052;
  wire popcount22_2p23_core_053;
  wire popcount22_2p23_core_054;
  wire popcount22_2p23_core_056_not;
  wire popcount22_2p23_core_058;
  wire popcount22_2p23_core_059;
  wire popcount22_2p23_core_061;
  wire popcount22_2p23_core_062;
  wire popcount22_2p23_core_063;
  wire popcount22_2p23_core_065;
  wire popcount22_2p23_core_068;
  wire popcount22_2p23_core_069;
  wire popcount22_2p23_core_070;
  wire popcount22_2p23_core_071;
  wire popcount22_2p23_core_072;
  wire popcount22_2p23_core_073;
  wire popcount22_2p23_core_074;
  wire popcount22_2p23_core_076;
  wire popcount22_2p23_core_081;
  wire popcount22_2p23_core_082;
  wire popcount22_2p23_core_084;
  wire popcount22_2p23_core_085;
  wire popcount22_2p23_core_087;
  wire popcount22_2p23_core_088;
  wire popcount22_2p23_core_090;
  wire popcount22_2p23_core_095;
  wire popcount22_2p23_core_096;
  wire popcount22_2p23_core_098;
  wire popcount22_2p23_core_099;
  wire popcount22_2p23_core_100;
  wire popcount22_2p23_core_101;
  wire popcount22_2p23_core_102;
  wire popcount22_2p23_core_104;
  wire popcount22_2p23_core_105;
  wire popcount22_2p23_core_107;
  wire popcount22_2p23_core_108_not;
  wire popcount22_2p23_core_111;
  wire popcount22_2p23_core_112;
  wire popcount22_2p23_core_113;
  wire popcount22_2p23_core_115;
  wire popcount22_2p23_core_116;
  wire popcount22_2p23_core_117;
  wire popcount22_2p23_core_118;
  wire popcount22_2p23_core_119;
  wire popcount22_2p23_core_121_not;
  wire popcount22_2p23_core_124;
  wire popcount22_2p23_core_125;
  wire popcount22_2p23_core_127_not;
  wire popcount22_2p23_core_129;
  wire popcount22_2p23_core_130;
  wire popcount22_2p23_core_131;
  wire popcount22_2p23_core_132;
  wire popcount22_2p23_core_136;
  wire popcount22_2p23_core_137;
  wire popcount22_2p23_core_138;
  wire popcount22_2p23_core_139;
  wire popcount22_2p23_core_140;
  wire popcount22_2p23_core_141;
  wire popcount22_2p23_core_142;
  wire popcount22_2p23_core_143;
  wire popcount22_2p23_core_145;
  wire popcount22_2p23_core_146;
  wire popcount22_2p23_core_148;
  wire popcount22_2p23_core_149;
  wire popcount22_2p23_core_152;
  wire popcount22_2p23_core_153;
  wire popcount22_2p23_core_155;
  wire popcount22_2p23_core_156;
  wire popcount22_2p23_core_159;
  wire popcount22_2p23_core_160;
  wire popcount22_2p23_core_161;

  assign popcount22_2p23_core_027 = ~(input_a[14] ^ input_a[13]);
  assign popcount22_2p23_core_028 = input_a[18] & input_a[15];
  assign popcount22_2p23_core_031 = input_a[17] ^ input_a[19];
  assign popcount22_2p23_core_032 = ~(input_a[19] ^ input_a[1]);
  assign popcount22_2p23_core_033 = ~(input_a[19] | input_a[9]);
  assign popcount22_2p23_core_035_not = ~input_a[17];
  assign popcount22_2p23_core_036 = input_a[9] ^ input_a[4];
  assign popcount22_2p23_core_037 = input_a[1] & input_a[21];
  assign popcount22_2p23_core_038 = ~(input_a[9] & input_a[2]);
  assign popcount22_2p23_core_039 = ~(input_a[12] ^ input_a[14]);
  assign popcount22_2p23_core_041 = ~(input_a[13] & input_a[4]);
  assign popcount22_2p23_core_042 = input_a[6] | input_a[12];
  assign popcount22_2p23_core_047 = ~(input_a[12] | input_a[14]);
  assign popcount22_2p23_core_048 = input_a[13] | input_a[15];
  assign popcount22_2p23_core_050_not = ~input_a[1];
  assign popcount22_2p23_core_052 = input_a[1] & input_a[13];
  assign popcount22_2p23_core_053 = ~input_a[17];
  assign popcount22_2p23_core_054 = ~(input_a[6] | input_a[0]);
  assign popcount22_2p23_core_056_not = ~input_a[2];
  assign popcount22_2p23_core_058 = ~(input_a[21] ^ input_a[18]);
  assign popcount22_2p23_core_059 = ~(input_a[13] & input_a[2]);
  assign popcount22_2p23_core_061 = ~(input_a[0] & input_a[19]);
  assign popcount22_2p23_core_062 = ~(input_a[4] & input_a[15]);
  assign popcount22_2p23_core_063 = ~(input_a[11] ^ input_a[12]);
  assign popcount22_2p23_core_065 = ~(input_a[5] | input_a[18]);
  assign popcount22_2p23_core_068 = input_a[3] ^ input_a[2];
  assign popcount22_2p23_core_069 = ~(input_a[9] ^ input_a[0]);
  assign popcount22_2p23_core_070 = input_a[17] ^ input_a[4];
  assign popcount22_2p23_core_071 = input_a[20] & input_a[8];
  assign popcount22_2p23_core_072 = ~input_a[14];
  assign popcount22_2p23_core_073 = input_a[17] & input_a[18];
  assign popcount22_2p23_core_074 = ~(input_a[3] ^ input_a[3]);
  assign popcount22_2p23_core_076 = input_a[20] | input_a[2];
  assign popcount22_2p23_core_081 = ~(input_a[7] ^ input_a[1]);
  assign popcount22_2p23_core_082 = input_a[19] & input_a[12];
  assign popcount22_2p23_core_084 = ~input_a[20];
  assign popcount22_2p23_core_085 = ~input_a[14];
  assign popcount22_2p23_core_087 = input_a[0] | input_a[5];
  assign popcount22_2p23_core_088 = input_a[11] & input_a[13];
  assign popcount22_2p23_core_090 = ~input_a[12];
  assign popcount22_2p23_core_095 = ~(input_a[2] | input_a[20]);
  assign popcount22_2p23_core_096 = ~(input_a[20] ^ input_a[6]);
  assign popcount22_2p23_core_098 = ~(input_a[9] ^ input_a[19]);
  assign popcount22_2p23_core_099 = input_a[18] ^ input_a[5];
  assign popcount22_2p23_core_100 = input_a[7] & input_a[9];
  assign popcount22_2p23_core_101 = input_a[10] ^ input_a[11];
  assign popcount22_2p23_core_102 = input_a[20] | input_a[17];
  assign popcount22_2p23_core_104 = ~(input_a[15] & input_a[19]);
  assign popcount22_2p23_core_105 = input_a[13] | input_a[2];
  assign popcount22_2p23_core_107 = ~(input_a[5] ^ input_a[15]);
  assign popcount22_2p23_core_108_not = ~input_a[17];
  assign popcount22_2p23_core_111 = ~(input_a[2] ^ input_a[18]);
  assign popcount22_2p23_core_112 = input_a[8] | input_a[20];
  assign popcount22_2p23_core_113 = input_a[3] ^ input_a[5];
  assign popcount22_2p23_core_115 = ~(input_a[9] | input_a[6]);
  assign popcount22_2p23_core_116 = ~(input_a[11] ^ input_a[1]);
  assign popcount22_2p23_core_117 = ~input_a[1];
  assign popcount22_2p23_core_118 = ~(input_a[8] ^ input_a[11]);
  assign popcount22_2p23_core_119 = input_a[16] & input_a[12];
  assign popcount22_2p23_core_121_not = ~input_a[10];
  assign popcount22_2p23_core_124 = ~input_a[14];
  assign popcount22_2p23_core_125 = input_a[16] ^ input_a[12];
  assign popcount22_2p23_core_127_not = ~input_a[17];
  assign popcount22_2p23_core_129 = input_a[4] ^ input_a[10];
  assign popcount22_2p23_core_130 = input_a[16] ^ input_a[15];
  assign popcount22_2p23_core_131 = ~input_a[10];
  assign popcount22_2p23_core_132 = input_a[6] ^ input_a[5];
  assign popcount22_2p23_core_136 = ~(input_a[13] ^ input_a[4]);
  assign popcount22_2p23_core_137 = ~(input_a[12] ^ input_a[9]);
  assign popcount22_2p23_core_138 = ~(input_a[1] ^ input_a[13]);
  assign popcount22_2p23_core_139 = ~(input_a[9] ^ input_a[4]);
  assign popcount22_2p23_core_140 = input_a[7] ^ input_a[19];
  assign popcount22_2p23_core_141 = ~(input_a[2] | input_a[11]);
  assign popcount22_2p23_core_142 = ~input_a[20];
  assign popcount22_2p23_core_143 = ~(input_a[2] | input_a[8]);
  assign popcount22_2p23_core_145 = input_a[21] & input_a[19];
  assign popcount22_2p23_core_146 = ~(input_a[15] & input_a[8]);
  assign popcount22_2p23_core_148 = ~input_a[3];
  assign popcount22_2p23_core_149 = ~(input_a[17] & input_a[0]);
  assign popcount22_2p23_core_152 = ~(input_a[0] | input_a[7]);
  assign popcount22_2p23_core_153 = input_a[15] & input_a[0];
  assign popcount22_2p23_core_155 = ~(input_a[13] & input_a[4]);
  assign popcount22_2p23_core_156 = input_a[18] | input_a[10];
  assign popcount22_2p23_core_159 = ~input_a[11];
  assign popcount22_2p23_core_160 = ~(input_a[4] | input_a[11]);
  assign popcount22_2p23_core_161 = ~(input_a[2] & input_a[15]);

  assign popcount22_2p23_out[0] = 1'b1;
  assign popcount22_2p23_out[1] = 1'b1;
  assign popcount22_2p23_out[2] = input_a[18];
  assign popcount22_2p23_out[3] = 1'b0;
  assign popcount22_2p23_out[4] = 1'b0;
endmodule