// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.16697
// WCE=15.0
// EP=0.855536%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_ihkh(input [29:0] input_a, output [4:0] popcount30_ihkh_out);
  wire popcount30_ihkh_core_032;
  wire popcount30_ihkh_core_033;
  wire popcount30_ihkh_core_034;
  wire popcount30_ihkh_core_036;
  wire popcount30_ihkh_core_037;
  wire popcount30_ihkh_core_038;
  wire popcount30_ihkh_core_040_not;
  wire popcount30_ihkh_core_042;
  wire popcount30_ihkh_core_043;
  wire popcount30_ihkh_core_044;
  wire popcount30_ihkh_core_046;
  wire popcount30_ihkh_core_047;
  wire popcount30_ihkh_core_050;
  wire popcount30_ihkh_core_051;
  wire popcount30_ihkh_core_052;
  wire popcount30_ihkh_core_053;
  wire popcount30_ihkh_core_054;
  wire popcount30_ihkh_core_055;
  wire popcount30_ihkh_core_056;
  wire popcount30_ihkh_core_057;
  wire popcount30_ihkh_core_058_not;
  wire popcount30_ihkh_core_060;
  wire popcount30_ihkh_core_061;
  wire popcount30_ihkh_core_065;
  wire popcount30_ihkh_core_069;
  wire popcount30_ihkh_core_070;
  wire popcount30_ihkh_core_071;
  wire popcount30_ihkh_core_074;
  wire popcount30_ihkh_core_075;
  wire popcount30_ihkh_core_077;
  wire popcount30_ihkh_core_078;
  wire popcount30_ihkh_core_079;
  wire popcount30_ihkh_core_080;
  wire popcount30_ihkh_core_082;
  wire popcount30_ihkh_core_083;
  wire popcount30_ihkh_core_085;
  wire popcount30_ihkh_core_086;
  wire popcount30_ihkh_core_087;
  wire popcount30_ihkh_core_089;
  wire popcount30_ihkh_core_090;
  wire popcount30_ihkh_core_092;
  wire popcount30_ihkh_core_094;
  wire popcount30_ihkh_core_095;
  wire popcount30_ihkh_core_096;
  wire popcount30_ihkh_core_097_not;
  wire popcount30_ihkh_core_098;
  wire popcount30_ihkh_core_099;
  wire popcount30_ihkh_core_100;
  wire popcount30_ihkh_core_101;
  wire popcount30_ihkh_core_102;
  wire popcount30_ihkh_core_103;
  wire popcount30_ihkh_core_104;
  wire popcount30_ihkh_core_106;
  wire popcount30_ihkh_core_107;
  wire popcount30_ihkh_core_108;
  wire popcount30_ihkh_core_109;
  wire popcount30_ihkh_core_110;
  wire popcount30_ihkh_core_111;
  wire popcount30_ihkh_core_112;
  wire popcount30_ihkh_core_113;
  wire popcount30_ihkh_core_114;
  wire popcount30_ihkh_core_115;
  wire popcount30_ihkh_core_116;
  wire popcount30_ihkh_core_117;
  wire popcount30_ihkh_core_118;
  wire popcount30_ihkh_core_119;
  wire popcount30_ihkh_core_122;
  wire popcount30_ihkh_core_123;
  wire popcount30_ihkh_core_128;
  wire popcount30_ihkh_core_130;
  wire popcount30_ihkh_core_132;
  wire popcount30_ihkh_core_133;
  wire popcount30_ihkh_core_134;
  wire popcount30_ihkh_core_135;
  wire popcount30_ihkh_core_136;
  wire popcount30_ihkh_core_137;
  wire popcount30_ihkh_core_138;
  wire popcount30_ihkh_core_139;
  wire popcount30_ihkh_core_140;
  wire popcount30_ihkh_core_143;
  wire popcount30_ihkh_core_144;
  wire popcount30_ihkh_core_145;
  wire popcount30_ihkh_core_148;
  wire popcount30_ihkh_core_149;
  wire popcount30_ihkh_core_151;
  wire popcount30_ihkh_core_152;
  wire popcount30_ihkh_core_156;
  wire popcount30_ihkh_core_158;
  wire popcount30_ihkh_core_159;
  wire popcount30_ihkh_core_160;
  wire popcount30_ihkh_core_162;
  wire popcount30_ihkh_core_163;
  wire popcount30_ihkh_core_164;
  wire popcount30_ihkh_core_165;
  wire popcount30_ihkh_core_167;
  wire popcount30_ihkh_core_168;
  wire popcount30_ihkh_core_171;
  wire popcount30_ihkh_core_173;
  wire popcount30_ihkh_core_174_not;
  wire popcount30_ihkh_core_176;
  wire popcount30_ihkh_core_177;
  wire popcount30_ihkh_core_178;
  wire popcount30_ihkh_core_180;
  wire popcount30_ihkh_core_181;
  wire popcount30_ihkh_core_183;
  wire popcount30_ihkh_core_184;
  wire popcount30_ihkh_core_186;
  wire popcount30_ihkh_core_187;
  wire popcount30_ihkh_core_188;
  wire popcount30_ihkh_core_190;
  wire popcount30_ihkh_core_196;
  wire popcount30_ihkh_core_197;
  wire popcount30_ihkh_core_198;
  wire popcount30_ihkh_core_201;
  wire popcount30_ihkh_core_202;
  wire popcount30_ihkh_core_204;
  wire popcount30_ihkh_core_206;
  wire popcount30_ihkh_core_209;
  wire popcount30_ihkh_core_210;
  wire popcount30_ihkh_core_211;
  wire popcount30_ihkh_core_212;
  wire popcount30_ihkh_core_213;

  assign popcount30_ihkh_core_032 = ~(input_a[23] ^ input_a[15]);
  assign popcount30_ihkh_core_033 = ~(input_a[5] ^ input_a[27]);
  assign popcount30_ihkh_core_034 = input_a[9] | input_a[12];
  assign popcount30_ihkh_core_036 = ~(input_a[3] & input_a[21]);
  assign popcount30_ihkh_core_037 = input_a[23] | input_a[17];
  assign popcount30_ihkh_core_038 = ~(input_a[8] & input_a[14]);
  assign popcount30_ihkh_core_040_not = ~input_a[15];
  assign popcount30_ihkh_core_042 = ~(input_a[3] & input_a[2]);
  assign popcount30_ihkh_core_043 = ~(input_a[27] ^ input_a[21]);
  assign popcount30_ihkh_core_044 = input_a[4] | input_a[20];
  assign popcount30_ihkh_core_046 = ~(input_a[26] | input_a[8]);
  assign popcount30_ihkh_core_047 = input_a[28] | input_a[0];
  assign popcount30_ihkh_core_050 = ~(input_a[27] ^ input_a[21]);
  assign popcount30_ihkh_core_051 = input_a[9] & input_a[23];
  assign popcount30_ihkh_core_052 = input_a[0] & input_a[25];
  assign popcount30_ihkh_core_053 = ~(input_a[4] | input_a[27]);
  assign popcount30_ihkh_core_054 = input_a[17] & input_a[14];
  assign popcount30_ihkh_core_055 = input_a[21] & input_a[24];
  assign popcount30_ihkh_core_056 = input_a[29] ^ input_a[22];
  assign popcount30_ihkh_core_057 = ~(input_a[15] ^ input_a[24]);
  assign popcount30_ihkh_core_058_not = ~input_a[17];
  assign popcount30_ihkh_core_060 = ~input_a[15];
  assign popcount30_ihkh_core_061 = ~(input_a[26] & input_a[2]);
  assign popcount30_ihkh_core_065 = input_a[25] ^ input_a[10];
  assign popcount30_ihkh_core_069 = ~(input_a[4] & input_a[21]);
  assign popcount30_ihkh_core_070 = input_a[25] ^ input_a[20];
  assign popcount30_ihkh_core_071 = input_a[17] & input_a[8];
  assign popcount30_ihkh_core_074 = ~(input_a[8] ^ input_a[10]);
  assign popcount30_ihkh_core_075 = input_a[28] ^ input_a[16];
  assign popcount30_ihkh_core_077 = ~(input_a[29] | input_a[16]);
  assign popcount30_ihkh_core_078 = input_a[18] & input_a[3];
  assign popcount30_ihkh_core_079 = ~(input_a[6] | input_a[5]);
  assign popcount30_ihkh_core_080 = input_a[17] ^ input_a[1];
  assign popcount30_ihkh_core_082 = input_a[3] & input_a[6];
  assign popcount30_ihkh_core_083 = ~(input_a[23] | input_a[16]);
  assign popcount30_ihkh_core_085 = ~(input_a[27] ^ input_a[10]);
  assign popcount30_ihkh_core_086 = ~(input_a[4] ^ input_a[11]);
  assign popcount30_ihkh_core_087 = ~(input_a[28] ^ input_a[1]);
  assign popcount30_ihkh_core_089 = ~input_a[19];
  assign popcount30_ihkh_core_090 = ~(input_a[18] ^ input_a[26]);
  assign popcount30_ihkh_core_092 = ~input_a[16];
  assign popcount30_ihkh_core_094 = ~(input_a[6] & input_a[16]);
  assign popcount30_ihkh_core_095 = ~(input_a[24] | input_a[28]);
  assign popcount30_ihkh_core_096 = ~(input_a[6] & input_a[0]);
  assign popcount30_ihkh_core_097_not = ~input_a[0];
  assign popcount30_ihkh_core_098 = ~(input_a[24] & input_a[20]);
  assign popcount30_ihkh_core_099 = input_a[26] ^ input_a[24];
  assign popcount30_ihkh_core_100 = ~(input_a[0] | input_a[8]);
  assign popcount30_ihkh_core_101 = ~(input_a[1] | input_a[13]);
  assign popcount30_ihkh_core_102 = ~input_a[7];
  assign popcount30_ihkh_core_103 = input_a[4] ^ input_a[12];
  assign popcount30_ihkh_core_104 = ~input_a[0];
  assign popcount30_ihkh_core_106 = ~(input_a[4] ^ input_a[25]);
  assign popcount30_ihkh_core_107 = ~(input_a[24] & input_a[1]);
  assign popcount30_ihkh_core_108 = ~(input_a[1] & input_a[15]);
  assign popcount30_ihkh_core_109 = ~(input_a[25] & input_a[12]);
  assign popcount30_ihkh_core_110 = input_a[0] ^ input_a[9];
  assign popcount30_ihkh_core_111 = input_a[10] & input_a[25];
  assign popcount30_ihkh_core_112 = input_a[29] ^ input_a[0];
  assign popcount30_ihkh_core_113 = ~(input_a[15] & input_a[6]);
  assign popcount30_ihkh_core_114 = input_a[14] | input_a[20];
  assign popcount30_ihkh_core_115 = input_a[21] & input_a[11];
  assign popcount30_ihkh_core_116 = ~(input_a[4] & input_a[3]);
  assign popcount30_ihkh_core_117 = ~(input_a[6] ^ input_a[5]);
  assign popcount30_ihkh_core_118 = ~(input_a[28] ^ input_a[13]);
  assign popcount30_ihkh_core_119 = ~input_a[8];
  assign popcount30_ihkh_core_122 = input_a[26] | input_a[28];
  assign popcount30_ihkh_core_123 = ~(input_a[12] | input_a[7]);
  assign popcount30_ihkh_core_128 = input_a[22] | input_a[24];
  assign popcount30_ihkh_core_130 = input_a[16] ^ input_a[8];
  assign popcount30_ihkh_core_132 = input_a[5] & input_a[26];
  assign popcount30_ihkh_core_133 = input_a[18] & input_a[10];
  assign popcount30_ihkh_core_134 = input_a[16] ^ input_a[24];
  assign popcount30_ihkh_core_135 = ~input_a[2];
  assign popcount30_ihkh_core_136 = input_a[24] & input_a[16];
  assign popcount30_ihkh_core_137 = ~(input_a[17] & input_a[1]);
  assign popcount30_ihkh_core_138 = input_a[29] ^ input_a[0];
  assign popcount30_ihkh_core_139 = ~(input_a[28] | input_a[4]);
  assign popcount30_ihkh_core_140 = input_a[8] & input_a[28];
  assign popcount30_ihkh_core_143 = ~(input_a[3] ^ input_a[27]);
  assign popcount30_ihkh_core_144 = ~input_a[29];
  assign popcount30_ihkh_core_145 = ~input_a[5];
  assign popcount30_ihkh_core_148 = ~input_a[15];
  assign popcount30_ihkh_core_149 = ~input_a[24];
  assign popcount30_ihkh_core_151 = ~input_a[16];
  assign popcount30_ihkh_core_152 = input_a[9] & input_a[18];
  assign popcount30_ihkh_core_156 = ~(input_a[10] | input_a[2]);
  assign popcount30_ihkh_core_158 = input_a[17] & input_a[22];
  assign popcount30_ihkh_core_159 = ~(input_a[8] | input_a[14]);
  assign popcount30_ihkh_core_160 = input_a[12] ^ input_a[13];
  assign popcount30_ihkh_core_162 = input_a[0] | input_a[13];
  assign popcount30_ihkh_core_163 = input_a[7] ^ input_a[0];
  assign popcount30_ihkh_core_164 = ~(input_a[5] | input_a[21]);
  assign popcount30_ihkh_core_165 = ~input_a[3];
  assign popcount30_ihkh_core_167 = ~(input_a[26] & input_a[11]);
  assign popcount30_ihkh_core_168 = ~input_a[28];
  assign popcount30_ihkh_core_171 = ~input_a[1];
  assign popcount30_ihkh_core_173 = ~input_a[15];
  assign popcount30_ihkh_core_174_not = ~input_a[17];
  assign popcount30_ihkh_core_176 = ~input_a[22];
  assign popcount30_ihkh_core_177 = input_a[13] ^ input_a[16];
  assign popcount30_ihkh_core_178 = ~(input_a[1] & input_a[9]);
  assign popcount30_ihkh_core_180 = ~input_a[19];
  assign popcount30_ihkh_core_181 = input_a[9] | input_a[2];
  assign popcount30_ihkh_core_183 = input_a[5] ^ input_a[5];
  assign popcount30_ihkh_core_184 = ~(input_a[6] | input_a[25]);
  assign popcount30_ihkh_core_186 = input_a[22] ^ input_a[22];
  assign popcount30_ihkh_core_187 = ~(input_a[14] & input_a[8]);
  assign popcount30_ihkh_core_188 = ~(input_a[24] | input_a[2]);
  assign popcount30_ihkh_core_190 = ~input_a[8];
  assign popcount30_ihkh_core_196 = ~(input_a[7] & input_a[27]);
  assign popcount30_ihkh_core_197 = input_a[28] & input_a[0];
  assign popcount30_ihkh_core_198 = input_a[0] ^ input_a[0];
  assign popcount30_ihkh_core_201 = ~(input_a[20] & input_a[12]);
  assign popcount30_ihkh_core_202 = ~(input_a[18] & input_a[14]);
  assign popcount30_ihkh_core_204 = input_a[13] ^ input_a[14];
  assign popcount30_ihkh_core_206 = ~(input_a[7] | input_a[16]);
  assign popcount30_ihkh_core_209 = input_a[24] & input_a[0];
  assign popcount30_ihkh_core_210 = input_a[26] & input_a[28];
  assign popcount30_ihkh_core_211 = ~(input_a[13] ^ input_a[13]);
  assign popcount30_ihkh_core_212 = input_a[26] & input_a[2];
  assign popcount30_ihkh_core_213 = input_a[1] ^ input_a[6];

  assign popcount30_ihkh_out[0] = input_a[23];
  assign popcount30_ihkh_out[1] = 1'b1;
  assign popcount30_ihkh_out[2] = 1'b1;
  assign popcount30_ihkh_out[3] = 1'b1;
  assign popcount30_ihkh_out[4] = 1'b0;
endmodule