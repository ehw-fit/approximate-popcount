// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.86165
// WCE=10.0
// EP=0.834037%
// Printed PDK parameters:
//  Area=94639173.0
//  Delay=91963824.0
//  Power=4061200.0

module popcount47_ubuz(input [46:0] input_a, output [5:0] popcount47_ubuz_out);
  wire popcount47_ubuz_core_049;
  wire popcount47_ubuz_core_050;
  wire popcount47_ubuz_core_051;
  wire popcount47_ubuz_core_052;
  wire popcount47_ubuz_core_054;
  wire popcount47_ubuz_core_057;
  wire popcount47_ubuz_core_058;
  wire popcount47_ubuz_core_059;
  wire popcount47_ubuz_core_061;
  wire popcount47_ubuz_core_062;
  wire popcount47_ubuz_core_063;
  wire popcount47_ubuz_core_066;
  wire popcount47_ubuz_core_067;
  wire popcount47_ubuz_core_068;
  wire popcount47_ubuz_core_069;
  wire popcount47_ubuz_core_070;
  wire popcount47_ubuz_core_072;
  wire popcount47_ubuz_core_073;
  wire popcount47_ubuz_core_074;
  wire popcount47_ubuz_core_075;
  wire popcount47_ubuz_core_076;
  wire popcount47_ubuz_core_078;
  wire popcount47_ubuz_core_079;
  wire popcount47_ubuz_core_080;
  wire popcount47_ubuz_core_081;
  wire popcount47_ubuz_core_083;
  wire popcount47_ubuz_core_084;
  wire popcount47_ubuz_core_088;
  wire popcount47_ubuz_core_089;
  wire popcount47_ubuz_core_099_not;
  wire popcount47_ubuz_core_103;
  wire popcount47_ubuz_core_106;
  wire popcount47_ubuz_core_107;
  wire popcount47_ubuz_core_108;
  wire popcount47_ubuz_core_110;
  wire popcount47_ubuz_core_111;
  wire popcount47_ubuz_core_113;
  wire popcount47_ubuz_core_114;
  wire popcount47_ubuz_core_115;
  wire popcount47_ubuz_core_116;
  wire popcount47_ubuz_core_117;
  wire popcount47_ubuz_core_118;
  wire popcount47_ubuz_core_119;
  wire popcount47_ubuz_core_120;
  wire popcount47_ubuz_core_121;
  wire popcount47_ubuz_core_122;
  wire popcount47_ubuz_core_123;
  wire popcount47_ubuz_core_124;
  wire popcount47_ubuz_core_125;
  wire popcount47_ubuz_core_127;
  wire popcount47_ubuz_core_129;
  wire popcount47_ubuz_core_131;
  wire popcount47_ubuz_core_132;
  wire popcount47_ubuz_core_133;
  wire popcount47_ubuz_core_134;
  wire popcount47_ubuz_core_135;
  wire popcount47_ubuz_core_136;
  wire popcount47_ubuz_core_137;
  wire popcount47_ubuz_core_138;
  wire popcount47_ubuz_core_139;
  wire popcount47_ubuz_core_140;
  wire popcount47_ubuz_core_141;
  wire popcount47_ubuz_core_142;
  wire popcount47_ubuz_core_143;
  wire popcount47_ubuz_core_144;
  wire popcount47_ubuz_core_145;
  wire popcount47_ubuz_core_146;
  wire popcount47_ubuz_core_147;
  wire popcount47_ubuz_core_148;
  wire popcount47_ubuz_core_149;
  wire popcount47_ubuz_core_151;
  wire popcount47_ubuz_core_153;
  wire popcount47_ubuz_core_154;
  wire popcount47_ubuz_core_155;
  wire popcount47_ubuz_core_156;
  wire popcount47_ubuz_core_157;
  wire popcount47_ubuz_core_158;
  wire popcount47_ubuz_core_159;
  wire popcount47_ubuz_core_160;
  wire popcount47_ubuz_core_161;
  wire popcount47_ubuz_core_162;
  wire popcount47_ubuz_core_163;
  wire popcount47_ubuz_core_164;
  wire popcount47_ubuz_core_165;
  wire popcount47_ubuz_core_166;
  wire popcount47_ubuz_core_170;
  wire popcount47_ubuz_core_171;
  wire popcount47_ubuz_core_172;
  wire popcount47_ubuz_core_173;
  wire popcount47_ubuz_core_176;
  wire popcount47_ubuz_core_177;
  wire popcount47_ubuz_core_179;
  wire popcount47_ubuz_core_180;
  wire popcount47_ubuz_core_181;
  wire popcount47_ubuz_core_182;
  wire popcount47_ubuz_core_183;
  wire popcount47_ubuz_core_184;
  wire popcount47_ubuz_core_185;
  wire popcount47_ubuz_core_186;
  wire popcount47_ubuz_core_187;
  wire popcount47_ubuz_core_188;
  wire popcount47_ubuz_core_190;
  wire popcount47_ubuz_core_193;
  wire popcount47_ubuz_core_194;
  wire popcount47_ubuz_core_195;
  wire popcount47_ubuz_core_199;
  wire popcount47_ubuz_core_200;
  wire popcount47_ubuz_core_201;
  wire popcount47_ubuz_core_202;
  wire popcount47_ubuz_core_203;
  wire popcount47_ubuz_core_204;
  wire popcount47_ubuz_core_205;
  wire popcount47_ubuz_core_207;
  wire popcount47_ubuz_core_210;
  wire popcount47_ubuz_core_211;
  wire popcount47_ubuz_core_216;
  wire popcount47_ubuz_core_218;
  wire popcount47_ubuz_core_219;
  wire popcount47_ubuz_core_220;
  wire popcount47_ubuz_core_221;
  wire popcount47_ubuz_core_222;
  wire popcount47_ubuz_core_223;
  wire popcount47_ubuz_core_224;
  wire popcount47_ubuz_core_225;
  wire popcount47_ubuz_core_226;
  wire popcount47_ubuz_core_227;
  wire popcount47_ubuz_core_230;
  wire popcount47_ubuz_core_232;
  wire popcount47_ubuz_core_233;
  wire popcount47_ubuz_core_234;
  wire popcount47_ubuz_core_235;
  wire popcount47_ubuz_core_236;
  wire popcount47_ubuz_core_238;
  wire popcount47_ubuz_core_240;
  wire popcount47_ubuz_core_241;
  wire popcount47_ubuz_core_243;
  wire popcount47_ubuz_core_244;
  wire popcount47_ubuz_core_245;
  wire popcount47_ubuz_core_246;
  wire popcount47_ubuz_core_247;
  wire popcount47_ubuz_core_248;
  wire popcount47_ubuz_core_249;
  wire popcount47_ubuz_core_250;
  wire popcount47_ubuz_core_251;
  wire popcount47_ubuz_core_252;
  wire popcount47_ubuz_core_253;
  wire popcount47_ubuz_core_255;
  wire popcount47_ubuz_core_260;
  wire popcount47_ubuz_core_269;
  wire popcount47_ubuz_core_270;
  wire popcount47_ubuz_core_272;
  wire popcount47_ubuz_core_273;
  wire popcount47_ubuz_core_274;
  wire popcount47_ubuz_core_275;
  wire popcount47_ubuz_core_276;
  wire popcount47_ubuz_core_277;
  wire popcount47_ubuz_core_280;
  wire popcount47_ubuz_core_281;
  wire popcount47_ubuz_core_283;
  wire popcount47_ubuz_core_284;
  wire popcount47_ubuz_core_285;
  wire popcount47_ubuz_core_286;
  wire popcount47_ubuz_core_287;
  wire popcount47_ubuz_core_288;
  wire popcount47_ubuz_core_289;
  wire popcount47_ubuz_core_291;
  wire popcount47_ubuz_core_292;
  wire popcount47_ubuz_core_293;
  wire popcount47_ubuz_core_295;
  wire popcount47_ubuz_core_296;
  wire popcount47_ubuz_core_298;
  wire popcount47_ubuz_core_301;
  wire popcount47_ubuz_core_304;
  wire popcount47_ubuz_core_307;
  wire popcount47_ubuz_core_309;
  wire popcount47_ubuz_core_310;
  wire popcount47_ubuz_core_316;
  wire popcount47_ubuz_core_317;
  wire popcount47_ubuz_core_321;
  wire popcount47_ubuz_core_322;
  wire popcount47_ubuz_core_323;
  wire popcount47_ubuz_core_325;
  wire popcount47_ubuz_core_326;
  wire popcount47_ubuz_core_327;
  wire popcount47_ubuz_core_328;
  wire popcount47_ubuz_core_329;
  wire popcount47_ubuz_core_330;
  wire popcount47_ubuz_core_331;
  wire popcount47_ubuz_core_332;
  wire popcount47_ubuz_core_333;
  wire popcount47_ubuz_core_334;
  wire popcount47_ubuz_core_335;
  wire popcount47_ubuz_core_336;
  wire popcount47_ubuz_core_337;
  wire popcount47_ubuz_core_338;
  wire popcount47_ubuz_core_339;
  wire popcount47_ubuz_core_340;
  wire popcount47_ubuz_core_344;
  wire popcount47_ubuz_core_345;
  wire popcount47_ubuz_core_347;
  wire popcount47_ubuz_core_348;
  wire popcount47_ubuz_core_349;
  wire popcount47_ubuz_core_350;
  wire popcount47_ubuz_core_351;
  wire popcount47_ubuz_core_352;
  wire popcount47_ubuz_core_353;
  wire popcount47_ubuz_core_354;
  wire popcount47_ubuz_core_355;
  wire popcount47_ubuz_core_356;
  wire popcount47_ubuz_core_357;
  wire popcount47_ubuz_core_358;
  wire popcount47_ubuz_core_359;
  wire popcount47_ubuz_core_360;
  wire popcount47_ubuz_core_361;
  wire popcount47_ubuz_core_362;
  wire popcount47_ubuz_core_363;
  wire popcount47_ubuz_core_364;
  wire popcount47_ubuz_core_365;
  wire popcount47_ubuz_core_366;
  wire popcount47_ubuz_core_367;
  wire popcount47_ubuz_core_369;
  wire popcount47_ubuz_core_372;

  assign popcount47_ubuz_core_049 = ~(input_a[19] | input_a[45]);
  assign popcount47_ubuz_core_050 = ~(input_a[1] ^ input_a[24]);
  assign popcount47_ubuz_core_051 = input_a[41] & input_a[43];
  assign popcount47_ubuz_core_052 = ~(input_a[19] & input_a[30]);
  assign popcount47_ubuz_core_054 = input_a[32] & input_a[3];
  assign popcount47_ubuz_core_057 = ~(input_a[27] | input_a[15]);
  assign popcount47_ubuz_core_058 = ~input_a[20];
  assign popcount47_ubuz_core_059 = input_a[38] & input_a[25];
  assign popcount47_ubuz_core_061 = ~(input_a[39] & input_a[11]);
  assign popcount47_ubuz_core_062 = ~(input_a[27] ^ input_a[43]);
  assign popcount47_ubuz_core_063 = ~input_a[42];
  assign popcount47_ubuz_core_066 = input_a[6] ^ input_a[7];
  assign popcount47_ubuz_core_067 = input_a[6] & input_a[7];
  assign popcount47_ubuz_core_068 = input_a[5] ^ popcount47_ubuz_core_066;
  assign popcount47_ubuz_core_069 = input_a[5] & popcount47_ubuz_core_066;
  assign popcount47_ubuz_core_070 = popcount47_ubuz_core_067 | popcount47_ubuz_core_069;
  assign popcount47_ubuz_core_072 = input_a[9] ^ input_a[10];
  assign popcount47_ubuz_core_073 = input_a[9] & input_a[10];
  assign popcount47_ubuz_core_074 = input_a[8] ^ popcount47_ubuz_core_072;
  assign popcount47_ubuz_core_075 = input_a[8] & popcount47_ubuz_core_072;
  assign popcount47_ubuz_core_076 = popcount47_ubuz_core_073 ^ popcount47_ubuz_core_075;
  assign popcount47_ubuz_core_078 = input_a[3] & input_a[25];
  assign popcount47_ubuz_core_079 = popcount47_ubuz_core_068 & popcount47_ubuz_core_074;
  assign popcount47_ubuz_core_080 = popcount47_ubuz_core_070 | popcount47_ubuz_core_076;
  assign popcount47_ubuz_core_081 = popcount47_ubuz_core_070 & popcount47_ubuz_core_076;
  assign popcount47_ubuz_core_083 = popcount47_ubuz_core_080 & popcount47_ubuz_core_079;
  assign popcount47_ubuz_core_084 = popcount47_ubuz_core_081 | popcount47_ubuz_core_083;
  assign popcount47_ubuz_core_088 = ~(input_a[25] & input_a[0]);
  assign popcount47_ubuz_core_089 = input_a[41] ^ input_a[34];
  assign popcount47_ubuz_core_099_not = ~popcount47_ubuz_core_084;
  assign popcount47_ubuz_core_103 = input_a[34] ^ input_a[6];
  assign popcount47_ubuz_core_106 = ~(input_a[0] & input_a[34]);
  assign popcount47_ubuz_core_107 = ~(input_a[24] | input_a[2]);
  assign popcount47_ubuz_core_108 = input_a[12] & input_a[35];
  assign popcount47_ubuz_core_110 = input_a[11] & input_a[23];
  assign popcount47_ubuz_core_111 = popcount47_ubuz_core_108 | popcount47_ubuz_core_110;
  assign popcount47_ubuz_core_113 = input_a[15] ^ input_a[16];
  assign popcount47_ubuz_core_114 = input_a[15] & input_a[16];
  assign popcount47_ubuz_core_115 = input_a[14] ^ popcount47_ubuz_core_113;
  assign popcount47_ubuz_core_116 = input_a[14] & popcount47_ubuz_core_113;
  assign popcount47_ubuz_core_117 = popcount47_ubuz_core_114 | popcount47_ubuz_core_116;
  assign popcount47_ubuz_core_118 = ~input_a[20];
  assign popcount47_ubuz_core_119 = input_a[45] | input_a[22];
  assign popcount47_ubuz_core_120 = input_a[4] & popcount47_ubuz_core_115;
  assign popcount47_ubuz_core_121 = popcount47_ubuz_core_111 ^ popcount47_ubuz_core_117;
  assign popcount47_ubuz_core_122 = popcount47_ubuz_core_111 & popcount47_ubuz_core_117;
  assign popcount47_ubuz_core_123 = popcount47_ubuz_core_121 ^ popcount47_ubuz_core_120;
  assign popcount47_ubuz_core_124 = popcount47_ubuz_core_121 & popcount47_ubuz_core_120;
  assign popcount47_ubuz_core_125 = popcount47_ubuz_core_122 | popcount47_ubuz_core_124;
  assign popcount47_ubuz_core_127 = input_a[29] ^ input_a[35];
  assign popcount47_ubuz_core_129 = ~input_a[29];
  assign popcount47_ubuz_core_131 = input_a[18] ^ input_a[19];
  assign popcount47_ubuz_core_132 = input_a[18] & input_a[19];
  assign popcount47_ubuz_core_133 = input_a[17] ^ popcount47_ubuz_core_131;
  assign popcount47_ubuz_core_134 = input_a[17] & popcount47_ubuz_core_131;
  assign popcount47_ubuz_core_135 = popcount47_ubuz_core_132 | popcount47_ubuz_core_134;
  assign popcount47_ubuz_core_136 = ~(input_a[43] | input_a[18]);
  assign popcount47_ubuz_core_137 = input_a[21] ^ input_a[22];
  assign popcount47_ubuz_core_138 = input_a[21] & input_a[22];
  assign popcount47_ubuz_core_139 = input_a[20] ^ popcount47_ubuz_core_137;
  assign popcount47_ubuz_core_140 = input_a[20] & popcount47_ubuz_core_137;
  assign popcount47_ubuz_core_141 = popcount47_ubuz_core_138 | popcount47_ubuz_core_140;
  assign popcount47_ubuz_core_142 = ~(input_a[38] & input_a[20]);
  assign popcount47_ubuz_core_143 = popcount47_ubuz_core_133 ^ popcount47_ubuz_core_139;
  assign popcount47_ubuz_core_144 = popcount47_ubuz_core_133 & popcount47_ubuz_core_139;
  assign popcount47_ubuz_core_145 = popcount47_ubuz_core_135 ^ popcount47_ubuz_core_141;
  assign popcount47_ubuz_core_146 = popcount47_ubuz_core_135 & popcount47_ubuz_core_141;
  assign popcount47_ubuz_core_147 = popcount47_ubuz_core_145 ^ popcount47_ubuz_core_144;
  assign popcount47_ubuz_core_148 = popcount47_ubuz_core_145 & popcount47_ubuz_core_144;
  assign popcount47_ubuz_core_149 = popcount47_ubuz_core_146 | popcount47_ubuz_core_148;
  assign popcount47_ubuz_core_151 = input_a[22] ^ input_a[10];
  assign popcount47_ubuz_core_153 = ~(input_a[16] ^ input_a[22]);
  assign popcount47_ubuz_core_154 = ~(input_a[21] & input_a[15]);
  assign popcount47_ubuz_core_155 = ~(input_a[39] | input_a[21]);
  assign popcount47_ubuz_core_156 = input_a[39] & popcount47_ubuz_core_143;
  assign popcount47_ubuz_core_157 = popcount47_ubuz_core_123 ^ popcount47_ubuz_core_147;
  assign popcount47_ubuz_core_158 = popcount47_ubuz_core_123 & popcount47_ubuz_core_147;
  assign popcount47_ubuz_core_159 = popcount47_ubuz_core_157 ^ popcount47_ubuz_core_156;
  assign popcount47_ubuz_core_160 = popcount47_ubuz_core_157 & popcount47_ubuz_core_156;
  assign popcount47_ubuz_core_161 = popcount47_ubuz_core_158 | popcount47_ubuz_core_160;
  assign popcount47_ubuz_core_162 = popcount47_ubuz_core_125 ^ popcount47_ubuz_core_149;
  assign popcount47_ubuz_core_163 = popcount47_ubuz_core_125 & popcount47_ubuz_core_149;
  assign popcount47_ubuz_core_164 = popcount47_ubuz_core_162 ^ popcount47_ubuz_core_161;
  assign popcount47_ubuz_core_165 = popcount47_ubuz_core_162 & popcount47_ubuz_core_161;
  assign popcount47_ubuz_core_166 = popcount47_ubuz_core_163 | popcount47_ubuz_core_165;
  assign popcount47_ubuz_core_170 = ~input_a[39];
  assign popcount47_ubuz_core_171 = input_a[6] ^ input_a[42];
  assign popcount47_ubuz_core_172 = input_a[5] & input_a[30];
  assign popcount47_ubuz_core_173 = ~(input_a[24] & input_a[25]);
  assign popcount47_ubuz_core_176 = ~(popcount47_ubuz_core_159 & popcount47_ubuz_core_173);
  assign popcount47_ubuz_core_177 = popcount47_ubuz_core_159 & popcount47_ubuz_core_173;
  assign popcount47_ubuz_core_179 = popcount47_ubuz_core_099_not ^ popcount47_ubuz_core_164;
  assign popcount47_ubuz_core_180 = popcount47_ubuz_core_099_not & popcount47_ubuz_core_164;
  assign popcount47_ubuz_core_181 = popcount47_ubuz_core_179 ^ popcount47_ubuz_core_177;
  assign popcount47_ubuz_core_182 = popcount47_ubuz_core_179 & popcount47_ubuz_core_177;
  assign popcount47_ubuz_core_183 = popcount47_ubuz_core_180 | popcount47_ubuz_core_182;
  assign popcount47_ubuz_core_184 = popcount47_ubuz_core_084 ^ popcount47_ubuz_core_166;
  assign popcount47_ubuz_core_185 = popcount47_ubuz_core_084 & popcount47_ubuz_core_166;
  assign popcount47_ubuz_core_186 = popcount47_ubuz_core_184 ^ popcount47_ubuz_core_183;
  assign popcount47_ubuz_core_187 = popcount47_ubuz_core_184 & popcount47_ubuz_core_183;
  assign popcount47_ubuz_core_188 = popcount47_ubuz_core_185 | popcount47_ubuz_core_187;
  assign popcount47_ubuz_core_190 = input_a[14] ^ input_a[28];
  assign popcount47_ubuz_core_193 = input_a[21] | input_a[5];
  assign popcount47_ubuz_core_194 = ~(input_a[23] | input_a[24]);
  assign popcount47_ubuz_core_195 = ~(input_a[4] & input_a[33]);
  assign popcount47_ubuz_core_199 = ~(input_a[28] & input_a[36]);
  assign popcount47_ubuz_core_200 = input_a[27] ^ input_a[28];
  assign popcount47_ubuz_core_201 = input_a[27] & input_a[28];
  assign popcount47_ubuz_core_202 = input_a[26] ^ popcount47_ubuz_core_200;
  assign popcount47_ubuz_core_203 = input_a[26] & popcount47_ubuz_core_200;
  assign popcount47_ubuz_core_204 = popcount47_ubuz_core_201 | popcount47_ubuz_core_203;
  assign popcount47_ubuz_core_205 = input_a[12] ^ input_a[0];
  assign popcount47_ubuz_core_207 = input_a[43] & popcount47_ubuz_core_202;
  assign popcount47_ubuz_core_210 = popcount47_ubuz_core_204 ^ popcount47_ubuz_core_207;
  assign popcount47_ubuz_core_211 = popcount47_ubuz_core_204 & popcount47_ubuz_core_207;
  assign popcount47_ubuz_core_216 = ~(input_a[4] ^ input_a[23]);
  assign popcount47_ubuz_core_218 = input_a[30] ^ input_a[31];
  assign popcount47_ubuz_core_219 = input_a[30] & input_a[31];
  assign popcount47_ubuz_core_220 = input_a[29] ^ popcount47_ubuz_core_218;
  assign popcount47_ubuz_core_221 = input_a[29] & popcount47_ubuz_core_218;
  assign popcount47_ubuz_core_222 = popcount47_ubuz_core_219 | popcount47_ubuz_core_221;
  assign popcount47_ubuz_core_223 = ~(input_a[36] | input_a[24]);
  assign popcount47_ubuz_core_224 = ~input_a[25];
  assign popcount47_ubuz_core_225 = input_a[33] & input_a[34];
  assign popcount47_ubuz_core_226 = input_a[13] & input_a[4];
  assign popcount47_ubuz_core_227 = input_a[10] ^ input_a[3];
  assign popcount47_ubuz_core_230 = ~popcount47_ubuz_core_220;
  assign popcount47_ubuz_core_232 = popcount47_ubuz_core_222 ^ popcount47_ubuz_core_225;
  assign popcount47_ubuz_core_233 = popcount47_ubuz_core_222 & popcount47_ubuz_core_225;
  assign popcount47_ubuz_core_234 = popcount47_ubuz_core_232 ^ popcount47_ubuz_core_220;
  assign popcount47_ubuz_core_235 = popcount47_ubuz_core_232 & popcount47_ubuz_core_220;
  assign popcount47_ubuz_core_236 = popcount47_ubuz_core_233 | popcount47_ubuz_core_235;
  assign popcount47_ubuz_core_238 = input_a[1] & input_a[18];
  assign popcount47_ubuz_core_240 = input_a[19] | input_a[38];
  assign popcount47_ubuz_core_241 = input_a[34] ^ input_a[26];
  assign popcount47_ubuz_core_243 = input_a[3] & popcount47_ubuz_core_230;
  assign popcount47_ubuz_core_244 = popcount47_ubuz_core_210 ^ popcount47_ubuz_core_234;
  assign popcount47_ubuz_core_245 = popcount47_ubuz_core_210 & popcount47_ubuz_core_234;
  assign popcount47_ubuz_core_246 = popcount47_ubuz_core_244 ^ popcount47_ubuz_core_243;
  assign popcount47_ubuz_core_247 = popcount47_ubuz_core_244 & popcount47_ubuz_core_243;
  assign popcount47_ubuz_core_248 = popcount47_ubuz_core_245 | popcount47_ubuz_core_247;
  assign popcount47_ubuz_core_249 = popcount47_ubuz_core_211 ^ popcount47_ubuz_core_236;
  assign popcount47_ubuz_core_250 = popcount47_ubuz_core_211 & popcount47_ubuz_core_236;
  assign popcount47_ubuz_core_251 = popcount47_ubuz_core_249 ^ popcount47_ubuz_core_248;
  assign popcount47_ubuz_core_252 = popcount47_ubuz_core_249 & popcount47_ubuz_core_248;
  assign popcount47_ubuz_core_253 = popcount47_ubuz_core_250 | popcount47_ubuz_core_252;
  assign popcount47_ubuz_core_255 = input_a[42] & input_a[42];
  assign popcount47_ubuz_core_260 = input_a[36] & input_a[46];
  assign popcount47_ubuz_core_269 = ~(input_a[1] & input_a[32]);
  assign popcount47_ubuz_core_270 = input_a[1] & input_a[32];
  assign popcount47_ubuz_core_272 = input_a[37] & input_a[40];
  assign popcount47_ubuz_core_273 = popcount47_ubuz_core_260 ^ popcount47_ubuz_core_269;
  assign popcount47_ubuz_core_274 = popcount47_ubuz_core_260 & popcount47_ubuz_core_269;
  assign popcount47_ubuz_core_275 = popcount47_ubuz_core_273 ^ popcount47_ubuz_core_272;
  assign popcount47_ubuz_core_276 = popcount47_ubuz_core_273 & popcount47_ubuz_core_272;
  assign popcount47_ubuz_core_277 = popcount47_ubuz_core_274 | popcount47_ubuz_core_276;
  assign popcount47_ubuz_core_280 = popcount47_ubuz_core_270 ^ popcount47_ubuz_core_277;
  assign popcount47_ubuz_core_281 = popcount47_ubuz_core_270 & popcount47_ubuz_core_277;
  assign popcount47_ubuz_core_283 = input_a[15] & input_a[13];
  assign popcount47_ubuz_core_284 = input_a[42] & input_a[45];
  assign popcount47_ubuz_core_285 = ~(input_a[6] & input_a[28]);
  assign popcount47_ubuz_core_286 = input_a[41] & input_a[0];
  assign popcount47_ubuz_core_287 = popcount47_ubuz_core_284 | popcount47_ubuz_core_286;
  assign popcount47_ubuz_core_288 = ~input_a[6];
  assign popcount47_ubuz_core_289 = input_a[29] ^ input_a[31];
  assign popcount47_ubuz_core_291 = ~(input_a[6] ^ input_a[24]);
  assign popcount47_ubuz_core_292 = input_a[41] ^ input_a[44];
  assign popcount47_ubuz_core_293 = ~(input_a[28] | input_a[29]);
  assign popcount47_ubuz_core_295 = input_a[26] | input_a[6];
  assign popcount47_ubuz_core_296 = ~input_a[9];
  assign popcount47_ubuz_core_298 = ~(input_a[9] | input_a[36]);
  assign popcount47_ubuz_core_301 = ~(input_a[1] | input_a[35]);
  assign popcount47_ubuz_core_304 = input_a[35] ^ input_a[9];
  assign popcount47_ubuz_core_307 = ~(input_a[36] & input_a[24]);
  assign popcount47_ubuz_core_309 = popcount47_ubuz_core_275 ^ popcount47_ubuz_core_287;
  assign popcount47_ubuz_core_310 = popcount47_ubuz_core_275 & popcount47_ubuz_core_287;
  assign popcount47_ubuz_core_316 = popcount47_ubuz_core_280 ^ popcount47_ubuz_core_310;
  assign popcount47_ubuz_core_317 = popcount47_ubuz_core_280 & popcount47_ubuz_core_310;
  assign popcount47_ubuz_core_321 = popcount47_ubuz_core_281 | popcount47_ubuz_core_317;
  assign popcount47_ubuz_core_322 = input_a[36] & input_a[41];
  assign popcount47_ubuz_core_323 = ~(input_a[17] & input_a[18]);
  assign popcount47_ubuz_core_325 = input_a[44] & input_a[44];
  assign popcount47_ubuz_core_326 = popcount47_ubuz_core_246 ^ popcount47_ubuz_core_309;
  assign popcount47_ubuz_core_327 = popcount47_ubuz_core_246 & popcount47_ubuz_core_309;
  assign popcount47_ubuz_core_328 = popcount47_ubuz_core_326 ^ input_a[44];
  assign popcount47_ubuz_core_329 = popcount47_ubuz_core_326 & popcount47_ubuz_core_325;
  assign popcount47_ubuz_core_330 = popcount47_ubuz_core_327 | popcount47_ubuz_core_329;
  assign popcount47_ubuz_core_331 = popcount47_ubuz_core_251 ^ popcount47_ubuz_core_316;
  assign popcount47_ubuz_core_332 = popcount47_ubuz_core_251 & popcount47_ubuz_core_316;
  assign popcount47_ubuz_core_333 = popcount47_ubuz_core_331 ^ popcount47_ubuz_core_330;
  assign popcount47_ubuz_core_334 = popcount47_ubuz_core_331 & popcount47_ubuz_core_330;
  assign popcount47_ubuz_core_335 = popcount47_ubuz_core_332 | popcount47_ubuz_core_334;
  assign popcount47_ubuz_core_336 = popcount47_ubuz_core_253 ^ popcount47_ubuz_core_321;
  assign popcount47_ubuz_core_337 = popcount47_ubuz_core_253 & popcount47_ubuz_core_321;
  assign popcount47_ubuz_core_338 = popcount47_ubuz_core_336 ^ popcount47_ubuz_core_335;
  assign popcount47_ubuz_core_339 = popcount47_ubuz_core_336 & popcount47_ubuz_core_335;
  assign popcount47_ubuz_core_340 = popcount47_ubuz_core_337 | popcount47_ubuz_core_339;
  assign popcount47_ubuz_core_344 = input_a[3] | input_a[35];
  assign popcount47_ubuz_core_345 = ~(input_a[36] ^ input_a[43]);
  assign popcount47_ubuz_core_347 = input_a[25] & input_a[24];
  assign popcount47_ubuz_core_348 = popcount47_ubuz_core_176 ^ popcount47_ubuz_core_328;
  assign popcount47_ubuz_core_349 = popcount47_ubuz_core_176 & popcount47_ubuz_core_328;
  assign popcount47_ubuz_core_350 = popcount47_ubuz_core_348 ^ popcount47_ubuz_core_347;
  assign popcount47_ubuz_core_351 = popcount47_ubuz_core_348 & popcount47_ubuz_core_347;
  assign popcount47_ubuz_core_352 = popcount47_ubuz_core_349 | popcount47_ubuz_core_351;
  assign popcount47_ubuz_core_353 = popcount47_ubuz_core_181 ^ popcount47_ubuz_core_333;
  assign popcount47_ubuz_core_354 = popcount47_ubuz_core_181 & popcount47_ubuz_core_333;
  assign popcount47_ubuz_core_355 = popcount47_ubuz_core_353 ^ popcount47_ubuz_core_352;
  assign popcount47_ubuz_core_356 = popcount47_ubuz_core_353 & popcount47_ubuz_core_352;
  assign popcount47_ubuz_core_357 = popcount47_ubuz_core_354 | popcount47_ubuz_core_356;
  assign popcount47_ubuz_core_358 = popcount47_ubuz_core_186 ^ popcount47_ubuz_core_338;
  assign popcount47_ubuz_core_359 = popcount47_ubuz_core_186 & popcount47_ubuz_core_338;
  assign popcount47_ubuz_core_360 = popcount47_ubuz_core_358 ^ popcount47_ubuz_core_357;
  assign popcount47_ubuz_core_361 = popcount47_ubuz_core_358 & popcount47_ubuz_core_357;
  assign popcount47_ubuz_core_362 = popcount47_ubuz_core_359 | popcount47_ubuz_core_361;
  assign popcount47_ubuz_core_363 = popcount47_ubuz_core_188 ^ popcount47_ubuz_core_340;
  assign popcount47_ubuz_core_364 = popcount47_ubuz_core_188 & popcount47_ubuz_core_340;
  assign popcount47_ubuz_core_365 = popcount47_ubuz_core_363 ^ popcount47_ubuz_core_362;
  assign popcount47_ubuz_core_366 = popcount47_ubuz_core_363 & popcount47_ubuz_core_362;
  assign popcount47_ubuz_core_367 = popcount47_ubuz_core_364 | popcount47_ubuz_core_366;
  assign popcount47_ubuz_core_369 = ~(input_a[46] | input_a[42]);
  assign popcount47_ubuz_core_372 = input_a[42] & input_a[4];

  assign popcount47_ubuz_out[0] = input_a[38];
  assign popcount47_ubuz_out[1] = popcount47_ubuz_core_350;
  assign popcount47_ubuz_out[2] = popcount47_ubuz_core_355;
  assign popcount47_ubuz_out[3] = popcount47_ubuz_core_360;
  assign popcount47_ubuz_out[4] = popcount47_ubuz_core_365;
  assign popcount47_ubuz_out[5] = popcount47_ubuz_core_367;
endmodule