// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=0.5
// WCE=1.0
// EP=0.5%
// Printed PDK parameters:
//  Area=81505128.0
//  Delay=69646880.0
//  Power=4604300.0

module popcount27_3ii0(input [26:0] input_a, output [4:0] popcount27_3ii0_out);
  wire popcount27_3ii0_core_029;
  wire popcount27_3ii0_core_030;
  wire popcount27_3ii0_core_031;
  wire popcount27_3ii0_core_032;
  wire popcount27_3ii0_core_033;
  wire popcount27_3ii0_core_034;
  wire popcount27_3ii0_core_035;
  wire popcount27_3ii0_core_036;
  wire popcount27_3ii0_core_037;
  wire popcount27_3ii0_core_038;
  wire popcount27_3ii0_core_039;
  wire popcount27_3ii0_core_041;
  wire popcount27_3ii0_core_042;
  wire popcount27_3ii0_core_043;
  wire popcount27_3ii0_core_044;
  wire popcount27_3ii0_core_045;
  wire popcount27_3ii0_core_046;
  wire popcount27_3ii0_core_047;
  wire popcount27_3ii0_core_049;
  wire popcount27_3ii0_core_053;
  wire popcount27_3ii0_core_054;
  wire popcount27_3ii0_core_055;
  wire popcount27_3ii0_core_056;
  wire popcount27_3ii0_core_057;
  wire popcount27_3ii0_core_059;
  wire popcount27_3ii0_core_060;
  wire popcount27_3ii0_core_061;
  wire popcount27_3ii0_core_062;
  wire popcount27_3ii0_core_063;
  wire popcount27_3ii0_core_064;
  wire popcount27_3ii0_core_065;
  wire popcount27_3ii0_core_066;
  wire popcount27_3ii0_core_067;
  wire popcount27_3ii0_core_068;
  wire popcount27_3ii0_core_070;
  wire popcount27_3ii0_core_071;
  wire popcount27_3ii0_core_072;
  wire popcount27_3ii0_core_073;
  wire popcount27_3ii0_core_074;
  wire popcount27_3ii0_core_075;
  wire popcount27_3ii0_core_076;
  wire popcount27_3ii0_core_079;
  wire popcount27_3ii0_core_080;
  wire popcount27_3ii0_core_081;
  wire popcount27_3ii0_core_082;
  wire popcount27_3ii0_core_083;
  wire popcount27_3ii0_core_084;
  wire popcount27_3ii0_core_085;
  wire popcount27_3ii0_core_086;
  wire popcount27_3ii0_core_087;
  wire popcount27_3ii0_core_088;
  wire popcount27_3ii0_core_089;
  wire popcount27_3ii0_core_090;
  wire popcount27_3ii0_core_091;
  wire popcount27_3ii0_core_092;
  wire popcount27_3ii0_core_093;
  wire popcount27_3ii0_core_097;
  wire popcount27_3ii0_core_099;
  wire popcount27_3ii0_core_100;
  wire popcount27_3ii0_core_101;
  wire popcount27_3ii0_core_102;
  wire popcount27_3ii0_core_103;
  wire popcount27_3ii0_core_105;
  wire popcount27_3ii0_core_106;
  wire popcount27_3ii0_core_107;
  wire popcount27_3ii0_core_108;
  wire popcount27_3ii0_core_109;
  wire popcount27_3ii0_core_110;
  wire popcount27_3ii0_core_111;
  wire popcount27_3ii0_core_112;
  wire popcount27_3ii0_core_113;
  wire popcount27_3ii0_core_116;
  wire popcount27_3ii0_core_117;
  wire popcount27_3ii0_core_118;
  wire popcount27_3ii0_core_119;
  wire popcount27_3ii0_core_120;
  wire popcount27_3ii0_core_121;
  wire popcount27_3ii0_core_122;
  wire popcount27_3ii0_core_124;
  wire popcount27_3ii0_core_125;
  wire popcount27_3ii0_core_126;
  wire popcount27_3ii0_core_128;
  wire popcount27_3ii0_core_129;
  wire popcount27_3ii0_core_130;
  wire popcount27_3ii0_core_131;
  wire popcount27_3ii0_core_132;
  wire popcount27_3ii0_core_134;
  wire popcount27_3ii0_core_135;
  wire popcount27_3ii0_core_136;
  wire popcount27_3ii0_core_137;
  wire popcount27_3ii0_core_138;
  wire popcount27_3ii0_core_139;
  wire popcount27_3ii0_core_140;
  wire popcount27_3ii0_core_141;
  wire popcount27_3ii0_core_142;
  wire popcount27_3ii0_core_143;
  wire popcount27_3ii0_core_145;
  wire popcount27_3ii0_core_146;
  wire popcount27_3ii0_core_147;
  wire popcount27_3ii0_core_148;
  wire popcount27_3ii0_core_149;
  wire popcount27_3ii0_core_150;
  wire popcount27_3ii0_core_151;
  wire popcount27_3ii0_core_154;
  wire popcount27_3ii0_core_156;
  wire popcount27_3ii0_core_157;
  wire popcount27_3ii0_core_158;
  wire popcount27_3ii0_core_159;
  wire popcount27_3ii0_core_160;
  wire popcount27_3ii0_core_161;
  wire popcount27_3ii0_core_162;
  wire popcount27_3ii0_core_163;
  wire popcount27_3ii0_core_164;
  wire popcount27_3ii0_core_165;
  wire popcount27_3ii0_core_166;
  wire popcount27_3ii0_core_167;
  wire popcount27_3ii0_core_168;
  wire popcount27_3ii0_core_172;
  wire popcount27_3ii0_core_174;
  wire popcount27_3ii0_core_175;
  wire popcount27_3ii0_core_176;
  wire popcount27_3ii0_core_177;
  wire popcount27_3ii0_core_178;
  wire popcount27_3ii0_core_179;
  wire popcount27_3ii0_core_180;
  wire popcount27_3ii0_core_181;
  wire popcount27_3ii0_core_182;
  wire popcount27_3ii0_core_183;
  wire popcount27_3ii0_core_184;
  wire popcount27_3ii0_core_185;
  wire popcount27_3ii0_core_186;
  wire popcount27_3ii0_core_187;
  wire popcount27_3ii0_core_188;
  wire popcount27_3ii0_core_189;
  wire popcount27_3ii0_core_190;
  wire popcount27_3ii0_core_194;
  wire popcount27_3ii0_core_195;

  assign popcount27_3ii0_core_029 = input_a[1] ^ input_a[2];
  assign popcount27_3ii0_core_030 = input_a[1] & input_a[2];
  assign popcount27_3ii0_core_031 = input_a[0] ^ popcount27_3ii0_core_029;
  assign popcount27_3ii0_core_032 = input_a[0] & popcount27_3ii0_core_029;
  assign popcount27_3ii0_core_033 = popcount27_3ii0_core_030 | popcount27_3ii0_core_032;
  assign popcount27_3ii0_core_034 = input_a[9] | input_a[16];
  assign popcount27_3ii0_core_035 = ~(input_a[4] & input_a[5]);
  assign popcount27_3ii0_core_036 = input_a[4] & input_a[5];
  assign popcount27_3ii0_core_037 = input_a[3] ^ popcount27_3ii0_core_035;
  assign popcount27_3ii0_core_038 = ~(input_a[25] & input_a[3]);
  assign popcount27_3ii0_core_039 = popcount27_3ii0_core_036 | input_a[3];
  assign popcount27_3ii0_core_041 = ~(input_a[23] & input_a[25]);
  assign popcount27_3ii0_core_042 = popcount27_3ii0_core_031 & popcount27_3ii0_core_037;
  assign popcount27_3ii0_core_043 = popcount27_3ii0_core_033 ^ popcount27_3ii0_core_039;
  assign popcount27_3ii0_core_044 = popcount27_3ii0_core_033 & popcount27_3ii0_core_039;
  assign popcount27_3ii0_core_045 = popcount27_3ii0_core_043 ^ popcount27_3ii0_core_042;
  assign popcount27_3ii0_core_046 = popcount27_3ii0_core_043 & popcount27_3ii0_core_042;
  assign popcount27_3ii0_core_047 = popcount27_3ii0_core_044 | popcount27_3ii0_core_046;
  assign popcount27_3ii0_core_049 = input_a[1] | input_a[15];
  assign popcount27_3ii0_core_053 = input_a[7] ^ input_a[8];
  assign popcount27_3ii0_core_054 = input_a[7] & input_a[8];
  assign popcount27_3ii0_core_055 = input_a[6] ^ popcount27_3ii0_core_053;
  assign popcount27_3ii0_core_056 = input_a[6] & popcount27_3ii0_core_053;
  assign popcount27_3ii0_core_057 = popcount27_3ii0_core_054 | popcount27_3ii0_core_056;
  assign popcount27_3ii0_core_059 = input_a[9] ^ input_a[10];
  assign popcount27_3ii0_core_060 = input_a[9] & input_a[10];
  assign popcount27_3ii0_core_061 = input_a[11] ^ input_a[12];
  assign popcount27_3ii0_core_062 = input_a[11] & input_a[12];
  assign popcount27_3ii0_core_063 = popcount27_3ii0_core_059 ^ popcount27_3ii0_core_061;
  assign popcount27_3ii0_core_064 = popcount27_3ii0_core_059 & popcount27_3ii0_core_061;
  assign popcount27_3ii0_core_065 = popcount27_3ii0_core_060 ^ popcount27_3ii0_core_062;
  assign popcount27_3ii0_core_066 = popcount27_3ii0_core_060 & popcount27_3ii0_core_062;
  assign popcount27_3ii0_core_067 = popcount27_3ii0_core_065 | popcount27_3ii0_core_064;
  assign popcount27_3ii0_core_068 = ~(input_a[6] & input_a[25]);
  assign popcount27_3ii0_core_070 = popcount27_3ii0_core_055 ^ popcount27_3ii0_core_063;
  assign popcount27_3ii0_core_071 = popcount27_3ii0_core_055 & popcount27_3ii0_core_063;
  assign popcount27_3ii0_core_072 = popcount27_3ii0_core_057 ^ popcount27_3ii0_core_067;
  assign popcount27_3ii0_core_073 = popcount27_3ii0_core_057 & popcount27_3ii0_core_067;
  assign popcount27_3ii0_core_074 = popcount27_3ii0_core_072 ^ popcount27_3ii0_core_071;
  assign popcount27_3ii0_core_075 = popcount27_3ii0_core_072 & popcount27_3ii0_core_071;
  assign popcount27_3ii0_core_076 = popcount27_3ii0_core_073 | popcount27_3ii0_core_075;
  assign popcount27_3ii0_core_079 = popcount27_3ii0_core_066 | popcount27_3ii0_core_076;
  assign popcount27_3ii0_core_080 = input_a[16] & input_a[11];
  assign popcount27_3ii0_core_081 = ~(input_a[9] ^ input_a[13]);
  assign popcount27_3ii0_core_082 = input_a[5] ^ popcount27_3ii0_core_070;
  assign popcount27_3ii0_core_083 = input_a[5] & popcount27_3ii0_core_070;
  assign popcount27_3ii0_core_084 = popcount27_3ii0_core_045 ^ popcount27_3ii0_core_074;
  assign popcount27_3ii0_core_085 = popcount27_3ii0_core_045 & popcount27_3ii0_core_074;
  assign popcount27_3ii0_core_086 = popcount27_3ii0_core_084 ^ popcount27_3ii0_core_083;
  assign popcount27_3ii0_core_087 = popcount27_3ii0_core_084 & popcount27_3ii0_core_083;
  assign popcount27_3ii0_core_088 = popcount27_3ii0_core_085 | popcount27_3ii0_core_087;
  assign popcount27_3ii0_core_089 = popcount27_3ii0_core_047 ^ popcount27_3ii0_core_079;
  assign popcount27_3ii0_core_090 = popcount27_3ii0_core_047 & popcount27_3ii0_core_079;
  assign popcount27_3ii0_core_091 = popcount27_3ii0_core_089 ^ popcount27_3ii0_core_088;
  assign popcount27_3ii0_core_092 = popcount27_3ii0_core_089 & popcount27_3ii0_core_088;
  assign popcount27_3ii0_core_093 = popcount27_3ii0_core_090 | popcount27_3ii0_core_092;
  assign popcount27_3ii0_core_097 = ~(input_a[4] & input_a[5]);
  assign popcount27_3ii0_core_099 = input_a[14] ^ input_a[15];
  assign popcount27_3ii0_core_100 = input_a[14] & input_a[15];
  assign popcount27_3ii0_core_101 = input_a[13] ^ popcount27_3ii0_core_099;
  assign popcount27_3ii0_core_102 = input_a[13] & popcount27_3ii0_core_099;
  assign popcount27_3ii0_core_103 = popcount27_3ii0_core_100 | popcount27_3ii0_core_102;
  assign popcount27_3ii0_core_105 = input_a[16] ^ input_a[17];
  assign popcount27_3ii0_core_106 = input_a[16] & input_a[17];
  assign popcount27_3ii0_core_107 = input_a[18] ^ input_a[19];
  assign popcount27_3ii0_core_108 = input_a[18] & input_a[19];
  assign popcount27_3ii0_core_109 = popcount27_3ii0_core_105 ^ popcount27_3ii0_core_107;
  assign popcount27_3ii0_core_110 = popcount27_3ii0_core_105 & popcount27_3ii0_core_107;
  assign popcount27_3ii0_core_111 = popcount27_3ii0_core_106 ^ popcount27_3ii0_core_108;
  assign popcount27_3ii0_core_112 = popcount27_3ii0_core_106 & popcount27_3ii0_core_108;
  assign popcount27_3ii0_core_113 = popcount27_3ii0_core_111 | popcount27_3ii0_core_110;
  assign popcount27_3ii0_core_116 = popcount27_3ii0_core_101 ^ popcount27_3ii0_core_109;
  assign popcount27_3ii0_core_117 = popcount27_3ii0_core_101 & popcount27_3ii0_core_109;
  assign popcount27_3ii0_core_118 = popcount27_3ii0_core_103 ^ popcount27_3ii0_core_113;
  assign popcount27_3ii0_core_119 = popcount27_3ii0_core_103 & popcount27_3ii0_core_113;
  assign popcount27_3ii0_core_120 = popcount27_3ii0_core_118 ^ popcount27_3ii0_core_117;
  assign popcount27_3ii0_core_121 = popcount27_3ii0_core_118 & popcount27_3ii0_core_117;
  assign popcount27_3ii0_core_122 = popcount27_3ii0_core_119 | popcount27_3ii0_core_121;
  assign popcount27_3ii0_core_124 = ~(input_a[16] & input_a[19]);
  assign popcount27_3ii0_core_125 = popcount27_3ii0_core_112 | popcount27_3ii0_core_122;
  assign popcount27_3ii0_core_126 = input_a[1] ^ input_a[21];
  assign popcount27_3ii0_core_128 = input_a[21] ^ input_a[22];
  assign popcount27_3ii0_core_129 = input_a[21] & input_a[22];
  assign popcount27_3ii0_core_130 = input_a[20] ^ popcount27_3ii0_core_128;
  assign popcount27_3ii0_core_131 = input_a[20] & popcount27_3ii0_core_128;
  assign popcount27_3ii0_core_132 = popcount27_3ii0_core_129 | popcount27_3ii0_core_131;
  assign popcount27_3ii0_core_134 = input_a[23] ^ input_a[24];
  assign popcount27_3ii0_core_135 = input_a[23] & input_a[24];
  assign popcount27_3ii0_core_136 = input_a[25] ^ input_a[26];
  assign popcount27_3ii0_core_137 = input_a[25] & input_a[26];
  assign popcount27_3ii0_core_138 = popcount27_3ii0_core_134 ^ popcount27_3ii0_core_136;
  assign popcount27_3ii0_core_139 = popcount27_3ii0_core_134 & popcount27_3ii0_core_136;
  assign popcount27_3ii0_core_140 = popcount27_3ii0_core_135 ^ popcount27_3ii0_core_137;
  assign popcount27_3ii0_core_141 = popcount27_3ii0_core_135 & popcount27_3ii0_core_137;
  assign popcount27_3ii0_core_142 = popcount27_3ii0_core_140 | popcount27_3ii0_core_139;
  assign popcount27_3ii0_core_143 = input_a[18] ^ input_a[17];
  assign popcount27_3ii0_core_145 = popcount27_3ii0_core_130 ^ popcount27_3ii0_core_138;
  assign popcount27_3ii0_core_146 = popcount27_3ii0_core_130 & popcount27_3ii0_core_138;
  assign popcount27_3ii0_core_147 = popcount27_3ii0_core_132 ^ popcount27_3ii0_core_142;
  assign popcount27_3ii0_core_148 = popcount27_3ii0_core_132 & popcount27_3ii0_core_142;
  assign popcount27_3ii0_core_149 = popcount27_3ii0_core_147 ^ popcount27_3ii0_core_146;
  assign popcount27_3ii0_core_150 = popcount27_3ii0_core_147 & popcount27_3ii0_core_146;
  assign popcount27_3ii0_core_151 = popcount27_3ii0_core_148 | popcount27_3ii0_core_150;
  assign popcount27_3ii0_core_154 = popcount27_3ii0_core_141 | popcount27_3ii0_core_151;
  assign popcount27_3ii0_core_156 = input_a[7] ^ input_a[25];
  assign popcount27_3ii0_core_157 = popcount27_3ii0_core_116 ^ popcount27_3ii0_core_145;
  assign popcount27_3ii0_core_158 = popcount27_3ii0_core_116 & popcount27_3ii0_core_145;
  assign popcount27_3ii0_core_159 = popcount27_3ii0_core_120 ^ popcount27_3ii0_core_149;
  assign popcount27_3ii0_core_160 = popcount27_3ii0_core_120 & popcount27_3ii0_core_149;
  assign popcount27_3ii0_core_161 = popcount27_3ii0_core_159 ^ popcount27_3ii0_core_158;
  assign popcount27_3ii0_core_162 = popcount27_3ii0_core_159 & popcount27_3ii0_core_158;
  assign popcount27_3ii0_core_163 = popcount27_3ii0_core_160 | popcount27_3ii0_core_162;
  assign popcount27_3ii0_core_164 = popcount27_3ii0_core_125 ^ popcount27_3ii0_core_154;
  assign popcount27_3ii0_core_165 = popcount27_3ii0_core_125 & popcount27_3ii0_core_154;
  assign popcount27_3ii0_core_166 = popcount27_3ii0_core_164 ^ popcount27_3ii0_core_163;
  assign popcount27_3ii0_core_167 = popcount27_3ii0_core_164 & popcount27_3ii0_core_163;
  assign popcount27_3ii0_core_168 = popcount27_3ii0_core_165 | popcount27_3ii0_core_167;
  assign popcount27_3ii0_core_172 = input_a[19] | input_a[10];
  assign popcount27_3ii0_core_174 = popcount27_3ii0_core_082 ^ popcount27_3ii0_core_157;
  assign popcount27_3ii0_core_175 = popcount27_3ii0_core_082 & popcount27_3ii0_core_157;
  assign popcount27_3ii0_core_176 = popcount27_3ii0_core_086 ^ popcount27_3ii0_core_161;
  assign popcount27_3ii0_core_177 = popcount27_3ii0_core_086 & popcount27_3ii0_core_161;
  assign popcount27_3ii0_core_178 = popcount27_3ii0_core_176 ^ popcount27_3ii0_core_175;
  assign popcount27_3ii0_core_179 = popcount27_3ii0_core_176 & popcount27_3ii0_core_175;
  assign popcount27_3ii0_core_180 = popcount27_3ii0_core_177 | popcount27_3ii0_core_179;
  assign popcount27_3ii0_core_181 = popcount27_3ii0_core_091 ^ popcount27_3ii0_core_166;
  assign popcount27_3ii0_core_182 = popcount27_3ii0_core_091 & popcount27_3ii0_core_166;
  assign popcount27_3ii0_core_183 = popcount27_3ii0_core_181 ^ popcount27_3ii0_core_180;
  assign popcount27_3ii0_core_184 = popcount27_3ii0_core_181 & popcount27_3ii0_core_180;
  assign popcount27_3ii0_core_185 = popcount27_3ii0_core_182 | popcount27_3ii0_core_184;
  assign popcount27_3ii0_core_186 = popcount27_3ii0_core_093 ^ popcount27_3ii0_core_168;
  assign popcount27_3ii0_core_187 = popcount27_3ii0_core_093 & popcount27_3ii0_core_168;
  assign popcount27_3ii0_core_188 = popcount27_3ii0_core_186 ^ popcount27_3ii0_core_185;
  assign popcount27_3ii0_core_189 = popcount27_3ii0_core_186 & popcount27_3ii0_core_185;
  assign popcount27_3ii0_core_190 = popcount27_3ii0_core_187 | popcount27_3ii0_core_189;
  assign popcount27_3ii0_core_194 = ~(input_a[20] ^ input_a[9]);
  assign popcount27_3ii0_core_195 = input_a[21] & input_a[18];

  assign popcount27_3ii0_out[0] = popcount27_3ii0_core_174;
  assign popcount27_3ii0_out[1] = popcount27_3ii0_core_178;
  assign popcount27_3ii0_out[2] = popcount27_3ii0_core_183;
  assign popcount27_3ii0_out[3] = popcount27_3ii0_core_188;
  assign popcount27_3ii0_out[4] = popcount27_3ii0_core_190;
endmodule