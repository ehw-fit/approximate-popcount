// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.46738
// WCE=6.0
// EP=0.792892%
// Printed PDK parameters:
//  Area=47898478.0
//  Delay=64143948.0
//  Power=2330500.0

module popcount28_b7nj(input [27:0] input_a, output [4:0] popcount28_b7nj_out);
  wire popcount28_b7nj_core_030;
  wire popcount28_b7nj_core_031;
  wire popcount28_b7nj_core_033;
  wire popcount28_b7nj_core_035;
  wire popcount28_b7nj_core_037;
  wire popcount28_b7nj_core_038;
  wire popcount28_b7nj_core_039;
  wire popcount28_b7nj_core_040;
  wire popcount28_b7nj_core_041;
  wire popcount28_b7nj_core_042;
  wire popcount28_b7nj_core_044;
  wire popcount28_b7nj_core_045;
  wire popcount28_b7nj_core_046;
  wire popcount28_b7nj_core_047;
  wire popcount28_b7nj_core_048;
  wire popcount28_b7nj_core_054;
  wire popcount28_b7nj_core_056;
  wire popcount28_b7nj_core_057;
  wire popcount28_b7nj_core_059;
  wire popcount28_b7nj_core_060;
  wire popcount28_b7nj_core_061;
  wire popcount28_b7nj_core_062;
  wire popcount28_b7nj_core_063;
  wire popcount28_b7nj_core_065;
  wire popcount28_b7nj_core_066;
  wire popcount28_b7nj_core_067;
  wire popcount28_b7nj_core_068;
  wire popcount28_b7nj_core_069;
  wire popcount28_b7nj_core_070;
  wire popcount28_b7nj_core_071;
  wire popcount28_b7nj_core_072;
  wire popcount28_b7nj_core_073;
  wire popcount28_b7nj_core_074;
  wire popcount28_b7nj_core_076;
  wire popcount28_b7nj_core_077;
  wire popcount28_b7nj_core_078;
  wire popcount28_b7nj_core_079;
  wire popcount28_b7nj_core_080;
  wire popcount28_b7nj_core_081;
  wire popcount28_b7nj_core_082;
  wire popcount28_b7nj_core_085;
  wire popcount28_b7nj_core_086;
  wire popcount28_b7nj_core_088;
  wire popcount28_b7nj_core_089;
  wire popcount28_b7nj_core_091;
  wire popcount28_b7nj_core_094;
  wire popcount28_b7nj_core_095;
  wire popcount28_b7nj_core_096;
  wire popcount28_b7nj_core_098;
  wire popcount28_b7nj_core_102;
  wire popcount28_b7nj_core_103;
  wire popcount28_b7nj_core_104;
  wire popcount28_b7nj_core_105;
  wire popcount28_b7nj_core_106;
  wire popcount28_b7nj_core_107;
  wire popcount28_b7nj_core_108;
  wire popcount28_b7nj_core_111;
  wire popcount28_b7nj_core_112;
  wire popcount28_b7nj_core_113;
  wire popcount28_b7nj_core_114;
  wire popcount28_b7nj_core_116;
  wire popcount28_b7nj_core_117;
  wire popcount28_b7nj_core_118;
  wire popcount28_b7nj_core_119;
  wire popcount28_b7nj_core_120;
  wire popcount28_b7nj_core_123;
  wire popcount28_b7nj_core_124;
  wire popcount28_b7nj_core_125;
  wire popcount28_b7nj_core_130;
  wire popcount28_b7nj_core_131;
  wire popcount28_b7nj_core_132;
  wire popcount28_b7nj_core_133;
  wire popcount28_b7nj_core_135;
  wire popcount28_b7nj_core_137;
  wire popcount28_b7nj_core_138;
  wire popcount28_b7nj_core_140;
  wire popcount28_b7nj_core_141;
  wire popcount28_b7nj_core_142;
  wire popcount28_b7nj_core_143;
  wire popcount28_b7nj_core_144;
  wire popcount28_b7nj_core_145;
  wire popcount28_b7nj_core_146;
  wire popcount28_b7nj_core_147;
  wire popcount28_b7nj_core_148;
  wire popcount28_b7nj_core_149;
  wire popcount28_b7nj_core_150;
  wire popcount28_b7nj_core_151;
  wire popcount28_b7nj_core_152;
  wire popcount28_b7nj_core_153;
  wire popcount28_b7nj_core_154;
  wire popcount28_b7nj_core_160;
  wire popcount28_b7nj_core_163;
  wire popcount28_b7nj_core_164;
  wire popcount28_b7nj_core_165;
  wire popcount28_b7nj_core_166;
  wire popcount28_b7nj_core_167;
  wire popcount28_b7nj_core_168;
  wire popcount28_b7nj_core_169;
  wire popcount28_b7nj_core_170;
  wire popcount28_b7nj_core_171;
  wire popcount28_b7nj_core_172;
  wire popcount28_b7nj_core_173;
  wire popcount28_b7nj_core_174;
  wire popcount28_b7nj_core_176;
  wire popcount28_b7nj_core_178;
  wire popcount28_b7nj_core_179;
  wire popcount28_b7nj_core_180;
  wire popcount28_b7nj_core_181;
  wire popcount28_b7nj_core_182;
  wire popcount28_b7nj_core_183;
  wire popcount28_b7nj_core_184;
  wire popcount28_b7nj_core_185;
  wire popcount28_b7nj_core_186;
  wire popcount28_b7nj_core_187;
  wire popcount28_b7nj_core_188;
  wire popcount28_b7nj_core_189;
  wire popcount28_b7nj_core_190;
  wire popcount28_b7nj_core_191;
  wire popcount28_b7nj_core_192;
  wire popcount28_b7nj_core_193;
  wire popcount28_b7nj_core_194;
  wire popcount28_b7nj_core_195;
  wire popcount28_b7nj_core_196;
  wire popcount28_b7nj_core_197;
  wire popcount28_b7nj_core_198;
  wire popcount28_b7nj_core_199;
  wire popcount28_b7nj_core_200;

  assign popcount28_b7nj_core_030 = input_a[11] & input_a[14];
  assign popcount28_b7nj_core_031 = input_a[9] ^ input_a[9];
  assign popcount28_b7nj_core_033 = ~(input_a[20] ^ input_a[7]);
  assign popcount28_b7nj_core_035 = ~(input_a[24] | input_a[3]);
  assign popcount28_b7nj_core_037 = input_a[15] & input_a[0];
  assign popcount28_b7nj_core_038 = ~(input_a[4] ^ input_a[21]);
  assign popcount28_b7nj_core_039 = input_a[5] & input_a[6];
  assign popcount28_b7nj_core_040 = ~input_a[21];
  assign popcount28_b7nj_core_041 = input_a[19] & input_a[2];
  assign popcount28_b7nj_core_042 = ~(input_a[2] & popcount28_b7nj_core_039);
  assign popcount28_b7nj_core_044 = ~popcount28_b7nj_core_042;
  assign popcount28_b7nj_core_045 = ~(input_a[5] ^ input_a[4]);
  assign popcount28_b7nj_core_046 = ~(input_a[3] | input_a[3]);
  assign popcount28_b7nj_core_047 = ~(input_a[27] ^ input_a[22]);
  assign popcount28_b7nj_core_048 = ~input_a[8];
  assign popcount28_b7nj_core_054 = ~(input_a[3] & input_a[22]);
  assign popcount28_b7nj_core_056 = ~(input_a[3] & popcount28_b7nj_core_044);
  assign popcount28_b7nj_core_057 = input_a[3] & popcount28_b7nj_core_044;
  assign popcount28_b7nj_core_059 = input_a[8] ^ input_a[9];
  assign popcount28_b7nj_core_060 = input_a[8] & input_a[9];
  assign popcount28_b7nj_core_061 = input_a[7] ^ popcount28_b7nj_core_059;
  assign popcount28_b7nj_core_062 = input_a[7] & popcount28_b7nj_core_059;
  assign popcount28_b7nj_core_063 = popcount28_b7nj_core_060 | popcount28_b7nj_core_062;
  assign popcount28_b7nj_core_065 = input_a[10] ^ input_a[11];
  assign popcount28_b7nj_core_066 = input_a[10] & input_a[11];
  assign popcount28_b7nj_core_067 = input_a[12] ^ input_a[13];
  assign popcount28_b7nj_core_068 = input_a[12] & input_a[13];
  assign popcount28_b7nj_core_069 = popcount28_b7nj_core_065 ^ popcount28_b7nj_core_067;
  assign popcount28_b7nj_core_070 = popcount28_b7nj_core_065 & popcount28_b7nj_core_067;
  assign popcount28_b7nj_core_071 = popcount28_b7nj_core_066 ^ popcount28_b7nj_core_068;
  assign popcount28_b7nj_core_072 = popcount28_b7nj_core_066 & popcount28_b7nj_core_068;
  assign popcount28_b7nj_core_073 = popcount28_b7nj_core_071 | popcount28_b7nj_core_070;
  assign popcount28_b7nj_core_074 = input_a[22] ^ input_a[22];
  assign popcount28_b7nj_core_076 = input_a[23] ^ input_a[7];
  assign popcount28_b7nj_core_077 = popcount28_b7nj_core_061 & popcount28_b7nj_core_069;
  assign popcount28_b7nj_core_078 = popcount28_b7nj_core_063 ^ popcount28_b7nj_core_073;
  assign popcount28_b7nj_core_079 = popcount28_b7nj_core_063 & popcount28_b7nj_core_073;
  assign popcount28_b7nj_core_080 = popcount28_b7nj_core_078 ^ popcount28_b7nj_core_077;
  assign popcount28_b7nj_core_081 = popcount28_b7nj_core_078 & popcount28_b7nj_core_077;
  assign popcount28_b7nj_core_082 = popcount28_b7nj_core_079 | popcount28_b7nj_core_081;
  assign popcount28_b7nj_core_085 = popcount28_b7nj_core_072 | popcount28_b7nj_core_082;
  assign popcount28_b7nj_core_086 = ~(input_a[0] ^ input_a[13]);
  assign popcount28_b7nj_core_088 = input_a[10] | input_a[8];
  assign popcount28_b7nj_core_089 = ~input_a[12];
  assign popcount28_b7nj_core_091 = ~input_a[18];
  assign popcount28_b7nj_core_094 = input_a[17] ^ input_a[14];
  assign popcount28_b7nj_core_095 = popcount28_b7nj_core_056 ^ popcount28_b7nj_core_085;
  assign popcount28_b7nj_core_096 = popcount28_b7nj_core_056 & popcount28_b7nj_core_085;
  assign popcount28_b7nj_core_098 = ~input_a[3];
  assign popcount28_b7nj_core_102 = popcount28_b7nj_core_057 | popcount28_b7nj_core_096;
  assign popcount28_b7nj_core_103 = input_a[15] & input_a[19];
  assign popcount28_b7nj_core_104 = ~(input_a[6] ^ input_a[3]);
  assign popcount28_b7nj_core_105 = ~(input_a[3] ^ input_a[10]);
  assign popcount28_b7nj_core_106 = ~input_a[26];
  assign popcount28_b7nj_core_107 = ~input_a[10];
  assign popcount28_b7nj_core_108 = input_a[0] & input_a[5];
  assign popcount28_b7nj_core_111 = input_a[17] | input_a[18];
  assign popcount28_b7nj_core_112 = input_a[17] & input_a[18];
  assign popcount28_b7nj_core_113 = ~input_a[23];
  assign popcount28_b7nj_core_114 = input_a[19] & input_a[20];
  assign popcount28_b7nj_core_116 = popcount28_b7nj_core_111 & input_a[25];
  assign popcount28_b7nj_core_117 = popcount28_b7nj_core_112 ^ popcount28_b7nj_core_114;
  assign popcount28_b7nj_core_118 = popcount28_b7nj_core_112 & popcount28_b7nj_core_114;
  assign popcount28_b7nj_core_119 = popcount28_b7nj_core_117 | popcount28_b7nj_core_116;
  assign popcount28_b7nj_core_120 = ~(input_a[4] ^ input_a[21]);
  assign popcount28_b7nj_core_123 = ~(input_a[14] & input_a[2]);
  assign popcount28_b7nj_core_124 = input_a[15] ^ popcount28_b7nj_core_119;
  assign popcount28_b7nj_core_125 = input_a[15] & popcount28_b7nj_core_119;
  assign popcount28_b7nj_core_130 = ~input_a[26];
  assign popcount28_b7nj_core_131 = popcount28_b7nj_core_118 | popcount28_b7nj_core_125;
  assign popcount28_b7nj_core_132 = input_a[25] | input_a[23];
  assign popcount28_b7nj_core_133 = ~input_a[20];
  assign popcount28_b7nj_core_135 = input_a[22] & input_a[23];
  assign popcount28_b7nj_core_137 = input_a[21] & input_a[16];
  assign popcount28_b7nj_core_138 = popcount28_b7nj_core_135 | popcount28_b7nj_core_137;
  assign popcount28_b7nj_core_140 = ~(input_a[19] ^ input_a[1]);
  assign popcount28_b7nj_core_141 = input_a[24] & input_a[0];
  assign popcount28_b7nj_core_142 = input_a[26] ^ input_a[27];
  assign popcount28_b7nj_core_143 = input_a[26] & input_a[27];
  assign popcount28_b7nj_core_144 = ~(input_a[4] & input_a[6]);
  assign popcount28_b7nj_core_145 = input_a[4] & popcount28_b7nj_core_142;
  assign popcount28_b7nj_core_146 = popcount28_b7nj_core_141 ^ popcount28_b7nj_core_143;
  assign popcount28_b7nj_core_147 = popcount28_b7nj_core_141 & popcount28_b7nj_core_143;
  assign popcount28_b7nj_core_148 = popcount28_b7nj_core_146 ^ popcount28_b7nj_core_145;
  assign popcount28_b7nj_core_149 = popcount28_b7nj_core_146 & popcount28_b7nj_core_145;
  assign popcount28_b7nj_core_150 = popcount28_b7nj_core_147 | popcount28_b7nj_core_149;
  assign popcount28_b7nj_core_151 = ~(input_a[11] & input_a[27]);
  assign popcount28_b7nj_core_152 = ~(input_a[7] | input_a[5]);
  assign popcount28_b7nj_core_153 = popcount28_b7nj_core_138 ^ popcount28_b7nj_core_148;
  assign popcount28_b7nj_core_154 = popcount28_b7nj_core_138 & popcount28_b7nj_core_148;
  assign popcount28_b7nj_core_160 = popcount28_b7nj_core_150 | popcount28_b7nj_core_154;
  assign popcount28_b7nj_core_163 = ~input_a[14];
  assign popcount28_b7nj_core_164 = ~(input_a[4] | input_a[12]);
  assign popcount28_b7nj_core_165 = popcount28_b7nj_core_124 ^ popcount28_b7nj_core_153;
  assign popcount28_b7nj_core_166 = popcount28_b7nj_core_124 & popcount28_b7nj_core_153;
  assign popcount28_b7nj_core_167 = popcount28_b7nj_core_165 ^ input_a[14];
  assign popcount28_b7nj_core_168 = popcount28_b7nj_core_165 & input_a[14];
  assign popcount28_b7nj_core_169 = popcount28_b7nj_core_166 | popcount28_b7nj_core_168;
  assign popcount28_b7nj_core_170 = popcount28_b7nj_core_131 ^ popcount28_b7nj_core_160;
  assign popcount28_b7nj_core_171 = popcount28_b7nj_core_131 & popcount28_b7nj_core_160;
  assign popcount28_b7nj_core_172 = popcount28_b7nj_core_170 ^ popcount28_b7nj_core_169;
  assign popcount28_b7nj_core_173 = popcount28_b7nj_core_170 & popcount28_b7nj_core_169;
  assign popcount28_b7nj_core_174 = popcount28_b7nj_core_171 | popcount28_b7nj_core_173;
  assign popcount28_b7nj_core_176 = ~input_a[19];
  assign popcount28_b7nj_core_178 = ~(input_a[9] ^ input_a[27]);
  assign popcount28_b7nj_core_179 = input_a[18] | input_a[8];
  assign popcount28_b7nj_core_180 = input_a[17] ^ input_a[10];
  assign popcount28_b7nj_core_181 = input_a[1] & popcount28_b7nj_core_163;
  assign popcount28_b7nj_core_182 = popcount28_b7nj_core_080 ^ popcount28_b7nj_core_167;
  assign popcount28_b7nj_core_183 = popcount28_b7nj_core_080 & popcount28_b7nj_core_167;
  assign popcount28_b7nj_core_184 = popcount28_b7nj_core_182 ^ popcount28_b7nj_core_181;
  assign popcount28_b7nj_core_185 = popcount28_b7nj_core_182 & popcount28_b7nj_core_181;
  assign popcount28_b7nj_core_186 = popcount28_b7nj_core_183 | popcount28_b7nj_core_185;
  assign popcount28_b7nj_core_187 = popcount28_b7nj_core_095 ^ popcount28_b7nj_core_172;
  assign popcount28_b7nj_core_188 = popcount28_b7nj_core_095 & popcount28_b7nj_core_172;
  assign popcount28_b7nj_core_189 = popcount28_b7nj_core_187 ^ popcount28_b7nj_core_186;
  assign popcount28_b7nj_core_190 = popcount28_b7nj_core_187 & popcount28_b7nj_core_186;
  assign popcount28_b7nj_core_191 = popcount28_b7nj_core_188 | popcount28_b7nj_core_190;
  assign popcount28_b7nj_core_192 = popcount28_b7nj_core_102 ^ popcount28_b7nj_core_174;
  assign popcount28_b7nj_core_193 = popcount28_b7nj_core_102 & popcount28_b7nj_core_174;
  assign popcount28_b7nj_core_194 = popcount28_b7nj_core_192 ^ popcount28_b7nj_core_191;
  assign popcount28_b7nj_core_195 = popcount28_b7nj_core_192 & popcount28_b7nj_core_191;
  assign popcount28_b7nj_core_196 = popcount28_b7nj_core_193 | popcount28_b7nj_core_195;
  assign popcount28_b7nj_core_197 = input_a[2] ^ input_a[8];
  assign popcount28_b7nj_core_198 = input_a[4] & input_a[22];
  assign popcount28_b7nj_core_199 = input_a[18] | input_a[9];
  assign popcount28_b7nj_core_200 = ~(input_a[10] | input_a[6]);

  assign popcount28_b7nj_out[0] = 1'b0;
  assign popcount28_b7nj_out[1] = popcount28_b7nj_core_184;
  assign popcount28_b7nj_out[2] = popcount28_b7nj_core_189;
  assign popcount28_b7nj_out[3] = popcount28_b7nj_core_194;
  assign popcount28_b7nj_out[4] = popcount28_b7nj_core_196;
endmodule