// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.89482
// WCE=16.0
// EP=0.92946%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount19_zvgu(input [18:0] input_a, output [4:0] popcount19_zvgu_out);
  wire popcount19_zvgu_core_021;
  wire popcount19_zvgu_core_023;
  wire popcount19_zvgu_core_024;
  wire popcount19_zvgu_core_025;
  wire popcount19_zvgu_core_026;
  wire popcount19_zvgu_core_027;
  wire popcount19_zvgu_core_029;
  wire popcount19_zvgu_core_032;
  wire popcount19_zvgu_core_034;
  wire popcount19_zvgu_core_036;
  wire popcount19_zvgu_core_037;
  wire popcount19_zvgu_core_039;
  wire popcount19_zvgu_core_041;
  wire popcount19_zvgu_core_042;
  wire popcount19_zvgu_core_045;
  wire popcount19_zvgu_core_049;
  wire popcount19_zvgu_core_052;
  wire popcount19_zvgu_core_054;
  wire popcount19_zvgu_core_056;
  wire popcount19_zvgu_core_058;
  wire popcount19_zvgu_core_059_not;
  wire popcount19_zvgu_core_061;
  wire popcount19_zvgu_core_063;
  wire popcount19_zvgu_core_064;
  wire popcount19_zvgu_core_065;
  wire popcount19_zvgu_core_066;
  wire popcount19_zvgu_core_068;
  wire popcount19_zvgu_core_069;
  wire popcount19_zvgu_core_071;
  wire popcount19_zvgu_core_072;
  wire popcount19_zvgu_core_075;
  wire popcount19_zvgu_core_076;
  wire popcount19_zvgu_core_077;
  wire popcount19_zvgu_core_078;
  wire popcount19_zvgu_core_080;
  wire popcount19_zvgu_core_082;
  wire popcount19_zvgu_core_083;
  wire popcount19_zvgu_core_084;
  wire popcount19_zvgu_core_085;
  wire popcount19_zvgu_core_087;
  wire popcount19_zvgu_core_088_not;
  wire popcount19_zvgu_core_089;
  wire popcount19_zvgu_core_091;
  wire popcount19_zvgu_core_092;
  wire popcount19_zvgu_core_094_not;
  wire popcount19_zvgu_core_096;
  wire popcount19_zvgu_core_097;
  wire popcount19_zvgu_core_098;
  wire popcount19_zvgu_core_099;
  wire popcount19_zvgu_core_100;
  wire popcount19_zvgu_core_102;
  wire popcount19_zvgu_core_103;
  wire popcount19_zvgu_core_104;
  wire popcount19_zvgu_core_105;
  wire popcount19_zvgu_core_106;
  wire popcount19_zvgu_core_107;
  wire popcount19_zvgu_core_108;
  wire popcount19_zvgu_core_109;
  wire popcount19_zvgu_core_110_not;
  wire popcount19_zvgu_core_111;
  wire popcount19_zvgu_core_114;
  wire popcount19_zvgu_core_116;
  wire popcount19_zvgu_core_117;
  wire popcount19_zvgu_core_122;
  wire popcount19_zvgu_core_123;
  wire popcount19_zvgu_core_124;
  wire popcount19_zvgu_core_126;
  wire popcount19_zvgu_core_128;
  wire popcount19_zvgu_core_129;
  wire popcount19_zvgu_core_130;
  wire popcount19_zvgu_core_131_not;
  wire popcount19_zvgu_core_132;
  wire popcount19_zvgu_core_133;
  wire popcount19_zvgu_core_135;

  assign popcount19_zvgu_core_021 = ~(input_a[18] | input_a[2]);
  assign popcount19_zvgu_core_023 = input_a[1] ^ input_a[7];
  assign popcount19_zvgu_core_024 = ~(input_a[11] & input_a[14]);
  assign popcount19_zvgu_core_025 = ~(input_a[10] ^ input_a[15]);
  assign popcount19_zvgu_core_026 = ~(input_a[4] & input_a[5]);
  assign popcount19_zvgu_core_027 = ~input_a[2];
  assign popcount19_zvgu_core_029 = input_a[14] ^ input_a[6];
  assign popcount19_zvgu_core_032 = ~(input_a[6] | input_a[18]);
  assign popcount19_zvgu_core_034 = ~(input_a[0] ^ input_a[11]);
  assign popcount19_zvgu_core_036 = input_a[7] | input_a[17];
  assign popcount19_zvgu_core_037 = ~(input_a[17] | input_a[17]);
  assign popcount19_zvgu_core_039 = ~(input_a[10] | input_a[4]);
  assign popcount19_zvgu_core_041 = input_a[12] ^ input_a[0];
  assign popcount19_zvgu_core_042 = ~input_a[12];
  assign popcount19_zvgu_core_045 = input_a[10] ^ input_a[15];
  assign popcount19_zvgu_core_049 = ~(input_a[11] ^ input_a[4]);
  assign popcount19_zvgu_core_052 = ~(input_a[16] ^ input_a[4]);
  assign popcount19_zvgu_core_054 = ~(input_a[1] & input_a[9]);
  assign popcount19_zvgu_core_056 = ~(input_a[1] & input_a[16]);
  assign popcount19_zvgu_core_058 = input_a[0] & input_a[6];
  assign popcount19_zvgu_core_059_not = ~input_a[13];
  assign popcount19_zvgu_core_061 = ~(input_a[12] | input_a[13]);
  assign popcount19_zvgu_core_063 = ~input_a[12];
  assign popcount19_zvgu_core_064 = input_a[0] ^ input_a[1];
  assign popcount19_zvgu_core_065 = ~(input_a[18] & input_a[10]);
  assign popcount19_zvgu_core_066 = ~(input_a[17] ^ input_a[0]);
  assign popcount19_zvgu_core_068 = ~input_a[17];
  assign popcount19_zvgu_core_069 = ~input_a[9];
  assign popcount19_zvgu_core_071 = ~(input_a[12] | input_a[4]);
  assign popcount19_zvgu_core_072 = input_a[14] & input_a[15];
  assign popcount19_zvgu_core_075 = ~(input_a[13] & input_a[13]);
  assign popcount19_zvgu_core_076 = ~input_a[8];
  assign popcount19_zvgu_core_077 = ~input_a[5];
  assign popcount19_zvgu_core_078 = ~input_a[6];
  assign popcount19_zvgu_core_080 = ~(input_a[12] & input_a[16]);
  assign popcount19_zvgu_core_082 = input_a[5] ^ input_a[11];
  assign popcount19_zvgu_core_083 = ~input_a[4];
  assign popcount19_zvgu_core_084 = ~input_a[18];
  assign popcount19_zvgu_core_085 = ~(input_a[8] ^ input_a[2]);
  assign popcount19_zvgu_core_087 = input_a[3] ^ input_a[17];
  assign popcount19_zvgu_core_088_not = ~input_a[15];
  assign popcount19_zvgu_core_089 = ~(input_a[2] | input_a[11]);
  assign popcount19_zvgu_core_091 = ~(input_a[16] ^ input_a[14]);
  assign popcount19_zvgu_core_092 = ~(input_a[15] | input_a[16]);
  assign popcount19_zvgu_core_094_not = ~input_a[18];
  assign popcount19_zvgu_core_096 = input_a[13] ^ input_a[0];
  assign popcount19_zvgu_core_097 = input_a[0] & input_a[18];
  assign popcount19_zvgu_core_098 = ~input_a[16];
  assign popcount19_zvgu_core_099 = input_a[6] & input_a[10];
  assign popcount19_zvgu_core_100 = ~(input_a[9] | input_a[14]);
  assign popcount19_zvgu_core_102 = input_a[0] & input_a[17];
  assign popcount19_zvgu_core_103 = ~input_a[7];
  assign popcount19_zvgu_core_104 = input_a[8] & input_a[5];
  assign popcount19_zvgu_core_105 = input_a[8] | input_a[10];
  assign popcount19_zvgu_core_106 = input_a[18] | input_a[14];
  assign popcount19_zvgu_core_107 = ~input_a[17];
  assign popcount19_zvgu_core_108 = input_a[12] | input_a[7];
  assign popcount19_zvgu_core_109 = input_a[12] & input_a[6];
  assign popcount19_zvgu_core_110_not = ~input_a[13];
  assign popcount19_zvgu_core_111 = ~(input_a[2] & input_a[5]);
  assign popcount19_zvgu_core_114 = ~(input_a[17] | input_a[18]);
  assign popcount19_zvgu_core_116 = input_a[15] & input_a[7];
  assign popcount19_zvgu_core_117 = ~input_a[7];
  assign popcount19_zvgu_core_122 = input_a[17] & input_a[8];
  assign popcount19_zvgu_core_123 = input_a[1] & input_a[3];
  assign popcount19_zvgu_core_124 = ~input_a[15];
  assign popcount19_zvgu_core_126 = ~input_a[11];
  assign popcount19_zvgu_core_128 = input_a[4] ^ input_a[7];
  assign popcount19_zvgu_core_129 = ~input_a[18];
  assign popcount19_zvgu_core_130 = ~(input_a[13] & input_a[0]);
  assign popcount19_zvgu_core_131_not = ~input_a[4];
  assign popcount19_zvgu_core_132 = input_a[3] ^ input_a[9];
  assign popcount19_zvgu_core_133 = ~(input_a[13] & input_a[18]);
  assign popcount19_zvgu_core_135 = ~(input_a[12] & input_a[4]);

  assign popcount19_zvgu_out[0] = 1'b1;
  assign popcount19_zvgu_out[1] = 1'b1;
  assign popcount19_zvgu_out[2] = input_a[2];
  assign popcount19_zvgu_out[3] = input_a[4];
  assign popcount19_zvgu_out[4] = 1'b0;
endmodule