// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.75816
// WCE=21.0
// EP=0.886569%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount40_w51f(input [39:0] input_a, output [5:0] popcount40_w51f_out);
  wire popcount40_w51f_core_043;
  wire popcount40_w51f_core_044;
  wire popcount40_w51f_core_045_not;
  wire popcount40_w51f_core_046;
  wire popcount40_w51f_core_047;
  wire popcount40_w51f_core_048;
  wire popcount40_w51f_core_049;
  wire popcount40_w51f_core_050;
  wire popcount40_w51f_core_051;
  wire popcount40_w51f_core_053;
  wire popcount40_w51f_core_055;
  wire popcount40_w51f_core_056;
  wire popcount40_w51f_core_058;
  wire popcount40_w51f_core_059;
  wire popcount40_w51f_core_060_not;
  wire popcount40_w51f_core_061;
  wire popcount40_w51f_core_062;
  wire popcount40_w51f_core_063;
  wire popcount40_w51f_core_064;
  wire popcount40_w51f_core_068;
  wire popcount40_w51f_core_069;
  wire popcount40_w51f_core_072;
  wire popcount40_w51f_core_074;
  wire popcount40_w51f_core_075;
  wire popcount40_w51f_core_076;
  wire popcount40_w51f_core_077;
  wire popcount40_w51f_core_078;
  wire popcount40_w51f_core_079;
  wire popcount40_w51f_core_080;
  wire popcount40_w51f_core_081;
  wire popcount40_w51f_core_082;
  wire popcount40_w51f_core_083_not;
  wire popcount40_w51f_core_084;
  wire popcount40_w51f_core_085;
  wire popcount40_w51f_core_087;
  wire popcount40_w51f_core_088;
  wire popcount40_w51f_core_090;
  wire popcount40_w51f_core_091;
  wire popcount40_w51f_core_093;
  wire popcount40_w51f_core_094_not;
  wire popcount40_w51f_core_095;
  wire popcount40_w51f_core_096;
  wire popcount40_w51f_core_097;
  wire popcount40_w51f_core_098;
  wire popcount40_w51f_core_100;
  wire popcount40_w51f_core_101;
  wire popcount40_w51f_core_102;
  wire popcount40_w51f_core_103;
  wire popcount40_w51f_core_104;
  wire popcount40_w51f_core_105;
  wire popcount40_w51f_core_106;
  wire popcount40_w51f_core_108;
  wire popcount40_w51f_core_111;
  wire popcount40_w51f_core_112;
  wire popcount40_w51f_core_113;
  wire popcount40_w51f_core_116;
  wire popcount40_w51f_core_117;
  wire popcount40_w51f_core_119;
  wire popcount40_w51f_core_120;
  wire popcount40_w51f_core_123;
  wire popcount40_w51f_core_124;
  wire popcount40_w51f_core_125;
  wire popcount40_w51f_core_126;
  wire popcount40_w51f_core_127;
  wire popcount40_w51f_core_128;
  wire popcount40_w51f_core_129;
  wire popcount40_w51f_core_131;
  wire popcount40_w51f_core_132;
  wire popcount40_w51f_core_135;
  wire popcount40_w51f_core_136;
  wire popcount40_w51f_core_138;
  wire popcount40_w51f_core_139;
  wire popcount40_w51f_core_140;
  wire popcount40_w51f_core_142;
  wire popcount40_w51f_core_143;
  wire popcount40_w51f_core_144;
  wire popcount40_w51f_core_145_not;
  wire popcount40_w51f_core_146;
  wire popcount40_w51f_core_147;
  wire popcount40_w51f_core_148;
  wire popcount40_w51f_core_150;
  wire popcount40_w51f_core_153;
  wire popcount40_w51f_core_154;
  wire popcount40_w51f_core_155;
  wire popcount40_w51f_core_156;
  wire popcount40_w51f_core_158;
  wire popcount40_w51f_core_159;
  wire popcount40_w51f_core_160;
  wire popcount40_w51f_core_161;
  wire popcount40_w51f_core_163;
  wire popcount40_w51f_core_164;
  wire popcount40_w51f_core_165;
  wire popcount40_w51f_core_166;
  wire popcount40_w51f_core_169;
  wire popcount40_w51f_core_170;
  wire popcount40_w51f_core_172;
  wire popcount40_w51f_core_175;
  wire popcount40_w51f_core_177;
  wire popcount40_w51f_core_179;
  wire popcount40_w51f_core_181;
  wire popcount40_w51f_core_182;
  wire popcount40_w51f_core_183;
  wire popcount40_w51f_core_185;
  wire popcount40_w51f_core_187;
  wire popcount40_w51f_core_188;
  wire popcount40_w51f_core_189;
  wire popcount40_w51f_core_190;
  wire popcount40_w51f_core_192;
  wire popcount40_w51f_core_194;
  wire popcount40_w51f_core_195;
  wire popcount40_w51f_core_196;
  wire popcount40_w51f_core_198;
  wire popcount40_w51f_core_199;
  wire popcount40_w51f_core_200;
  wire popcount40_w51f_core_201;
  wire popcount40_w51f_core_202;
  wire popcount40_w51f_core_205;
  wire popcount40_w51f_core_206;
  wire popcount40_w51f_core_207_not;
  wire popcount40_w51f_core_208;
  wire popcount40_w51f_core_209;
  wire popcount40_w51f_core_210;
  wire popcount40_w51f_core_211;
  wire popcount40_w51f_core_214;
  wire popcount40_w51f_core_215;
  wire popcount40_w51f_core_216;
  wire popcount40_w51f_core_217;
  wire popcount40_w51f_core_218;
  wire popcount40_w51f_core_219;
  wire popcount40_w51f_core_220;
  wire popcount40_w51f_core_223;
  wire popcount40_w51f_core_227;
  wire popcount40_w51f_core_228;
  wire popcount40_w51f_core_230;
  wire popcount40_w51f_core_231;
  wire popcount40_w51f_core_232;
  wire popcount40_w51f_core_233;
  wire popcount40_w51f_core_234;
  wire popcount40_w51f_core_235;
  wire popcount40_w51f_core_236;
  wire popcount40_w51f_core_238;
  wire popcount40_w51f_core_241;
  wire popcount40_w51f_core_242;
  wire popcount40_w51f_core_243;
  wire popcount40_w51f_core_246;
  wire popcount40_w51f_core_247;
  wire popcount40_w51f_core_249;
  wire popcount40_w51f_core_250;
  wire popcount40_w51f_core_251;
  wire popcount40_w51f_core_252;
  wire popcount40_w51f_core_255;
  wire popcount40_w51f_core_256;
  wire popcount40_w51f_core_257;
  wire popcount40_w51f_core_258;
  wire popcount40_w51f_core_261;
  wire popcount40_w51f_core_262_not;
  wire popcount40_w51f_core_263;
  wire popcount40_w51f_core_265;
  wire popcount40_w51f_core_266;
  wire popcount40_w51f_core_267;
  wire popcount40_w51f_core_268;
  wire popcount40_w51f_core_269;
  wire popcount40_w51f_core_274;
  wire popcount40_w51f_core_275;
  wire popcount40_w51f_core_276;
  wire popcount40_w51f_core_277_not;
  wire popcount40_w51f_core_279;
  wire popcount40_w51f_core_282;
  wire popcount40_w51f_core_284;
  wire popcount40_w51f_core_286;
  wire popcount40_w51f_core_289;
  wire popcount40_w51f_core_290;
  wire popcount40_w51f_core_291;
  wire popcount40_w51f_core_292;
  wire popcount40_w51f_core_294;
  wire popcount40_w51f_core_295;
  wire popcount40_w51f_core_296;
  wire popcount40_w51f_core_297;
  wire popcount40_w51f_core_298;
  wire popcount40_w51f_core_299;
  wire popcount40_w51f_core_300;
  wire popcount40_w51f_core_303;
  wire popcount40_w51f_core_304;
  wire popcount40_w51f_core_306;
  wire popcount40_w51f_core_308;
  wire popcount40_w51f_core_309;
  wire popcount40_w51f_core_310;
  wire popcount40_w51f_core_313;
  wire popcount40_w51f_core_314;
  wire popcount40_w51f_core_315;
  wire popcount40_w51f_core_316;

  assign popcount40_w51f_core_043 = input_a[13] & input_a[23];
  assign popcount40_w51f_core_044 = ~input_a[34];
  assign popcount40_w51f_core_045_not = ~input_a[31];
  assign popcount40_w51f_core_046 = ~(input_a[18] & input_a[4]);
  assign popcount40_w51f_core_047 = input_a[38] | input_a[23];
  assign popcount40_w51f_core_048 = ~(input_a[14] & input_a[23]);
  assign popcount40_w51f_core_049 = ~(input_a[29] ^ input_a[8]);
  assign popcount40_w51f_core_050 = input_a[8] | input_a[12];
  assign popcount40_w51f_core_051 = input_a[14] & input_a[14];
  assign popcount40_w51f_core_053 = ~(input_a[31] | input_a[29]);
  assign popcount40_w51f_core_055 = ~input_a[12];
  assign popcount40_w51f_core_056 = input_a[8] & input_a[30];
  assign popcount40_w51f_core_058 = ~input_a[12];
  assign popcount40_w51f_core_059 = ~(input_a[6] ^ input_a[8]);
  assign popcount40_w51f_core_060_not = ~input_a[7];
  assign popcount40_w51f_core_061 = ~input_a[19];
  assign popcount40_w51f_core_062 = ~input_a[13];
  assign popcount40_w51f_core_063 = ~(input_a[10] ^ input_a[19]);
  assign popcount40_w51f_core_064 = input_a[29] | input_a[35];
  assign popcount40_w51f_core_068 = input_a[33] | input_a[31];
  assign popcount40_w51f_core_069 = ~(input_a[15] | input_a[31]);
  assign popcount40_w51f_core_072 = input_a[11] & input_a[19];
  assign popcount40_w51f_core_074 = input_a[21] | input_a[3];
  assign popcount40_w51f_core_075 = input_a[23] | input_a[7];
  assign popcount40_w51f_core_076 = ~(input_a[35] & input_a[33]);
  assign popcount40_w51f_core_077 = ~input_a[26];
  assign popcount40_w51f_core_078 = input_a[9] & input_a[17];
  assign popcount40_w51f_core_079 = input_a[35] & input_a[16];
  assign popcount40_w51f_core_080 = ~(input_a[26] & input_a[32]);
  assign popcount40_w51f_core_081 = input_a[9] ^ input_a[10];
  assign popcount40_w51f_core_082 = ~(input_a[13] & input_a[8]);
  assign popcount40_w51f_core_083_not = ~input_a[25];
  assign popcount40_w51f_core_084 = input_a[13] ^ input_a[24];
  assign popcount40_w51f_core_085 = ~input_a[17];
  assign popcount40_w51f_core_087 = ~(input_a[10] | input_a[34]);
  assign popcount40_w51f_core_088 = ~(input_a[0] & input_a[28]);
  assign popcount40_w51f_core_090 = input_a[3] | input_a[18];
  assign popcount40_w51f_core_091 = input_a[0] & input_a[14];
  assign popcount40_w51f_core_093 = ~(input_a[12] | input_a[4]);
  assign popcount40_w51f_core_094_not = ~input_a[37];
  assign popcount40_w51f_core_095 = input_a[17] ^ input_a[26];
  assign popcount40_w51f_core_096 = ~(input_a[24] | input_a[17]);
  assign popcount40_w51f_core_097 = input_a[9] ^ input_a[10];
  assign popcount40_w51f_core_098 = ~(input_a[38] | input_a[32]);
  assign popcount40_w51f_core_100 = input_a[33] ^ input_a[28];
  assign popcount40_w51f_core_101 = input_a[15] & input_a[38];
  assign popcount40_w51f_core_102 = ~(input_a[22] & input_a[5]);
  assign popcount40_w51f_core_103 = input_a[7] | input_a[18];
  assign popcount40_w51f_core_104 = ~(input_a[14] | input_a[31]);
  assign popcount40_w51f_core_105 = ~input_a[8];
  assign popcount40_w51f_core_106 = ~(input_a[19] ^ input_a[12]);
  assign popcount40_w51f_core_108 = input_a[39] ^ input_a[20];
  assign popcount40_w51f_core_111 = input_a[30] & input_a[5];
  assign popcount40_w51f_core_112 = input_a[8] | input_a[33];
  assign popcount40_w51f_core_113 = ~(input_a[23] ^ input_a[5]);
  assign popcount40_w51f_core_116 = ~input_a[38];
  assign popcount40_w51f_core_117 = ~(input_a[11] | input_a[24]);
  assign popcount40_w51f_core_119 = ~(input_a[12] ^ input_a[10]);
  assign popcount40_w51f_core_120 = ~(input_a[15] | input_a[7]);
  assign popcount40_w51f_core_123 = ~(input_a[30] | input_a[5]);
  assign popcount40_w51f_core_124 = ~(input_a[34] ^ input_a[26]);
  assign popcount40_w51f_core_125 = ~(input_a[29] | input_a[1]);
  assign popcount40_w51f_core_126 = input_a[22] | input_a[29];
  assign popcount40_w51f_core_127 = input_a[9] ^ input_a[13];
  assign popcount40_w51f_core_128 = ~input_a[18];
  assign popcount40_w51f_core_129 = ~(input_a[33] ^ input_a[26]);
  assign popcount40_w51f_core_131 = ~(input_a[20] | input_a[21]);
  assign popcount40_w51f_core_132 = ~(input_a[18] ^ input_a[29]);
  assign popcount40_w51f_core_135 = ~(input_a[26] ^ input_a[27]);
  assign popcount40_w51f_core_136 = ~(input_a[22] ^ input_a[17]);
  assign popcount40_w51f_core_138 = ~input_a[7];
  assign popcount40_w51f_core_139 = input_a[3] & input_a[39];
  assign popcount40_w51f_core_140 = ~(input_a[23] ^ input_a[17]);
  assign popcount40_w51f_core_142 = ~(input_a[28] | input_a[14]);
  assign popcount40_w51f_core_143 = ~(input_a[1] | input_a[7]);
  assign popcount40_w51f_core_144 = input_a[5] | input_a[39];
  assign popcount40_w51f_core_145_not = ~input_a[30];
  assign popcount40_w51f_core_146 = ~(input_a[9] | input_a[28]);
  assign popcount40_w51f_core_147 = ~(input_a[0] ^ input_a[4]);
  assign popcount40_w51f_core_148 = ~(input_a[28] & input_a[14]);
  assign popcount40_w51f_core_150 = ~input_a[10];
  assign popcount40_w51f_core_153 = ~(input_a[6] & input_a[13]);
  assign popcount40_w51f_core_154 = ~(input_a[36] | input_a[22]);
  assign popcount40_w51f_core_155 = ~(input_a[29] ^ input_a[5]);
  assign popcount40_w51f_core_156 = input_a[24] ^ input_a[3];
  assign popcount40_w51f_core_158 = input_a[6] ^ input_a[1];
  assign popcount40_w51f_core_159 = ~(input_a[35] | input_a[24]);
  assign popcount40_w51f_core_160 = ~input_a[23];
  assign popcount40_w51f_core_161 = ~input_a[22];
  assign popcount40_w51f_core_163 = input_a[8] & input_a[3];
  assign popcount40_w51f_core_164 = ~input_a[25];
  assign popcount40_w51f_core_165 = input_a[18] ^ input_a[23];
  assign popcount40_w51f_core_166 = input_a[13] & input_a[33];
  assign popcount40_w51f_core_169 = input_a[18] & input_a[20];
  assign popcount40_w51f_core_170 = input_a[20] & input_a[4];
  assign popcount40_w51f_core_172 = ~(input_a[21] | input_a[17]);
  assign popcount40_w51f_core_175 = input_a[14] ^ input_a[38];
  assign popcount40_w51f_core_177 = ~(input_a[31] | input_a[24]);
  assign popcount40_w51f_core_179 = input_a[25] & input_a[24];
  assign popcount40_w51f_core_181 = ~(input_a[1] ^ input_a[1]);
  assign popcount40_w51f_core_182 = ~(input_a[7] | input_a[11]);
  assign popcount40_w51f_core_183 = ~(input_a[2] & input_a[0]);
  assign popcount40_w51f_core_185 = input_a[11] & input_a[29];
  assign popcount40_w51f_core_187 = input_a[37] ^ input_a[22];
  assign popcount40_w51f_core_188 = ~(input_a[19] ^ input_a[16]);
  assign popcount40_w51f_core_189 = ~input_a[8];
  assign popcount40_w51f_core_190 = input_a[29] & input_a[5];
  assign popcount40_w51f_core_192 = input_a[2] & input_a[6];
  assign popcount40_w51f_core_194 = input_a[8] | input_a[33];
  assign popcount40_w51f_core_195 = ~(input_a[30] & input_a[15]);
  assign popcount40_w51f_core_196 = input_a[39] | input_a[23];
  assign popcount40_w51f_core_198 = input_a[34] & input_a[25];
  assign popcount40_w51f_core_199 = ~(input_a[18] | input_a[11]);
  assign popcount40_w51f_core_200 = ~input_a[14];
  assign popcount40_w51f_core_201 = input_a[28] ^ input_a[23];
  assign popcount40_w51f_core_202 = ~(input_a[18] | input_a[29]);
  assign popcount40_w51f_core_205 = ~(input_a[38] & input_a[30]);
  assign popcount40_w51f_core_206 = ~(input_a[25] ^ input_a[37]);
  assign popcount40_w51f_core_207_not = ~input_a[11];
  assign popcount40_w51f_core_208 = input_a[18] & input_a[5];
  assign popcount40_w51f_core_209 = input_a[29] ^ input_a[16];
  assign popcount40_w51f_core_210 = ~(input_a[32] ^ input_a[15]);
  assign popcount40_w51f_core_211 = ~input_a[39];
  assign popcount40_w51f_core_214 = ~(input_a[19] | input_a[7]);
  assign popcount40_w51f_core_215 = input_a[15] & input_a[33];
  assign popcount40_w51f_core_216 = input_a[23] | input_a[28];
  assign popcount40_w51f_core_217 = input_a[22] ^ input_a[11];
  assign popcount40_w51f_core_218 = ~(input_a[11] & input_a[28]);
  assign popcount40_w51f_core_219 = input_a[38] ^ input_a[4];
  assign popcount40_w51f_core_220 = ~(input_a[1] | input_a[7]);
  assign popcount40_w51f_core_223 = ~(input_a[30] ^ input_a[30]);
  assign popcount40_w51f_core_227 = input_a[36] | input_a[26];
  assign popcount40_w51f_core_228 = ~(input_a[20] & input_a[10]);
  assign popcount40_w51f_core_230 = ~input_a[12];
  assign popcount40_w51f_core_231 = ~(input_a[29] & input_a[38]);
  assign popcount40_w51f_core_232 = ~(input_a[33] | input_a[10]);
  assign popcount40_w51f_core_233 = input_a[36] | input_a[6];
  assign popcount40_w51f_core_234 = input_a[18] | input_a[27];
  assign popcount40_w51f_core_235 = ~input_a[9];
  assign popcount40_w51f_core_236 = input_a[9] ^ input_a[8];
  assign popcount40_w51f_core_238 = input_a[8] ^ input_a[26];
  assign popcount40_w51f_core_241 = ~(input_a[15] | input_a[14]);
  assign popcount40_w51f_core_242 = ~(input_a[9] ^ input_a[8]);
  assign popcount40_w51f_core_243 = input_a[6] & input_a[36];
  assign popcount40_w51f_core_246 = ~(input_a[3] ^ input_a[10]);
  assign popcount40_w51f_core_247 = ~input_a[9];
  assign popcount40_w51f_core_249 = input_a[5] & input_a[5];
  assign popcount40_w51f_core_250 = input_a[17] & input_a[4];
  assign popcount40_w51f_core_251 = input_a[24] ^ input_a[0];
  assign popcount40_w51f_core_252 = input_a[13] | input_a[19];
  assign popcount40_w51f_core_255 = ~(input_a[29] | input_a[39]);
  assign popcount40_w51f_core_256 = input_a[29] & input_a[12];
  assign popcount40_w51f_core_257 = ~input_a[38];
  assign popcount40_w51f_core_258 = input_a[30] ^ input_a[3];
  assign popcount40_w51f_core_261 = input_a[39] | input_a[10];
  assign popcount40_w51f_core_262_not = ~input_a[38];
  assign popcount40_w51f_core_263 = input_a[22] & input_a[4];
  assign popcount40_w51f_core_265 = input_a[7] ^ input_a[14];
  assign popcount40_w51f_core_266 = ~(input_a[27] | input_a[38]);
  assign popcount40_w51f_core_267 = ~(input_a[30] & input_a[22]);
  assign popcount40_w51f_core_268 = ~(input_a[13] ^ input_a[2]);
  assign popcount40_w51f_core_269 = ~input_a[11];
  assign popcount40_w51f_core_274 = ~(input_a[4] ^ input_a[36]);
  assign popcount40_w51f_core_275 = ~(input_a[21] | input_a[10]);
  assign popcount40_w51f_core_276 = ~input_a[10];
  assign popcount40_w51f_core_277_not = ~input_a[8];
  assign popcount40_w51f_core_279 = input_a[31] & input_a[32];
  assign popcount40_w51f_core_282 = ~input_a[29];
  assign popcount40_w51f_core_284 = input_a[3] ^ input_a[28];
  assign popcount40_w51f_core_286 = ~input_a[32];
  assign popcount40_w51f_core_289 = ~(input_a[11] | input_a[36]);
  assign popcount40_w51f_core_290 = input_a[13] | input_a[3];
  assign popcount40_w51f_core_291 = input_a[7] | input_a[17];
  assign popcount40_w51f_core_292 = ~(input_a[19] | input_a[2]);
  assign popcount40_w51f_core_294 = ~input_a[39];
  assign popcount40_w51f_core_295 = input_a[17] | input_a[2];
  assign popcount40_w51f_core_296 = input_a[19] | input_a[23];
  assign popcount40_w51f_core_297 = ~(input_a[8] ^ input_a[36]);
  assign popcount40_w51f_core_298 = ~(input_a[23] & input_a[19]);
  assign popcount40_w51f_core_299 = input_a[39] ^ input_a[11];
  assign popcount40_w51f_core_300 = input_a[26] ^ input_a[9];
  assign popcount40_w51f_core_303 = ~input_a[18];
  assign popcount40_w51f_core_304 = input_a[28] & input_a[7];
  assign popcount40_w51f_core_306 = ~(input_a[4] ^ input_a[8]);
  assign popcount40_w51f_core_308 = ~(input_a[9] | input_a[12]);
  assign popcount40_w51f_core_309 = ~(input_a[9] ^ input_a[20]);
  assign popcount40_w51f_core_310 = ~(input_a[32] & input_a[9]);
  assign popcount40_w51f_core_313 = input_a[25] | input_a[7];
  assign popcount40_w51f_core_314 = input_a[9] | input_a[26];
  assign popcount40_w51f_core_315 = ~(input_a[9] | input_a[20]);
  assign popcount40_w51f_core_316 = ~(input_a[6] ^ input_a[37]);

  assign popcount40_w51f_out[0] = input_a[14];
  assign popcount40_w51f_out[1] = input_a[16];
  assign popcount40_w51f_out[2] = input_a[17];
  assign popcount40_w51f_out[3] = 1'b0;
  assign popcount40_w51f_out[4] = 1'b1;
  assign popcount40_w51f_out[5] = 1'b0;
endmodule