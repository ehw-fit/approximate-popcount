// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.85317
// WCE=17.0
// EP=0.894307%
// Printed PDK parameters:
//  Area=627920.0
//  Delay=2618200.0
//  Power=30372.0

module popcount31_qr3w(input [30:0] input_a, output [4:0] popcount31_qr3w_out);
  wire popcount31_qr3w_core_033;
  wire popcount31_qr3w_core_034;
  wire popcount31_qr3w_core_035;
  wire popcount31_qr3w_core_037;
  wire popcount31_qr3w_core_039;
  wire popcount31_qr3w_core_040;
  wire popcount31_qr3w_core_042;
  wire popcount31_qr3w_core_043;
  wire popcount31_qr3w_core_044;
  wire popcount31_qr3w_core_045;
  wire popcount31_qr3w_core_046;
  wire popcount31_qr3w_core_048;
  wire popcount31_qr3w_core_049;
  wire popcount31_qr3w_core_050;
  wire popcount31_qr3w_core_051;
  wire popcount31_qr3w_core_052;
  wire popcount31_qr3w_core_053;
  wire popcount31_qr3w_core_054;
  wire popcount31_qr3w_core_058;
  wire popcount31_qr3w_core_059;
  wire popcount31_qr3w_core_060;
  wire popcount31_qr3w_core_062;
  wire popcount31_qr3w_core_064;
  wire popcount31_qr3w_core_066;
  wire popcount31_qr3w_core_069;
  wire popcount31_qr3w_core_073;
  wire popcount31_qr3w_core_075;
  wire popcount31_qr3w_core_076;
  wire popcount31_qr3w_core_078;
  wire popcount31_qr3w_core_079;
  wire popcount31_qr3w_core_081;
  wire popcount31_qr3w_core_082;
  wire popcount31_qr3w_core_086;
  wire popcount31_qr3w_core_088;
  wire popcount31_qr3w_core_091;
  wire popcount31_qr3w_core_093;
  wire popcount31_qr3w_core_096;
  wire popcount31_qr3w_core_098;
  wire popcount31_qr3w_core_099;
  wire popcount31_qr3w_core_100;
  wire popcount31_qr3w_core_101;
  wire popcount31_qr3w_core_102;
  wire popcount31_qr3w_core_103;
  wire popcount31_qr3w_core_104;
  wire popcount31_qr3w_core_105;
  wire popcount31_qr3w_core_106;
  wire popcount31_qr3w_core_107;
  wire popcount31_qr3w_core_108;
  wire popcount31_qr3w_core_111;
  wire popcount31_qr3w_core_113;
  wire popcount31_qr3w_core_114;
  wire popcount31_qr3w_core_115;
  wire popcount31_qr3w_core_116;
  wire popcount31_qr3w_core_119;
  wire popcount31_qr3w_core_120;
  wire popcount31_qr3w_core_122;
  wire popcount31_qr3w_core_125;
  wire popcount31_qr3w_core_126;
  wire popcount31_qr3w_core_128;
  wire popcount31_qr3w_core_129;
  wire popcount31_qr3w_core_130;
  wire popcount31_qr3w_core_131;
  wire popcount31_qr3w_core_132;
  wire popcount31_qr3w_core_134;
  wire popcount31_qr3w_core_135;
  wire popcount31_qr3w_core_136;
  wire popcount31_qr3w_core_137;
  wire popcount31_qr3w_core_140;
  wire popcount31_qr3w_core_141;
  wire popcount31_qr3w_core_143;
  wire popcount31_qr3w_core_152;
  wire popcount31_qr3w_core_154_not;
  wire popcount31_qr3w_core_156;
  wire popcount31_qr3w_core_158;
  wire popcount31_qr3w_core_160;
  wire popcount31_qr3w_core_161;
  wire popcount31_qr3w_core_164;
  wire popcount31_qr3w_core_165;
  wire popcount31_qr3w_core_167;
  wire popcount31_qr3w_core_169;
  wire popcount31_qr3w_core_170;
  wire popcount31_qr3w_core_172;
  wire popcount31_qr3w_core_173;
  wire popcount31_qr3w_core_174;
  wire popcount31_qr3w_core_176;
  wire popcount31_qr3w_core_178;
  wire popcount31_qr3w_core_180;
  wire popcount31_qr3w_core_182;
  wire popcount31_qr3w_core_184;
  wire popcount31_qr3w_core_188;
  wire popcount31_qr3w_core_189;
  wire popcount31_qr3w_core_190;
  wire popcount31_qr3w_core_194;
  wire popcount31_qr3w_core_196;
  wire popcount31_qr3w_core_197;
  wire popcount31_qr3w_core_199;
  wire popcount31_qr3w_core_201;
  wire popcount31_qr3w_core_202;
  wire popcount31_qr3w_core_205;
  wire popcount31_qr3w_core_207;
  wire popcount31_qr3w_core_210;
  wire popcount31_qr3w_core_212;
  wire popcount31_qr3w_core_213;
  wire popcount31_qr3w_core_214_not;
  wire popcount31_qr3w_core_217;

  assign popcount31_qr3w_core_033 = ~(input_a[19] | input_a[4]);
  assign popcount31_qr3w_core_034 = ~(input_a[17] & input_a[4]);
  assign popcount31_qr3w_core_035 = input_a[30] | input_a[6];
  assign popcount31_qr3w_core_037 = input_a[21] ^ input_a[21];
  assign popcount31_qr3w_core_039 = ~(input_a[26] & input_a[15]);
  assign popcount31_qr3w_core_040 = input_a[13] ^ input_a[23];
  assign popcount31_qr3w_core_042 = input_a[21] | input_a[13];
  assign popcount31_qr3w_core_043 = ~(input_a[20] & input_a[24]);
  assign popcount31_qr3w_core_044 = input_a[26] ^ input_a[0];
  assign popcount31_qr3w_core_045 = input_a[30] | input_a[19];
  assign popcount31_qr3w_core_046 = input_a[12] | input_a[28];
  assign popcount31_qr3w_core_048 = ~(input_a[23] ^ input_a[7]);
  assign popcount31_qr3w_core_049 = ~(input_a[13] & input_a[1]);
  assign popcount31_qr3w_core_050 = input_a[26] ^ input_a[10];
  assign popcount31_qr3w_core_051 = input_a[9] | input_a[9];
  assign popcount31_qr3w_core_052 = input_a[24] & input_a[10];
  assign popcount31_qr3w_core_053 = ~(input_a[0] | input_a[30]);
  assign popcount31_qr3w_core_054 = ~input_a[19];
  assign popcount31_qr3w_core_058 = ~(input_a[9] & input_a[9]);
  assign popcount31_qr3w_core_059 = ~input_a[2];
  assign popcount31_qr3w_core_060 = ~input_a[8];
  assign popcount31_qr3w_core_062 = input_a[7] & input_a[27];
  assign popcount31_qr3w_core_064 = input_a[18] ^ input_a[26];
  assign popcount31_qr3w_core_066 = input_a[8] & input_a[21];
  assign popcount31_qr3w_core_069 = ~(input_a[5] | input_a[14]);
  assign popcount31_qr3w_core_073 = input_a[10] ^ input_a[20];
  assign popcount31_qr3w_core_075 = ~input_a[24];
  assign popcount31_qr3w_core_076 = ~input_a[24];
  assign popcount31_qr3w_core_078 = ~(input_a[22] ^ input_a[24]);
  assign popcount31_qr3w_core_079 = input_a[13] & input_a[8];
  assign popcount31_qr3w_core_081 = input_a[2] & input_a[12];
  assign popcount31_qr3w_core_082 = input_a[8] & input_a[1];
  assign popcount31_qr3w_core_086 = ~(input_a[30] ^ input_a[7]);
  assign popcount31_qr3w_core_088 = input_a[29] | input_a[10];
  assign popcount31_qr3w_core_091 = input_a[15] & input_a[8];
  assign popcount31_qr3w_core_093 = ~(input_a[28] & input_a[4]);
  assign popcount31_qr3w_core_096 = ~(input_a[20] | input_a[21]);
  assign popcount31_qr3w_core_098 = ~(input_a[28] ^ input_a[18]);
  assign popcount31_qr3w_core_099 = ~(input_a[17] & input_a[3]);
  assign popcount31_qr3w_core_100 = ~(input_a[27] & input_a[10]);
  assign popcount31_qr3w_core_101 = input_a[20] | input_a[10];
  assign popcount31_qr3w_core_102 = ~input_a[5];
  assign popcount31_qr3w_core_103 = ~(input_a[6] ^ input_a[19]);
  assign popcount31_qr3w_core_104 = ~(input_a[1] ^ input_a[2]);
  assign popcount31_qr3w_core_105 = ~input_a[25];
  assign popcount31_qr3w_core_106 = input_a[1] | input_a[7];
  assign popcount31_qr3w_core_107 = input_a[27] & input_a[3];
  assign popcount31_qr3w_core_108 = input_a[20] | input_a[26];
  assign popcount31_qr3w_core_111 = ~input_a[25];
  assign popcount31_qr3w_core_113 = input_a[27] & input_a[11];
  assign popcount31_qr3w_core_114 = ~input_a[14];
  assign popcount31_qr3w_core_115 = ~(input_a[17] | input_a[15]);
  assign popcount31_qr3w_core_116 = input_a[24] & input_a[11];
  assign popcount31_qr3w_core_119 = ~(input_a[2] | input_a[11]);
  assign popcount31_qr3w_core_120 = ~(input_a[17] ^ input_a[24]);
  assign popcount31_qr3w_core_122 = input_a[25] & input_a[15];
  assign popcount31_qr3w_core_125 = input_a[23] ^ input_a[16];
  assign popcount31_qr3w_core_126 = ~(input_a[28] ^ input_a[6]);
  assign popcount31_qr3w_core_128 = input_a[1] & input_a[11];
  assign popcount31_qr3w_core_129 = input_a[2] | input_a[20];
  assign popcount31_qr3w_core_130 = input_a[11] ^ input_a[5];
  assign popcount31_qr3w_core_131 = ~(input_a[25] ^ input_a[21]);
  assign popcount31_qr3w_core_132 = ~input_a[18];
  assign popcount31_qr3w_core_134 = ~(input_a[13] ^ input_a[26]);
  assign popcount31_qr3w_core_135 = ~(input_a[24] | input_a[7]);
  assign popcount31_qr3w_core_136 = ~(input_a[23] & input_a[2]);
  assign popcount31_qr3w_core_137 = ~(input_a[28] & input_a[4]);
  assign popcount31_qr3w_core_140 = ~(input_a[12] | input_a[23]);
  assign popcount31_qr3w_core_141 = input_a[20] ^ input_a[27];
  assign popcount31_qr3w_core_143 = ~(input_a[16] | input_a[23]);
  assign popcount31_qr3w_core_152 = input_a[14] | input_a[16];
  assign popcount31_qr3w_core_154_not = ~input_a[13];
  assign popcount31_qr3w_core_156 = input_a[3] ^ input_a[4];
  assign popcount31_qr3w_core_158 = input_a[4] ^ input_a[8];
  assign popcount31_qr3w_core_160 = ~(input_a[8] | input_a[21]);
  assign popcount31_qr3w_core_161 = ~(input_a[5] ^ input_a[14]);
  assign popcount31_qr3w_core_164 = input_a[21] | input_a[2];
  assign popcount31_qr3w_core_165 = input_a[17] | input_a[17];
  assign popcount31_qr3w_core_167 = ~(input_a[22] | input_a[25]);
  assign popcount31_qr3w_core_169 = input_a[26] | input_a[9];
  assign popcount31_qr3w_core_170 = ~(input_a[11] ^ input_a[25]);
  assign popcount31_qr3w_core_172 = ~(input_a[17] | input_a[13]);
  assign popcount31_qr3w_core_173 = input_a[25] ^ input_a[9];
  assign popcount31_qr3w_core_174 = input_a[0] ^ input_a[17];
  assign popcount31_qr3w_core_176 = ~(input_a[27] | input_a[24]);
  assign popcount31_qr3w_core_178 = ~input_a[26];
  assign popcount31_qr3w_core_180 = ~(input_a[1] | input_a[3]);
  assign popcount31_qr3w_core_182 = ~(input_a[24] & input_a[14]);
  assign popcount31_qr3w_core_184 = input_a[8] | input_a[13];
  assign popcount31_qr3w_core_188 = input_a[8] | input_a[29];
  assign popcount31_qr3w_core_189 = input_a[20] ^ input_a[11];
  assign popcount31_qr3w_core_190 = ~input_a[27];
  assign popcount31_qr3w_core_194 = input_a[13] & input_a[9];
  assign popcount31_qr3w_core_196 = ~(input_a[3] & input_a[10]);
  assign popcount31_qr3w_core_197 = ~input_a[8];
  assign popcount31_qr3w_core_199 = ~(input_a[8] ^ input_a[18]);
  assign popcount31_qr3w_core_201 = input_a[28] ^ input_a[25];
  assign popcount31_qr3w_core_202 = ~(input_a[14] | input_a[25]);
  assign popcount31_qr3w_core_205 = popcount31_qr3w_core_105 | popcount31_qr3w_core_190;
  assign popcount31_qr3w_core_207 = ~(input_a[22] | input_a[19]);
  assign popcount31_qr3w_core_210 = input_a[25] ^ input_a[27];
  assign popcount31_qr3w_core_212 = popcount31_qr3w_core_210 ^ popcount31_qr3w_core_205;
  assign popcount31_qr3w_core_213 = ~(input_a[2] ^ input_a[26]);
  assign popcount31_qr3w_core_214_not = ~input_a[13];
  assign popcount31_qr3w_core_217 = input_a[27] | input_a[25];

  assign popcount31_qr3w_out[0] = input_a[2];
  assign popcount31_qr3w_out[1] = 1'b1;
  assign popcount31_qr3w_out[2] = popcount31_qr3w_core_212;
  assign popcount31_qr3w_out[3] = popcount31_qr3w_core_212;
  assign popcount31_qr3w_out[4] = popcount31_qr3w_core_217;
endmodule