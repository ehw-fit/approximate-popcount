// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.51489
// WCE=21.0
// EP=0.938456%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_6x39(input [24:0] input_a, output [4:0] popcount25_6x39_out);
  wire popcount25_6x39_core_028;
  wire popcount25_6x39_core_029;
  wire popcount25_6x39_core_030;
  wire popcount25_6x39_core_032;
  wire popcount25_6x39_core_033;
  wire popcount25_6x39_core_035;
  wire popcount25_6x39_core_036;
  wire popcount25_6x39_core_037;
  wire popcount25_6x39_core_041;
  wire popcount25_6x39_core_043;
  wire popcount25_6x39_core_044;
  wire popcount25_6x39_core_048;
  wire popcount25_6x39_core_051;
  wire popcount25_6x39_core_052_not;
  wire popcount25_6x39_core_057;
  wire popcount25_6x39_core_058;
  wire popcount25_6x39_core_064;
  wire popcount25_6x39_core_065;
  wire popcount25_6x39_core_067;
  wire popcount25_6x39_core_069;
  wire popcount25_6x39_core_070;
  wire popcount25_6x39_core_071;
  wire popcount25_6x39_core_072;
  wire popcount25_6x39_core_073;
  wire popcount25_6x39_core_076;
  wire popcount25_6x39_core_077;
  wire popcount25_6x39_core_078;
  wire popcount25_6x39_core_079;
  wire popcount25_6x39_core_080;
  wire popcount25_6x39_core_083;
  wire popcount25_6x39_core_086;
  wire popcount25_6x39_core_087;
  wire popcount25_6x39_core_088;
  wire popcount25_6x39_core_090;
  wire popcount25_6x39_core_092;
  wire popcount25_6x39_core_093;
  wire popcount25_6x39_core_097;
  wire popcount25_6x39_core_098;
  wire popcount25_6x39_core_100;
  wire popcount25_6x39_core_103;
  wire popcount25_6x39_core_104;
  wire popcount25_6x39_core_105;
  wire popcount25_6x39_core_106;
  wire popcount25_6x39_core_107;
  wire popcount25_6x39_core_108;
  wire popcount25_6x39_core_111;
  wire popcount25_6x39_core_112;
  wire popcount25_6x39_core_115;
  wire popcount25_6x39_core_116;
  wire popcount25_6x39_core_118;
  wire popcount25_6x39_core_119;
  wire popcount25_6x39_core_120;
  wire popcount25_6x39_core_122;
  wire popcount25_6x39_core_123;
  wire popcount25_6x39_core_125;
  wire popcount25_6x39_core_126;
  wire popcount25_6x39_core_127;
  wire popcount25_6x39_core_128;
  wire popcount25_6x39_core_129;
  wire popcount25_6x39_core_130;
  wire popcount25_6x39_core_131;
  wire popcount25_6x39_core_132;
  wire popcount25_6x39_core_133;
  wire popcount25_6x39_core_137_not;
  wire popcount25_6x39_core_138;
  wire popcount25_6x39_core_139;
  wire popcount25_6x39_core_140;
  wire popcount25_6x39_core_142;
  wire popcount25_6x39_core_143;
  wire popcount25_6x39_core_144;
  wire popcount25_6x39_core_147;
  wire popcount25_6x39_core_150;
  wire popcount25_6x39_core_152;
  wire popcount25_6x39_core_157;
  wire popcount25_6x39_core_158;
  wire popcount25_6x39_core_159_not;
  wire popcount25_6x39_core_163;
  wire popcount25_6x39_core_165;
  wire popcount25_6x39_core_166;
  wire popcount25_6x39_core_167;
  wire popcount25_6x39_core_168;
  wire popcount25_6x39_core_170;
  wire popcount25_6x39_core_172;
  wire popcount25_6x39_core_173;
  wire popcount25_6x39_core_175;
  wire popcount25_6x39_core_176;
  wire popcount25_6x39_core_178;
  wire popcount25_6x39_core_179;
  wire popcount25_6x39_core_180;
  wire popcount25_6x39_core_181;
  wire popcount25_6x39_core_182;

  assign popcount25_6x39_core_028 = ~(input_a[11] ^ input_a[18]);
  assign popcount25_6x39_core_029 = input_a[6] & input_a[18];
  assign popcount25_6x39_core_030 = ~(input_a[21] ^ input_a[1]);
  assign popcount25_6x39_core_032 = ~(input_a[12] & input_a[2]);
  assign popcount25_6x39_core_033 = ~(input_a[23] | input_a[9]);
  assign popcount25_6x39_core_035 = ~(input_a[21] & input_a[5]);
  assign popcount25_6x39_core_036 = ~(input_a[16] & input_a[16]);
  assign popcount25_6x39_core_037 = input_a[4] & input_a[24];
  assign popcount25_6x39_core_041 = input_a[3] | input_a[16];
  assign popcount25_6x39_core_043 = input_a[7] & input_a[13];
  assign popcount25_6x39_core_044 = ~(input_a[4] | input_a[9]);
  assign popcount25_6x39_core_048 = ~(input_a[6] ^ input_a[18]);
  assign popcount25_6x39_core_051 = input_a[5] & input_a[17];
  assign popcount25_6x39_core_052_not = ~input_a[21];
  assign popcount25_6x39_core_057 = input_a[0] & input_a[17];
  assign popcount25_6x39_core_058 = ~input_a[11];
  assign popcount25_6x39_core_064 = ~(input_a[16] & input_a[1]);
  assign popcount25_6x39_core_065 = ~(input_a[1] ^ input_a[6]);
  assign popcount25_6x39_core_067 = input_a[14] ^ input_a[17];
  assign popcount25_6x39_core_069 = ~(input_a[16] | input_a[0]);
  assign popcount25_6x39_core_070 = ~input_a[23];
  assign popcount25_6x39_core_071 = ~(input_a[12] & input_a[19]);
  assign popcount25_6x39_core_072 = ~input_a[10];
  assign popcount25_6x39_core_073 = ~(input_a[18] | input_a[7]);
  assign popcount25_6x39_core_076 = ~(input_a[2] & input_a[23]);
  assign popcount25_6x39_core_077 = input_a[16] ^ input_a[3];
  assign popcount25_6x39_core_078 = input_a[6] & input_a[3];
  assign popcount25_6x39_core_079 = ~(input_a[23] & input_a[12]);
  assign popcount25_6x39_core_080 = ~(input_a[17] | input_a[13]);
  assign popcount25_6x39_core_083 = ~input_a[11];
  assign popcount25_6x39_core_086 = input_a[24] & input_a[9];
  assign popcount25_6x39_core_087 = input_a[18] ^ input_a[14];
  assign popcount25_6x39_core_088 = ~(input_a[2] ^ input_a[11]);
  assign popcount25_6x39_core_090 = input_a[5] ^ input_a[17];
  assign popcount25_6x39_core_092 = ~(input_a[15] | input_a[15]);
  assign popcount25_6x39_core_093 = ~(input_a[8] | input_a[22]);
  assign popcount25_6x39_core_097 = ~(input_a[8] ^ input_a[13]);
  assign popcount25_6x39_core_098 = input_a[13] ^ input_a[6];
  assign popcount25_6x39_core_100 = ~(input_a[4] | input_a[15]);
  assign popcount25_6x39_core_103 = input_a[19] ^ input_a[6];
  assign popcount25_6x39_core_104 = input_a[12] ^ input_a[0];
  assign popcount25_6x39_core_105 = input_a[4] & input_a[18];
  assign popcount25_6x39_core_106 = ~(input_a[9] | input_a[19]);
  assign popcount25_6x39_core_107 = ~(input_a[5] | input_a[15]);
  assign popcount25_6x39_core_108 = ~(input_a[20] ^ input_a[11]);
  assign popcount25_6x39_core_111 = ~input_a[17];
  assign popcount25_6x39_core_112 = input_a[23] & input_a[16];
  assign popcount25_6x39_core_115 = ~(input_a[20] ^ input_a[10]);
  assign popcount25_6x39_core_116 = input_a[24] ^ input_a[8];
  assign popcount25_6x39_core_118 = ~(input_a[12] | input_a[0]);
  assign popcount25_6x39_core_119 = ~(input_a[23] ^ input_a[18]);
  assign popcount25_6x39_core_120 = ~(input_a[6] | input_a[22]);
  assign popcount25_6x39_core_122 = ~(input_a[14] ^ input_a[23]);
  assign popcount25_6x39_core_123 = ~(input_a[11] ^ input_a[13]);
  assign popcount25_6x39_core_125 = input_a[22] ^ input_a[5];
  assign popcount25_6x39_core_126 = ~(input_a[4] ^ input_a[23]);
  assign popcount25_6x39_core_127 = input_a[19] | input_a[18];
  assign popcount25_6x39_core_128 = ~(input_a[8] ^ input_a[13]);
  assign popcount25_6x39_core_129 = input_a[16] | input_a[10];
  assign popcount25_6x39_core_130 = ~(input_a[3] & input_a[15]);
  assign popcount25_6x39_core_131 = input_a[20] ^ input_a[17];
  assign popcount25_6x39_core_132 = ~input_a[12];
  assign popcount25_6x39_core_133 = input_a[0] & input_a[19];
  assign popcount25_6x39_core_137_not = ~input_a[13];
  assign popcount25_6x39_core_138 = input_a[15] | input_a[8];
  assign popcount25_6x39_core_139 = input_a[0] & input_a[23];
  assign popcount25_6x39_core_140 = input_a[5] & input_a[23];
  assign popcount25_6x39_core_142 = input_a[6] ^ input_a[24];
  assign popcount25_6x39_core_143 = input_a[8] ^ input_a[21];
  assign popcount25_6x39_core_144 = ~input_a[2];
  assign popcount25_6x39_core_147 = input_a[8] ^ input_a[20];
  assign popcount25_6x39_core_150 = ~(input_a[21] ^ input_a[17]);
  assign popcount25_6x39_core_152 = input_a[5] | input_a[1];
  assign popcount25_6x39_core_157 = ~(input_a[8] ^ input_a[21]);
  assign popcount25_6x39_core_158 = ~(input_a[22] ^ input_a[2]);
  assign popcount25_6x39_core_159_not = ~input_a[7];
  assign popcount25_6x39_core_163 = ~(input_a[19] & input_a[10]);
  assign popcount25_6x39_core_165 = input_a[6] | input_a[2];
  assign popcount25_6x39_core_166 = ~(input_a[19] & input_a[13]);
  assign popcount25_6x39_core_167 = input_a[11] | input_a[3];
  assign popcount25_6x39_core_168 = ~(input_a[2] & input_a[2]);
  assign popcount25_6x39_core_170 = input_a[9] | input_a[2];
  assign popcount25_6x39_core_172 = ~(input_a[19] | input_a[17]);
  assign popcount25_6x39_core_173 = input_a[20] & input_a[21];
  assign popcount25_6x39_core_175 = ~(input_a[6] | input_a[20]);
  assign popcount25_6x39_core_176 = ~(input_a[17] ^ input_a[7]);
  assign popcount25_6x39_core_178 = ~(input_a[9] ^ input_a[3]);
  assign popcount25_6x39_core_179 = ~(input_a[13] ^ input_a[11]);
  assign popcount25_6x39_core_180 = input_a[6] & input_a[8];
  assign popcount25_6x39_core_181 = input_a[10] & input_a[0];
  assign popcount25_6x39_core_182 = ~(input_a[7] | input_a[7]);

  assign popcount25_6x39_out[0] = input_a[12];
  assign popcount25_6x39_out[1] = input_a[1];
  assign popcount25_6x39_out[2] = input_a[24];
  assign popcount25_6x39_out[3] = input_a[17];
  assign popcount25_6x39_out[4] = 1'b0;
endmodule