// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.6455
// WCE=14.0
// EP=0.810564%
// Printed PDK parameters:
//  Area=38692770.0
//  Delay=63379108.0
//  Power=1762300.0

module popcount33_t3tt(input [32:0] input_a, output [5:0] popcount33_t3tt_out);
  wire popcount33_t3tt_core_035;
  wire popcount33_t3tt_core_036;
  wire popcount33_t3tt_core_037;
  wire popcount33_t3tt_core_038;
  wire popcount33_t3tt_core_041;
  wire popcount33_t3tt_core_042;
  wire popcount33_t3tt_core_043;
  wire popcount33_t3tt_core_044;
  wire popcount33_t3tt_core_045;
  wire popcount33_t3tt_core_046;
  wire popcount33_t3tt_core_047;
  wire popcount33_t3tt_core_049;
  wire popcount33_t3tt_core_050;
  wire popcount33_t3tt_core_052;
  wire popcount33_t3tt_core_053;
  wire popcount33_t3tt_core_055;
  wire popcount33_t3tt_core_058;
  wire popcount33_t3tt_core_059;
  wire popcount33_t3tt_core_060;
  wire popcount33_t3tt_core_061;
  wire popcount33_t3tt_core_062;
  wire popcount33_t3tt_core_063;
  wire popcount33_t3tt_core_066;
  wire popcount33_t3tt_core_067;
  wire popcount33_t3tt_core_069;
  wire popcount33_t3tt_core_070;
  wire popcount33_t3tt_core_073;
  wire popcount33_t3tt_core_076;
  wire popcount33_t3tt_core_081;
  wire popcount33_t3tt_core_082;
  wire popcount33_t3tt_core_083;
  wire popcount33_t3tt_core_084;
  wire popcount33_t3tt_core_085;
  wire popcount33_t3tt_core_086;
  wire popcount33_t3tt_core_087;
  wire popcount33_t3tt_core_088;
  wire popcount33_t3tt_core_089;
  wire popcount33_t3tt_core_092;
  wire popcount33_t3tt_core_093;
  wire popcount33_t3tt_core_094;
  wire popcount33_t3tt_core_095;
  wire popcount33_t3tt_core_096;
  wire popcount33_t3tt_core_097;
  wire popcount33_t3tt_core_100;
  wire popcount33_t3tt_core_101;
  wire popcount33_t3tt_core_102;
  wire popcount33_t3tt_core_104;
  wire popcount33_t3tt_core_105;
  wire popcount33_t3tt_core_106;
  wire popcount33_t3tt_core_107;
  wire popcount33_t3tt_core_108;
  wire popcount33_t3tt_core_109;
  wire popcount33_t3tt_core_110;
  wire popcount33_t3tt_core_111;
  wire popcount33_t3tt_core_112;
  wire popcount33_t3tt_core_113;
  wire popcount33_t3tt_core_114;
  wire popcount33_t3tt_core_117;
  wire popcount33_t3tt_core_119;
  wire popcount33_t3tt_core_120;
  wire popcount33_t3tt_core_121;
  wire popcount33_t3tt_core_123;
  wire popcount33_t3tt_core_125;
  wire popcount33_t3tt_core_126;
  wire popcount33_t3tt_core_127;
  wire popcount33_t3tt_core_129;
  wire popcount33_t3tt_core_130;
  wire popcount33_t3tt_core_131;
  wire popcount33_t3tt_core_132;
  wire popcount33_t3tt_core_133;
  wire popcount33_t3tt_core_134;
  wire popcount33_t3tt_core_135;
  wire popcount33_t3tt_core_136;
  wire popcount33_t3tt_core_138;
  wire popcount33_t3tt_core_139;
  wire popcount33_t3tt_core_141;
  wire popcount33_t3tt_core_142;
  wire popcount33_t3tt_core_143;
  wire popcount33_t3tt_core_144;
  wire popcount33_t3tt_core_152;
  wire popcount33_t3tt_core_153;
  wire popcount33_t3tt_core_154;
  wire popcount33_t3tt_core_155;
  wire popcount33_t3tt_core_156;
  wire popcount33_t3tt_core_160;
  wire popcount33_t3tt_core_162;
  wire popcount33_t3tt_core_163;
  wire popcount33_t3tt_core_165;
  wire popcount33_t3tt_core_167;
  wire popcount33_t3tt_core_169;
  wire popcount33_t3tt_core_171;
  wire popcount33_t3tt_core_173;
  wire popcount33_t3tt_core_174;
  wire popcount33_t3tt_core_175;
  wire popcount33_t3tt_core_176;
  wire popcount33_t3tt_core_177;
  wire popcount33_t3tt_core_179;
  wire popcount33_t3tt_core_180;
  wire popcount33_t3tt_core_182;
  wire popcount33_t3tt_core_183;
  wire popcount33_t3tt_core_184;
  wire popcount33_t3tt_core_187;
  wire popcount33_t3tt_core_189;
  wire popcount33_t3tt_core_190;
  wire popcount33_t3tt_core_192;
  wire popcount33_t3tt_core_193;
  wire popcount33_t3tt_core_197;
  wire popcount33_t3tt_core_198;
  wire popcount33_t3tt_core_199;
  wire popcount33_t3tt_core_201;
  wire popcount33_t3tt_core_203;
  wire popcount33_t3tt_core_204;
  wire popcount33_t3tt_core_205;
  wire popcount33_t3tt_core_206;
  wire popcount33_t3tt_core_207;
  wire popcount33_t3tt_core_209;
  wire popcount33_t3tt_core_213;
  wire popcount33_t3tt_core_215;
  wire popcount33_t3tt_core_217;
  wire popcount33_t3tt_core_218;
  wire popcount33_t3tt_core_219;
  wire popcount33_t3tt_core_220;
  wire popcount33_t3tt_core_221;
  wire popcount33_t3tt_core_222;
  wire popcount33_t3tt_core_223;
  wire popcount33_t3tt_core_224;
  wire popcount33_t3tt_core_225;
  wire popcount33_t3tt_core_226;
  wire popcount33_t3tt_core_227;
  wire popcount33_t3tt_core_228;
  wire popcount33_t3tt_core_229;
  wire popcount33_t3tt_core_230;
  wire popcount33_t3tt_core_231;
  wire popcount33_t3tt_core_232_not;
  wire popcount33_t3tt_core_233;
  wire popcount33_t3tt_core_234;
  wire popcount33_t3tt_core_235;
  wire popcount33_t3tt_core_237;
  wire popcount33_t3tt_core_238;

  assign popcount33_t3tt_core_035 = input_a[0] ^ input_a[1];
  assign popcount33_t3tt_core_036 = input_a[0] & input_a[1];
  assign popcount33_t3tt_core_037 = input_a[20] | input_a[1];
  assign popcount33_t3tt_core_038 = input_a[11] & input_a[7];
  assign popcount33_t3tt_core_041 = popcount33_t3tt_core_036 ^ popcount33_t3tt_core_038;
  assign popcount33_t3tt_core_042 = input_a[0] & popcount33_t3tt_core_038;
  assign popcount33_t3tt_core_043 = popcount33_t3tt_core_041 ^ popcount33_t3tt_core_035;
  assign popcount33_t3tt_core_044 = popcount33_t3tt_core_041 & popcount33_t3tt_core_035;
  assign popcount33_t3tt_core_045 = popcount33_t3tt_core_042 | popcount33_t3tt_core_044;
  assign popcount33_t3tt_core_046 = ~(input_a[20] & input_a[5]);
  assign popcount33_t3tt_core_047 = ~(input_a[10] & input_a[16]);
  assign popcount33_t3tt_core_049 = input_a[17] & input_a[6];
  assign popcount33_t3tt_core_050 = ~(input_a[15] | input_a[17]);
  assign popcount33_t3tt_core_052 = input_a[8] | popcount33_t3tt_core_049;
  assign popcount33_t3tt_core_053 = input_a[21] ^ input_a[7];
  assign popcount33_t3tt_core_055 = ~input_a[21];
  assign popcount33_t3tt_core_058 = input_a[28] & input_a[3];
  assign popcount33_t3tt_core_059 = popcount33_t3tt_core_043 ^ popcount33_t3tt_core_052;
  assign popcount33_t3tt_core_060 = popcount33_t3tt_core_043 & popcount33_t3tt_core_052;
  assign popcount33_t3tt_core_061 = popcount33_t3tt_core_059 ^ popcount33_t3tt_core_058;
  assign popcount33_t3tt_core_062 = popcount33_t3tt_core_059 & popcount33_t3tt_core_058;
  assign popcount33_t3tt_core_063 = popcount33_t3tt_core_060 | popcount33_t3tt_core_062;
  assign popcount33_t3tt_core_066 = popcount33_t3tt_core_045 ^ popcount33_t3tt_core_063;
  assign popcount33_t3tt_core_067 = popcount33_t3tt_core_045 & popcount33_t3tt_core_063;
  assign popcount33_t3tt_core_069 = input_a[4] ^ input_a[9];
  assign popcount33_t3tt_core_070 = input_a[10] & input_a[22];
  assign popcount33_t3tt_core_073 = input_a[5] ^ input_a[6];
  assign popcount33_t3tt_core_076 = ~input_a[0];
  assign popcount33_t3tt_core_081 = input_a[2] ^ input_a[16];
  assign popcount33_t3tt_core_082 = ~(input_a[13] ^ input_a[2]);
  assign popcount33_t3tt_core_083 = input_a[24] & input_a[30];
  assign popcount33_t3tt_core_084 = ~input_a[25];
  assign popcount33_t3tt_core_085 = input_a[16] & input_a[20];
  assign popcount33_t3tt_core_086 = input_a[9] ^ popcount33_t3tt_core_083;
  assign popcount33_t3tt_core_087 = input_a[9] & popcount33_t3tt_core_083;
  assign popcount33_t3tt_core_088 = popcount33_t3tt_core_086 | popcount33_t3tt_core_085;
  assign popcount33_t3tt_core_089 = ~input_a[4];
  assign popcount33_t3tt_core_092 = input_a[32] & input_a[2];
  assign popcount33_t3tt_core_093 = popcount33_t3tt_core_070 ^ popcount33_t3tt_core_088;
  assign popcount33_t3tt_core_094 = popcount33_t3tt_core_070 & popcount33_t3tt_core_088;
  assign popcount33_t3tt_core_095 = popcount33_t3tt_core_093 ^ popcount33_t3tt_core_092;
  assign popcount33_t3tt_core_096 = popcount33_t3tt_core_093 & popcount33_t3tt_core_092;
  assign popcount33_t3tt_core_097 = popcount33_t3tt_core_094 | popcount33_t3tt_core_096;
  assign popcount33_t3tt_core_100 = popcount33_t3tt_core_087 | popcount33_t3tt_core_097;
  assign popcount33_t3tt_core_101 = ~(input_a[23] | input_a[16]);
  assign popcount33_t3tt_core_102 = input_a[4] ^ input_a[12];
  assign popcount33_t3tt_core_104 = input_a[26] & input_a[18];
  assign popcount33_t3tt_core_105 = popcount33_t3tt_core_061 ^ popcount33_t3tt_core_095;
  assign popcount33_t3tt_core_106 = popcount33_t3tt_core_061 & popcount33_t3tt_core_095;
  assign popcount33_t3tt_core_107 = popcount33_t3tt_core_105 ^ popcount33_t3tt_core_104;
  assign popcount33_t3tt_core_108 = popcount33_t3tt_core_105 & popcount33_t3tt_core_104;
  assign popcount33_t3tt_core_109 = popcount33_t3tt_core_106 | popcount33_t3tt_core_108;
  assign popcount33_t3tt_core_110 = popcount33_t3tt_core_066 ^ popcount33_t3tt_core_100;
  assign popcount33_t3tt_core_111 = popcount33_t3tt_core_066 & popcount33_t3tt_core_100;
  assign popcount33_t3tt_core_112 = popcount33_t3tt_core_110 ^ popcount33_t3tt_core_109;
  assign popcount33_t3tt_core_113 = popcount33_t3tt_core_110 & popcount33_t3tt_core_109;
  assign popcount33_t3tt_core_114 = popcount33_t3tt_core_111 | popcount33_t3tt_core_113;
  assign popcount33_t3tt_core_117 = popcount33_t3tt_core_067 | popcount33_t3tt_core_114;
  assign popcount33_t3tt_core_119 = input_a[26] & input_a[23];
  assign popcount33_t3tt_core_120 = ~input_a[11];
  assign popcount33_t3tt_core_121 = input_a[23] & input_a[14];
  assign popcount33_t3tt_core_123 = input_a[19] & input_a[15];
  assign popcount33_t3tt_core_125 = input_a[25] ^ input_a[30];
  assign popcount33_t3tt_core_126 = popcount33_t3tt_core_121 | popcount33_t3tt_core_123;
  assign popcount33_t3tt_core_127 = ~(input_a[6] & input_a[10]);
  assign popcount33_t3tt_core_129 = input_a[21] | input_a[25];
  assign popcount33_t3tt_core_130 = ~(input_a[30] ^ input_a[2]);
  assign popcount33_t3tt_core_131 = ~(input_a[29] & input_a[0]);
  assign popcount33_t3tt_core_132 = input_a[14] & input_a[7];
  assign popcount33_t3tt_core_133 = ~input_a[24];
  assign popcount33_t3tt_core_134 = ~(input_a[17] ^ input_a[12]);
  assign popcount33_t3tt_core_135 = ~(input_a[29] ^ input_a[12]);
  assign popcount33_t3tt_core_136 = ~(input_a[6] ^ input_a[17]);
  assign popcount33_t3tt_core_138 = ~(input_a[28] | input_a[25]);
  assign popcount33_t3tt_core_139 = ~(input_a[14] | input_a[32]);
  assign popcount33_t3tt_core_141 = ~input_a[19];
  assign popcount33_t3tt_core_142 = ~(input_a[15] & input_a[13]);
  assign popcount33_t3tt_core_143 = ~(input_a[27] ^ input_a[17]);
  assign popcount33_t3tt_core_144 = ~popcount33_t3tt_core_126;
  assign popcount33_t3tt_core_152 = ~(input_a[27] | input_a[3]);
  assign popcount33_t3tt_core_153 = input_a[3] ^ input_a[9];
  assign popcount33_t3tt_core_154 = ~(input_a[21] | input_a[11]);
  assign popcount33_t3tt_core_155 = ~(input_a[32] & input_a[32]);
  assign popcount33_t3tt_core_156 = input_a[3] & input_a[20];
  assign popcount33_t3tt_core_160 = ~(input_a[13] ^ input_a[23]);
  assign popcount33_t3tt_core_162 = input_a[21] | input_a[4];
  assign popcount33_t3tt_core_163 = ~input_a[16];
  assign popcount33_t3tt_core_165 = ~(input_a[23] ^ input_a[9]);
  assign popcount33_t3tt_core_167 = input_a[9] | input_a[9];
  assign popcount33_t3tt_core_169 = input_a[29] ^ input_a[11];
  assign popcount33_t3tt_core_171 = input_a[29] | input_a[5];
  assign popcount33_t3tt_core_173 = ~(input_a[3] ^ input_a[11]);
  assign popcount33_t3tt_core_174 = input_a[20] ^ input_a[15];
  assign popcount33_t3tt_core_175 = input_a[31] | popcount33_t3tt_core_171;
  assign popcount33_t3tt_core_176 = input_a[27] ^ input_a[19];
  assign popcount33_t3tt_core_177 = ~popcount33_t3tt_core_175;
  assign popcount33_t3tt_core_179 = input_a[4] | popcount33_t3tt_core_175;
  assign popcount33_t3tt_core_180 = input_a[4] | popcount33_t3tt_core_179;
  assign popcount33_t3tt_core_182 = ~(input_a[23] | input_a[16]);
  assign popcount33_t3tt_core_183 = ~input_a[0];
  assign popcount33_t3tt_core_184 = popcount33_t3tt_core_162 ^ popcount33_t3tt_core_177;
  assign popcount33_t3tt_core_187 = ~(input_a[31] & input_a[13]);
  assign popcount33_t3tt_core_189 = input_a[21] | popcount33_t3tt_core_180;
  assign popcount33_t3tt_core_190 = input_a[32] & input_a[4];
  assign popcount33_t3tt_core_192 = input_a[22] ^ input_a[23];
  assign popcount33_t3tt_core_193 = ~(input_a[28] ^ input_a[31]);
  assign popcount33_t3tt_core_197 = ~(input_a[15] & input_a[9]);
  assign popcount33_t3tt_core_198 = popcount33_t3tt_core_144 ^ popcount33_t3tt_core_184;
  assign popcount33_t3tt_core_199 = popcount33_t3tt_core_144 & popcount33_t3tt_core_184;
  assign popcount33_t3tt_core_201 = ~(input_a[21] | input_a[7]);
  assign popcount33_t3tt_core_203 = popcount33_t3tt_core_126 ^ popcount33_t3tt_core_189;
  assign popcount33_t3tt_core_204 = popcount33_t3tt_core_126 & popcount33_t3tt_core_189;
  assign popcount33_t3tt_core_205 = popcount33_t3tt_core_203 ^ popcount33_t3tt_core_199;
  assign popcount33_t3tt_core_206 = popcount33_t3tt_core_203 & popcount33_t3tt_core_199;
  assign popcount33_t3tt_core_207 = popcount33_t3tt_core_204 | popcount33_t3tt_core_206;
  assign popcount33_t3tt_core_209 = ~input_a[14];
  assign popcount33_t3tt_core_213 = input_a[24] | input_a[22];
  assign popcount33_t3tt_core_215 = ~(input_a[16] ^ input_a[8]);
  assign popcount33_t3tt_core_217 = popcount33_t3tt_core_107 ^ popcount33_t3tt_core_198;
  assign popcount33_t3tt_core_218 = popcount33_t3tt_core_107 & popcount33_t3tt_core_198;
  assign popcount33_t3tt_core_219 = popcount33_t3tt_core_217 ^ input_a[27];
  assign popcount33_t3tt_core_220 = popcount33_t3tt_core_217 & input_a[27];
  assign popcount33_t3tt_core_221 = popcount33_t3tt_core_218 | popcount33_t3tt_core_220;
  assign popcount33_t3tt_core_222 = popcount33_t3tt_core_112 ^ popcount33_t3tt_core_205;
  assign popcount33_t3tt_core_223 = popcount33_t3tt_core_112 & popcount33_t3tt_core_205;
  assign popcount33_t3tt_core_224 = popcount33_t3tt_core_222 ^ popcount33_t3tt_core_221;
  assign popcount33_t3tt_core_225 = popcount33_t3tt_core_222 & popcount33_t3tt_core_221;
  assign popcount33_t3tt_core_226 = popcount33_t3tt_core_223 | popcount33_t3tt_core_225;
  assign popcount33_t3tt_core_227 = popcount33_t3tt_core_117 ^ popcount33_t3tt_core_207;
  assign popcount33_t3tt_core_228 = popcount33_t3tt_core_117 & popcount33_t3tt_core_207;
  assign popcount33_t3tt_core_229 = popcount33_t3tt_core_227 ^ popcount33_t3tt_core_226;
  assign popcount33_t3tt_core_230 = popcount33_t3tt_core_227 & popcount33_t3tt_core_226;
  assign popcount33_t3tt_core_231 = popcount33_t3tt_core_228 | popcount33_t3tt_core_230;
  assign popcount33_t3tt_core_232_not = ~input_a[14];
  assign popcount33_t3tt_core_233 = ~(input_a[1] | input_a[28]);
  assign popcount33_t3tt_core_234 = ~(input_a[15] ^ input_a[28]);
  assign popcount33_t3tt_core_235 = input_a[30] ^ input_a[1];
  assign popcount33_t3tt_core_237 = ~input_a[9];
  assign popcount33_t3tt_core_238 = ~(input_a[5] ^ input_a[4]);

  assign popcount33_t3tt_out[0] = popcount33_t3tt_core_229;
  assign popcount33_t3tt_out[1] = popcount33_t3tt_core_219;
  assign popcount33_t3tt_out[2] = popcount33_t3tt_core_224;
  assign popcount33_t3tt_out[3] = popcount33_t3tt_core_229;
  assign popcount33_t3tt_out[4] = popcount33_t3tt_core_231;
  assign popcount33_t3tt_out[5] = 1'b0;
endmodule