// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.2561
// WCE=5.0
// EP=0.759033%
// Printed PDK parameters:
//  Area=32040143.0
//  Delay=52919116.0
//  Power=1390900.0

module popcount24_8px4(input [23:0] input_a, output [4:0] popcount24_8px4_out);
  wire popcount24_8px4_core_026;
  wire popcount24_8px4_core_028;
  wire popcount24_8px4_core_029;
  wire popcount24_8px4_core_030;
  wire popcount24_8px4_core_033;
  wire popcount24_8px4_core_034;
  wire popcount24_8px4_core_035;
  wire popcount24_8px4_core_036;
  wire popcount24_8px4_core_038;
  wire popcount24_8px4_core_039;
  wire popcount24_8px4_core_040;
  wire popcount24_8px4_core_042;
  wire popcount24_8px4_core_044;
  wire popcount24_8px4_core_045;
  wire popcount24_8px4_core_048;
  wire popcount24_8px4_core_049;
  wire popcount24_8px4_core_051;
  wire popcount24_8px4_core_054;
  wire popcount24_8px4_core_055;
  wire popcount24_8px4_core_056;
  wire popcount24_8px4_core_057;
  wire popcount24_8px4_core_059;
  wire popcount24_8px4_core_060;
  wire popcount24_8px4_core_062;
  wire popcount24_8px4_core_063;
  wire popcount24_8px4_core_064;
  wire popcount24_8px4_core_066;
  wire popcount24_8px4_core_067;
  wire popcount24_8px4_core_068;
  wire popcount24_8px4_core_069;
  wire popcount24_8px4_core_071;
  wire popcount24_8px4_core_072;
  wire popcount24_8px4_core_073;
  wire popcount24_8px4_core_074;
  wire popcount24_8px4_core_076;
  wire popcount24_8px4_core_077;
  wire popcount24_8px4_core_078;
  wire popcount24_8px4_core_081;
  wire popcount24_8px4_core_083;
  wire popcount24_8px4_core_084;
  wire popcount24_8px4_core_087;
  wire popcount24_8px4_core_091;
  wire popcount24_8px4_core_092;
  wire popcount24_8px4_core_093;
  wire popcount24_8px4_core_094;
  wire popcount24_8px4_core_095;
  wire popcount24_8px4_core_096;
  wire popcount24_8px4_core_097;
  wire popcount24_8px4_core_098;
  wire popcount24_8px4_core_099;
  wire popcount24_8px4_core_100;
  wire popcount24_8px4_core_101;
  wire popcount24_8px4_core_102;
  wire popcount24_8px4_core_103;
  wire popcount24_8px4_core_104;
  wire popcount24_8px4_core_105;
  wire popcount24_8px4_core_106;
  wire popcount24_8px4_core_107;
  wire popcount24_8px4_core_108;
  wire popcount24_8px4_core_109;
  wire popcount24_8px4_core_111_not;
  wire popcount24_8px4_core_113;
  wire popcount24_8px4_core_114;
  wire popcount24_8px4_core_115;
  wire popcount24_8px4_core_116;
  wire popcount24_8px4_core_117;
  wire popcount24_8px4_core_118;
  wire popcount24_8px4_core_119;
  wire popcount24_8px4_core_120;
  wire popcount24_8px4_core_121;
  wire popcount24_8px4_core_122;
  wire popcount24_8px4_core_124;
  wire popcount24_8px4_core_125;
  wire popcount24_8px4_core_128;
  wire popcount24_8px4_core_129;
  wire popcount24_8px4_core_130;
  wire popcount24_8px4_core_131;
  wire popcount24_8px4_core_132;
  wire popcount24_8px4_core_133;
  wire popcount24_8px4_core_135;
  wire popcount24_8px4_core_137;
  wire popcount24_8px4_core_140;
  wire popcount24_8px4_core_141;
  wire popcount24_8px4_core_142;
  wire popcount24_8px4_core_144;
  wire popcount24_8px4_core_146;
  wire popcount24_8px4_core_147;
  wire popcount24_8px4_core_148;
  wire popcount24_8px4_core_149;
  wire popcount24_8px4_core_150;
  wire popcount24_8px4_core_152;
  wire popcount24_8px4_core_154;
  wire popcount24_8px4_core_155;
  wire popcount24_8px4_core_156;
  wire popcount24_8px4_core_157;
  wire popcount24_8px4_core_158;
  wire popcount24_8px4_core_159;
  wire popcount24_8px4_core_160;
  wire popcount24_8px4_core_161;
  wire popcount24_8px4_core_162;
  wire popcount24_8px4_core_163;
  wire popcount24_8px4_core_164;
  wire popcount24_8px4_core_165;
  wire popcount24_8px4_core_166;
  wire popcount24_8px4_core_167;
  wire popcount24_8px4_core_168;
  wire popcount24_8px4_core_169;
  wire popcount24_8px4_core_170;
  wire popcount24_8px4_core_171;
  wire popcount24_8px4_core_172;
  wire popcount24_8px4_core_174;
  wire popcount24_8px4_core_177_not;

  assign popcount24_8px4_core_026 = input_a[15] | input_a[5];
  assign popcount24_8px4_core_028 = input_a[5] ^ input_a[5];
  assign popcount24_8px4_core_029 = input_a[2] ^ input_a[9];
  assign popcount24_8px4_core_030 = input_a[19] | input_a[18];
  assign popcount24_8px4_core_033 = input_a[3] | input_a[23];
  assign popcount24_8px4_core_034 = ~(input_a[16] & input_a[7]);
  assign popcount24_8px4_core_035 = ~input_a[14];
  assign popcount24_8px4_core_036 = ~(input_a[11] ^ input_a[20]);
  assign popcount24_8px4_core_038 = input_a[0] ^ input_a[5];
  assign popcount24_8px4_core_039 = ~(input_a[1] & input_a[16]);
  assign popcount24_8px4_core_040 = ~input_a[14];
  assign popcount24_8px4_core_042 = ~(input_a[16] & input_a[13]);
  assign popcount24_8px4_core_044 = input_a[19] | input_a[10];
  assign popcount24_8px4_core_045 = ~input_a[7];
  assign popcount24_8px4_core_048 = ~(input_a[16] ^ input_a[5]);
  assign popcount24_8px4_core_049 = ~input_a[3];
  assign popcount24_8px4_core_051 = input_a[12] ^ input_a[0];
  assign popcount24_8px4_core_054 = ~input_a[16];
  assign popcount24_8px4_core_055 = ~(input_a[15] ^ input_a[6]);
  assign popcount24_8px4_core_056 = input_a[9] & input_a[5];
  assign popcount24_8px4_core_057 = ~(input_a[15] | input_a[16]);
  assign popcount24_8px4_core_059 = ~input_a[8];
  assign popcount24_8px4_core_060 = input_a[14] ^ input_a[19];
  assign popcount24_8px4_core_062 = ~input_a[6];
  assign popcount24_8px4_core_063 = ~input_a[17];
  assign popcount24_8px4_core_064 = input_a[3] ^ input_a[16];
  assign popcount24_8px4_core_066 = input_a[2] & input_a[9];
  assign popcount24_8px4_core_067 = input_a[17] & input_a[3];
  assign popcount24_8px4_core_068 = input_a[11] & input_a[9];
  assign popcount24_8px4_core_069 = input_a[9] & input_a[12];
  assign popcount24_8px4_core_071 = input_a[6] & input_a[2];
  assign popcount24_8px4_core_072 = input_a[1] & input_a[18];
  assign popcount24_8px4_core_073 = ~input_a[19];
  assign popcount24_8px4_core_074 = popcount24_8px4_core_038 ^ popcount24_8px4_core_062;
  assign popcount24_8px4_core_076 = input_a[0] ^ input_a[6];
  assign popcount24_8px4_core_077 = input_a[0] & input_a[6];
  assign popcount24_8px4_core_078 = popcount24_8px4_core_076 | popcount24_8px4_core_038;
  assign popcount24_8px4_core_081 = ~(input_a[4] ^ input_a[20]);
  assign popcount24_8px4_core_083 = ~(input_a[5] & popcount24_8px4_core_077);
  assign popcount24_8px4_core_084 = input_a[5] & popcount24_8px4_core_077;
  assign popcount24_8px4_core_087 = ~(input_a[3] | input_a[2]);
  assign popcount24_8px4_core_091 = input_a[23] ^ input_a[6];
  assign popcount24_8px4_core_092 = input_a[13] & input_a[19];
  assign popcount24_8px4_core_093 = ~input_a[4];
  assign popcount24_8px4_core_094 = input_a[12] & input_a[9];
  assign popcount24_8px4_core_095 = popcount24_8px4_core_092 | popcount24_8px4_core_094;
  assign popcount24_8px4_core_096 = ~(input_a[11] & input_a[3]);
  assign popcount24_8px4_core_097 = input_a[16] | input_a[17];
  assign popcount24_8px4_core_098 = input_a[16] & input_a[17];
  assign popcount24_8px4_core_099 = input_a[23] & input_a[16];
  assign popcount24_8px4_core_100 = input_a[15] & popcount24_8px4_core_097;
  assign popcount24_8px4_core_101 = popcount24_8px4_core_098 | popcount24_8px4_core_100;
  assign popcount24_8px4_core_102 = ~(input_a[10] | input_a[3]);
  assign popcount24_8px4_core_103 = ~(input_a[12] ^ input_a[10]);
  assign popcount24_8px4_core_104 = input_a[2] & input_a[8];
  assign popcount24_8px4_core_105 = popcount24_8px4_core_095 ^ popcount24_8px4_core_101;
  assign popcount24_8px4_core_106 = popcount24_8px4_core_095 & popcount24_8px4_core_101;
  assign popcount24_8px4_core_107 = popcount24_8px4_core_105 ^ popcount24_8px4_core_104;
  assign popcount24_8px4_core_108 = popcount24_8px4_core_105 & popcount24_8px4_core_104;
  assign popcount24_8px4_core_109 = popcount24_8px4_core_106 | popcount24_8px4_core_108;
  assign popcount24_8px4_core_111_not = ~input_a[11];
  assign popcount24_8px4_core_113 = ~(input_a[0] | input_a[9]);
  assign popcount24_8px4_core_114 = ~(input_a[22] & input_a[7]);
  assign popcount24_8px4_core_115 = input_a[11] & input_a[18];
  assign popcount24_8px4_core_116 = input_a[3] & input_a[20];
  assign popcount24_8px4_core_117 = ~(input_a[14] | input_a[15]);
  assign popcount24_8px4_core_118 = input_a[18] & input_a[1];
  assign popcount24_8px4_core_119 = popcount24_8px4_core_116 | popcount24_8px4_core_118;
  assign popcount24_8px4_core_120 = input_a[15] ^ input_a[11];
  assign popcount24_8px4_core_121 = input_a[13] ^ input_a[15];
  assign popcount24_8px4_core_122 = input_a[22] & input_a[23];
  assign popcount24_8px4_core_124 = input_a[21] & input_a[10];
  assign popcount24_8px4_core_125 = popcount24_8px4_core_122 | popcount24_8px4_core_124;
  assign popcount24_8px4_core_128 = input_a[11] & input_a[7];
  assign popcount24_8px4_core_129 = popcount24_8px4_core_119 ^ popcount24_8px4_core_125;
  assign popcount24_8px4_core_130 = popcount24_8px4_core_119 & popcount24_8px4_core_125;
  assign popcount24_8px4_core_131 = popcount24_8px4_core_129 ^ popcount24_8px4_core_128;
  assign popcount24_8px4_core_132 = popcount24_8px4_core_129 & popcount24_8px4_core_128;
  assign popcount24_8px4_core_133 = popcount24_8px4_core_130 | popcount24_8px4_core_132;
  assign popcount24_8px4_core_135 = ~input_a[11];
  assign popcount24_8px4_core_137 = input_a[16] ^ input_a[19];
  assign popcount24_8px4_core_140 = ~(input_a[11] | input_a[14]);
  assign popcount24_8px4_core_141 = popcount24_8px4_core_107 ^ popcount24_8px4_core_131;
  assign popcount24_8px4_core_142 = popcount24_8px4_core_107 & popcount24_8px4_core_131;
  assign popcount24_8px4_core_144 = ~(input_a[8] ^ input_a[21]);
  assign popcount24_8px4_core_146 = popcount24_8px4_core_109 ^ popcount24_8px4_core_133;
  assign popcount24_8px4_core_147 = popcount24_8px4_core_109 & popcount24_8px4_core_133;
  assign popcount24_8px4_core_148 = popcount24_8px4_core_146 ^ popcount24_8px4_core_142;
  assign popcount24_8px4_core_149 = popcount24_8px4_core_146 & popcount24_8px4_core_142;
  assign popcount24_8px4_core_150 = popcount24_8px4_core_147 | popcount24_8px4_core_149;
  assign popcount24_8px4_core_152 = input_a[17] ^ input_a[14];
  assign popcount24_8px4_core_154 = ~input_a[11];
  assign popcount24_8px4_core_155 = ~input_a[1];
  assign popcount24_8px4_core_156 = input_a[5] | input_a[19];
  assign popcount24_8px4_core_157 = popcount24_8px4_core_074 & input_a[4];
  assign popcount24_8px4_core_158 = popcount24_8px4_core_078 ^ popcount24_8px4_core_141;
  assign popcount24_8px4_core_159 = popcount24_8px4_core_078 & popcount24_8px4_core_141;
  assign popcount24_8px4_core_160 = popcount24_8px4_core_158 ^ popcount24_8px4_core_157;
  assign popcount24_8px4_core_161 = popcount24_8px4_core_158 & popcount24_8px4_core_157;
  assign popcount24_8px4_core_162 = popcount24_8px4_core_159 | popcount24_8px4_core_161;
  assign popcount24_8px4_core_163 = popcount24_8px4_core_083 ^ popcount24_8px4_core_148;
  assign popcount24_8px4_core_164 = popcount24_8px4_core_083 & popcount24_8px4_core_148;
  assign popcount24_8px4_core_165 = popcount24_8px4_core_163 ^ popcount24_8px4_core_162;
  assign popcount24_8px4_core_166 = popcount24_8px4_core_163 & popcount24_8px4_core_162;
  assign popcount24_8px4_core_167 = popcount24_8px4_core_164 | popcount24_8px4_core_166;
  assign popcount24_8px4_core_168 = popcount24_8px4_core_084 ^ popcount24_8px4_core_150;
  assign popcount24_8px4_core_169 = popcount24_8px4_core_084 & popcount24_8px4_core_150;
  assign popcount24_8px4_core_170 = popcount24_8px4_core_168 ^ popcount24_8px4_core_167;
  assign popcount24_8px4_core_171 = popcount24_8px4_core_168 & popcount24_8px4_core_167;
  assign popcount24_8px4_core_172 = popcount24_8px4_core_169 | popcount24_8px4_core_171;
  assign popcount24_8px4_core_174 = ~input_a[9];
  assign popcount24_8px4_core_177_not = ~input_a[10];

  assign popcount24_8px4_out[0] = input_a[14];
  assign popcount24_8px4_out[1] = popcount24_8px4_core_160;
  assign popcount24_8px4_out[2] = popcount24_8px4_core_165;
  assign popcount24_8px4_out[3] = popcount24_8px4_core_170;
  assign popcount24_8px4_out[4] = popcount24_8px4_core_172;
endmodule