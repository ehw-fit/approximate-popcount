// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.44133
// WCE=23.0
// EP=0.908798%
// Printed PDK parameters:
//  Area=65340486.0
//  Delay=67018788.0
//  Power=2878200.0

module popcount35_c6d4(input [34:0] input_a, output [5:0] popcount35_c6d4_out);
  wire popcount35_c6d4_core_037;
  wire popcount35_c6d4_core_039;
  wire popcount35_c6d4_core_043;
  wire popcount35_c6d4_core_045;
  wire popcount35_c6d4_core_046;
  wire popcount35_c6d4_core_047;
  wire popcount35_c6d4_core_048;
  wire popcount35_c6d4_core_050;
  wire popcount35_c6d4_core_051;
  wire popcount35_c6d4_core_052;
  wire popcount35_c6d4_core_053;
  wire popcount35_c6d4_core_056;
  wire popcount35_c6d4_core_057;
  wire popcount35_c6d4_core_059_not;
  wire popcount35_c6d4_core_062;
  wire popcount35_c6d4_core_063;
  wire popcount35_c6d4_core_064;
  wire popcount35_c6d4_core_065;
  wire popcount35_c6d4_core_066;
  wire popcount35_c6d4_core_067;
  wire popcount35_c6d4_core_068;
  wire popcount35_c6d4_core_069;
  wire popcount35_c6d4_core_070;
  wire popcount35_c6d4_core_071;
  wire popcount35_c6d4_core_072;
  wire popcount35_c6d4_core_073;
  wire popcount35_c6d4_core_074;
  wire popcount35_c6d4_core_075;
  wire popcount35_c6d4_core_076;
  wire popcount35_c6d4_core_077;
  wire popcount35_c6d4_core_078;
  wire popcount35_c6d4_core_079;
  wire popcount35_c6d4_core_080;
  wire popcount35_c6d4_core_082;
  wire popcount35_c6d4_core_083;
  wire popcount35_c6d4_core_085;
  wire popcount35_c6d4_core_090;
  wire popcount35_c6d4_core_091;
  wire popcount35_c6d4_core_092;
  wire popcount35_c6d4_core_093;
  wire popcount35_c6d4_core_100;
  wire popcount35_c6d4_core_103;
  wire popcount35_c6d4_core_104;
  wire popcount35_c6d4_core_108;
  wire popcount35_c6d4_core_109;
  wire popcount35_c6d4_core_112;
  wire popcount35_c6d4_core_113;
  wire popcount35_c6d4_core_115;
  wire popcount35_c6d4_core_116;
  wire popcount35_c6d4_core_117;
  wire popcount35_c6d4_core_118;
  wire popcount35_c6d4_core_119;
  wire popcount35_c6d4_core_120;
  wire popcount35_c6d4_core_121;
  wire popcount35_c6d4_core_122;
  wire popcount35_c6d4_core_123;
  wire popcount35_c6d4_core_124;
  wire popcount35_c6d4_core_125;
  wire popcount35_c6d4_core_126;
  wire popcount35_c6d4_core_127;
  wire popcount35_c6d4_core_128;
  wire popcount35_c6d4_core_129;
  wire popcount35_c6d4_core_130;
  wire popcount35_c6d4_core_131;
  wire popcount35_c6d4_core_132;
  wire popcount35_c6d4_core_133;
  wire popcount35_c6d4_core_134_not;
  wire popcount35_c6d4_core_135;
  wire popcount35_c6d4_core_136;
  wire popcount35_c6d4_core_137;
  wire popcount35_c6d4_core_138;
  wire popcount35_c6d4_core_139;
  wire popcount35_c6d4_core_140;
  wire popcount35_c6d4_core_141;
  wire popcount35_c6d4_core_142;
  wire popcount35_c6d4_core_143;
  wire popcount35_c6d4_core_145;
  wire popcount35_c6d4_core_146;
  wire popcount35_c6d4_core_147;
  wire popcount35_c6d4_core_148;
  wire popcount35_c6d4_core_149;
  wire popcount35_c6d4_core_150;
  wire popcount35_c6d4_core_151;
  wire popcount35_c6d4_core_152;
  wire popcount35_c6d4_core_155;
  wire popcount35_c6d4_core_156;
  wire popcount35_c6d4_core_158;
  wire popcount35_c6d4_core_159;
  wire popcount35_c6d4_core_161;
  wire popcount35_c6d4_core_162;
  wire popcount35_c6d4_core_163;
  wire popcount35_c6d4_core_164;
  wire popcount35_c6d4_core_165;
  wire popcount35_c6d4_core_166;
  wire popcount35_c6d4_core_167;
  wire popcount35_c6d4_core_168;
  wire popcount35_c6d4_core_169;
  wire popcount35_c6d4_core_170;
  wire popcount35_c6d4_core_171;
  wire popcount35_c6d4_core_172;
  wire popcount35_c6d4_core_173;
  wire popcount35_c6d4_core_174;
  wire popcount35_c6d4_core_175;
  wire popcount35_c6d4_core_177;
  wire popcount35_c6d4_core_178;
  wire popcount35_c6d4_core_179;
  wire popcount35_c6d4_core_181;
  wire popcount35_c6d4_core_182;
  wire popcount35_c6d4_core_183;
  wire popcount35_c6d4_core_184;
  wire popcount35_c6d4_core_185;
  wire popcount35_c6d4_core_186;
  wire popcount35_c6d4_core_188;
  wire popcount35_c6d4_core_189_not;
  wire popcount35_c6d4_core_191;
  wire popcount35_c6d4_core_192;
  wire popcount35_c6d4_core_193;
  wire popcount35_c6d4_core_194;
  wire popcount35_c6d4_core_196;
  wire popcount35_c6d4_core_197;
  wire popcount35_c6d4_core_198;
  wire popcount35_c6d4_core_199;
  wire popcount35_c6d4_core_200;
  wire popcount35_c6d4_core_201;
  wire popcount35_c6d4_core_203;
  wire popcount35_c6d4_core_209;
  wire popcount35_c6d4_core_210;
  wire popcount35_c6d4_core_211;
  wire popcount35_c6d4_core_212;
  wire popcount35_c6d4_core_213;
  wire popcount35_c6d4_core_214;
  wire popcount35_c6d4_core_215;
  wire popcount35_c6d4_core_216_not;
  wire popcount35_c6d4_core_218;
  wire popcount35_c6d4_core_220;
  wire popcount35_c6d4_core_221;
  wire popcount35_c6d4_core_223;
  wire popcount35_c6d4_core_224;
  wire popcount35_c6d4_core_225;
  wire popcount35_c6d4_core_226;
  wire popcount35_c6d4_core_227;
  wire popcount35_c6d4_core_228;
  wire popcount35_c6d4_core_229;
  wire popcount35_c6d4_core_230;
  wire popcount35_c6d4_core_231;
  wire popcount35_c6d4_core_232;
  wire popcount35_c6d4_core_233;
  wire popcount35_c6d4_core_235;
  wire popcount35_c6d4_core_236;
  wire popcount35_c6d4_core_238;
  wire popcount35_c6d4_core_239;
  wire popcount35_c6d4_core_240;
  wire popcount35_c6d4_core_241;
  wire popcount35_c6d4_core_242;
  wire popcount35_c6d4_core_243;
  wire popcount35_c6d4_core_244;
  wire popcount35_c6d4_core_245;
  wire popcount35_c6d4_core_246;
  wire popcount35_c6d4_core_247;
  wire popcount35_c6d4_core_248;
  wire popcount35_c6d4_core_249;
  wire popcount35_c6d4_core_250;
  wire popcount35_c6d4_core_251;
  wire popcount35_c6d4_core_252;
  wire popcount35_c6d4_core_253;
  wire popcount35_c6d4_core_254;
  wire popcount35_c6d4_core_255;
  wire popcount35_c6d4_core_256;
  wire popcount35_c6d4_core_257;
  wire popcount35_c6d4_core_258;
  wire popcount35_c6d4_core_259;
  wire popcount35_c6d4_core_260;
  wire popcount35_c6d4_core_262;
  wire popcount35_c6d4_core_263;

  assign popcount35_c6d4_core_037 = input_a[28] ^ input_a[1];
  assign popcount35_c6d4_core_039 = input_a[5] ^ input_a[3];
  assign popcount35_c6d4_core_043 = input_a[14] ^ input_a[16];
  assign popcount35_c6d4_core_045 = input_a[24] ^ input_a[30];
  assign popcount35_c6d4_core_046 = popcount35_c6d4_core_043 & input_a[18];
  assign popcount35_c6d4_core_047 = input_a[16] | input_a[5];
  assign popcount35_c6d4_core_048 = input_a[20] ^ input_a[5];
  assign popcount35_c6d4_core_050 = ~(input_a[6] | input_a[7]);
  assign popcount35_c6d4_core_051 = input_a[6] & input_a[7];
  assign popcount35_c6d4_core_052 = ~input_a[15];
  assign popcount35_c6d4_core_053 = popcount35_c6d4_core_048 & popcount35_c6d4_core_050;
  assign popcount35_c6d4_core_056 = popcount35_c6d4_core_051 ^ popcount35_c6d4_core_053;
  assign popcount35_c6d4_core_057 = popcount35_c6d4_core_051 & popcount35_c6d4_core_053;
  assign popcount35_c6d4_core_059_not = ~popcount35_c6d4_core_052;
  assign popcount35_c6d4_core_062 = popcount35_c6d4_core_045 & popcount35_c6d4_core_056;
  assign popcount35_c6d4_core_063 = input_a[23] ^ input_a[30];
  assign popcount35_c6d4_core_064 = input_a[3] & input_a[16];
  assign popcount35_c6d4_core_065 = popcount35_c6d4_core_062 | popcount35_c6d4_core_064;
  assign popcount35_c6d4_core_066 = ~(input_a[26] | popcount35_c6d4_core_057);
  assign popcount35_c6d4_core_067 = input_a[16] & popcount35_c6d4_core_057;
  assign popcount35_c6d4_core_068 = popcount35_c6d4_core_066 ^ popcount35_c6d4_core_065;
  assign popcount35_c6d4_core_069 = popcount35_c6d4_core_066 & popcount35_c6d4_core_065;
  assign popcount35_c6d4_core_070 = popcount35_c6d4_core_067 | popcount35_c6d4_core_069;
  assign popcount35_c6d4_core_071 = input_a[8] ^ input_a[9];
  assign popcount35_c6d4_core_072 = input_a[8] & input_a[9];
  assign popcount35_c6d4_core_073 = input_a[2] ^ input_a[14];
  assign popcount35_c6d4_core_074 = input_a[10] & input_a[12];
  assign popcount35_c6d4_core_075 = popcount35_c6d4_core_071 ^ input_a[9];
  assign popcount35_c6d4_core_076 = popcount35_c6d4_core_071 & input_a[32];
  assign popcount35_c6d4_core_077 = popcount35_c6d4_core_072 ^ popcount35_c6d4_core_074;
  assign popcount35_c6d4_core_078 = popcount35_c6d4_core_072 & popcount35_c6d4_core_074;
  assign popcount35_c6d4_core_079 = popcount35_c6d4_core_077 ^ popcount35_c6d4_core_076;
  assign popcount35_c6d4_core_080 = popcount35_c6d4_core_077 & popcount35_c6d4_core_076;
  assign popcount35_c6d4_core_082 = input_a[21] & input_a[13];
  assign popcount35_c6d4_core_083 = ~input_a[12];
  assign popcount35_c6d4_core_085 = input_a[15] & input_a[16];
  assign popcount35_c6d4_core_090 = input_a[24] ^ input_a[13];
  assign popcount35_c6d4_core_091 = popcount35_c6d4_core_082 & input_a[10];
  assign popcount35_c6d4_core_092 = input_a[8] ^ input_a[12];
  assign popcount35_c6d4_core_093 = popcount35_c6d4_core_083 & input_a[2];
  assign popcount35_c6d4_core_100 = popcount35_c6d4_core_075 & popcount35_c6d4_core_090;
  assign popcount35_c6d4_core_103 = popcount35_c6d4_core_079 ^ popcount35_c6d4_core_100;
  assign popcount35_c6d4_core_104 = popcount35_c6d4_core_079 & popcount35_c6d4_core_100;
  assign popcount35_c6d4_core_108 = popcount35_c6d4_core_078 ^ popcount35_c6d4_core_104;
  assign popcount35_c6d4_core_109 = popcount35_c6d4_core_078 & popcount35_c6d4_core_104;
  assign popcount35_c6d4_core_112 = input_a[30] & popcount35_c6d4_core_109;
  assign popcount35_c6d4_core_113 = popcount35_c6d4_core_059_not ^ popcount35_c6d4_core_075;
  assign popcount35_c6d4_core_115 = popcount35_c6d4_core_063 ^ popcount35_c6d4_core_103;
  assign popcount35_c6d4_core_116 = popcount35_c6d4_core_063 & popcount35_c6d4_core_103;
  assign popcount35_c6d4_core_117 = popcount35_c6d4_core_115 ^ input_a[19];
  assign popcount35_c6d4_core_118 = popcount35_c6d4_core_115 & input_a[19];
  assign popcount35_c6d4_core_119 = popcount35_c6d4_core_116 | popcount35_c6d4_core_118;
  assign popcount35_c6d4_core_120 = popcount35_c6d4_core_068 ^ popcount35_c6d4_core_108;
  assign popcount35_c6d4_core_121 = popcount35_c6d4_core_068 & popcount35_c6d4_core_108;
  assign popcount35_c6d4_core_122 = popcount35_c6d4_core_120 ^ popcount35_c6d4_core_119;
  assign popcount35_c6d4_core_123 = popcount35_c6d4_core_120 & popcount35_c6d4_core_119;
  assign popcount35_c6d4_core_124 = popcount35_c6d4_core_121 | popcount35_c6d4_core_123;
  assign popcount35_c6d4_core_125 = popcount35_c6d4_core_070 ^ popcount35_c6d4_core_109;
  assign popcount35_c6d4_core_126 = input_a[0] & popcount35_c6d4_core_109;
  assign popcount35_c6d4_core_127 = popcount35_c6d4_core_125 ^ popcount35_c6d4_core_124;
  assign popcount35_c6d4_core_128 = popcount35_c6d4_core_125 & popcount35_c6d4_core_124;
  assign popcount35_c6d4_core_129 = popcount35_c6d4_core_126 | popcount35_c6d4_core_128;
  assign popcount35_c6d4_core_130 = popcount35_c6d4_core_112 ^ popcount35_c6d4_core_129;
  assign popcount35_c6d4_core_131 = popcount35_c6d4_core_112 & input_a[15];
  assign popcount35_c6d4_core_132 = input_a[25] ^ input_a[18];
  assign popcount35_c6d4_core_133 = input_a[2] & input_a[18];
  assign popcount35_c6d4_core_134_not = ~input_a[20];
  assign popcount35_c6d4_core_135 = input_a[15] & input_a[20];
  assign popcount35_c6d4_core_136 = popcount35_c6d4_core_132 ^ input_a[16];
  assign popcount35_c6d4_core_137 = input_a[5] & popcount35_c6d4_core_134_not;
  assign popcount35_c6d4_core_138 = popcount35_c6d4_core_133 ^ popcount35_c6d4_core_135;
  assign popcount35_c6d4_core_139 = popcount35_c6d4_core_133 & popcount35_c6d4_core_135;
  assign popcount35_c6d4_core_140 = popcount35_c6d4_core_138 ^ popcount35_c6d4_core_137;
  assign popcount35_c6d4_core_141 = popcount35_c6d4_core_138 & popcount35_c6d4_core_137;
  assign popcount35_c6d4_core_142 = popcount35_c6d4_core_139 | popcount35_c6d4_core_141;
  assign popcount35_c6d4_core_143 = ~(input_a[21] & input_a[0]);
  assign popcount35_c6d4_core_145 = input_a[24] ^ input_a[2];
  assign popcount35_c6d4_core_146 = input_a[14] & input_a[25];
  assign popcount35_c6d4_core_147 = ~(input_a[23] & popcount35_c6d4_core_145);
  assign popcount35_c6d4_core_148 = input_a[23] & popcount35_c6d4_core_145;
  assign popcount35_c6d4_core_149 = popcount35_c6d4_core_146 ^ popcount35_c6d4_core_148;
  assign popcount35_c6d4_core_150 = popcount35_c6d4_core_146 & popcount35_c6d4_core_148;
  assign popcount35_c6d4_core_151 = popcount35_c6d4_core_143 ^ popcount35_c6d4_core_147;
  assign popcount35_c6d4_core_152 = popcount35_c6d4_core_143 & popcount35_c6d4_core_147;
  assign popcount35_c6d4_core_155 = popcount35_c6d4_core_149 ^ popcount35_c6d4_core_152;
  assign popcount35_c6d4_core_156 = popcount35_c6d4_core_149 & popcount35_c6d4_core_152;
  assign popcount35_c6d4_core_158 = popcount35_c6d4_core_150 ^ popcount35_c6d4_core_156;
  assign popcount35_c6d4_core_159 = popcount35_c6d4_core_150 & popcount35_c6d4_core_156;
  assign popcount35_c6d4_core_161 = input_a[30] & popcount35_c6d4_core_151;
  assign popcount35_c6d4_core_162 = popcount35_c6d4_core_140 ^ popcount35_c6d4_core_155;
  assign popcount35_c6d4_core_163 = popcount35_c6d4_core_140 & popcount35_c6d4_core_155;
  assign popcount35_c6d4_core_164 = popcount35_c6d4_core_162 ^ popcount35_c6d4_core_161;
  assign popcount35_c6d4_core_165 = input_a[27] & popcount35_c6d4_core_161;
  assign popcount35_c6d4_core_166 = popcount35_c6d4_core_163 | popcount35_c6d4_core_165;
  assign popcount35_c6d4_core_167 = popcount35_c6d4_core_142 ^ popcount35_c6d4_core_158;
  assign popcount35_c6d4_core_168 = popcount35_c6d4_core_142 & popcount35_c6d4_core_158;
  assign popcount35_c6d4_core_169 = popcount35_c6d4_core_167 ^ popcount35_c6d4_core_166;
  assign popcount35_c6d4_core_170 = popcount35_c6d4_core_167 & popcount35_c6d4_core_166;
  assign popcount35_c6d4_core_171 = ~popcount35_c6d4_core_168;
  assign popcount35_c6d4_core_172 = popcount35_c6d4_core_159 & popcount35_c6d4_core_171;
  assign popcount35_c6d4_core_173 = popcount35_c6d4_core_159 & popcount35_c6d4_core_171;
  assign popcount35_c6d4_core_174 = input_a[26] ^ input_a[13];
  assign popcount35_c6d4_core_175 = input_a[26] & input_a[27];
  assign popcount35_c6d4_core_177 = ~(input_a[28] ^ input_a[23]);
  assign popcount35_c6d4_core_178 = popcount35_c6d4_core_174 ^ input_a[3];
  assign popcount35_c6d4_core_179 = input_a[14] & input_a[3];
  assign popcount35_c6d4_core_181 = popcount35_c6d4_core_175 & input_a[26];
  assign popcount35_c6d4_core_182 = input_a[22] & input_a[22];
  assign popcount35_c6d4_core_183 = input_a[22] & popcount35_c6d4_core_179;
  assign popcount35_c6d4_core_184 = popcount35_c6d4_core_181 | popcount35_c6d4_core_183;
  assign popcount35_c6d4_core_185 = ~input_a[19];
  assign popcount35_c6d4_core_186 = input_a[12] & input_a[4];
  assign popcount35_c6d4_core_188 = input_a[33] & input_a[34];
  assign popcount35_c6d4_core_189_not = ~input_a[32];
  assign popcount35_c6d4_core_191 = popcount35_c6d4_core_188 ^ input_a[32];
  assign popcount35_c6d4_core_192 = popcount35_c6d4_core_188 & input_a[32];
  assign popcount35_c6d4_core_193 = popcount35_c6d4_core_185 ^ popcount35_c6d4_core_189_not;
  assign popcount35_c6d4_core_194 = input_a[9] & popcount35_c6d4_core_189_not;
  assign popcount35_c6d4_core_196 = popcount35_c6d4_core_186 & popcount35_c6d4_core_191;
  assign popcount35_c6d4_core_197 = popcount35_c6d4_core_186 ^ popcount35_c6d4_core_194;
  assign popcount35_c6d4_core_198 = popcount35_c6d4_core_186 & popcount35_c6d4_core_194;
  assign popcount35_c6d4_core_199 = popcount35_c6d4_core_196 | popcount35_c6d4_core_198;
  assign popcount35_c6d4_core_200 = popcount35_c6d4_core_192 ^ popcount35_c6d4_core_199;
  assign popcount35_c6d4_core_201 = popcount35_c6d4_core_192 & popcount35_c6d4_core_199;
  assign popcount35_c6d4_core_203 = ~popcount35_c6d4_core_178;
  assign popcount35_c6d4_core_209 = popcount35_c6d4_core_184 ^ popcount35_c6d4_core_200;
  assign popcount35_c6d4_core_210 = popcount35_c6d4_core_184 & popcount35_c6d4_core_200;
  assign popcount35_c6d4_core_211 = popcount35_c6d4_core_209 ^ input_a[26];
  assign popcount35_c6d4_core_212 = popcount35_c6d4_core_209 & input_a[26];
  assign popcount35_c6d4_core_213 = popcount35_c6d4_core_210 | popcount35_c6d4_core_212;
  assign popcount35_c6d4_core_214 = popcount35_c6d4_core_201 ^ popcount35_c6d4_core_213;
  assign popcount35_c6d4_core_215 = popcount35_c6d4_core_201 & popcount35_c6d4_core_213;
  assign popcount35_c6d4_core_216_not = ~input_a[20];
  assign popcount35_c6d4_core_218 = input_a[0] ^ input_a[17];
  assign popcount35_c6d4_core_220 = popcount35_c6d4_core_218 ^ input_a[20];
  assign popcount35_c6d4_core_221 = popcount35_c6d4_core_218 & input_a[20];
  assign popcount35_c6d4_core_223 = popcount35_c6d4_core_169 ^ popcount35_c6d4_core_211;
  assign popcount35_c6d4_core_224 = popcount35_c6d4_core_169 & popcount35_c6d4_core_211;
  assign popcount35_c6d4_core_225 = popcount35_c6d4_core_223 ^ popcount35_c6d4_core_221;
  assign popcount35_c6d4_core_226 = popcount35_c6d4_core_223 & popcount35_c6d4_core_221;
  assign popcount35_c6d4_core_227 = popcount35_c6d4_core_224 | popcount35_c6d4_core_226;
  assign popcount35_c6d4_core_228 = popcount35_c6d4_core_172 ^ popcount35_c6d4_core_214;
  assign popcount35_c6d4_core_229 = popcount35_c6d4_core_172 & popcount35_c6d4_core_214;
  assign popcount35_c6d4_core_230 = popcount35_c6d4_core_228 ^ popcount35_c6d4_core_227;
  assign popcount35_c6d4_core_231 = popcount35_c6d4_core_228 & popcount35_c6d4_core_227;
  assign popcount35_c6d4_core_232 = popcount35_c6d4_core_229 | popcount35_c6d4_core_231;
  assign popcount35_c6d4_core_233 = popcount35_c6d4_core_173 ^ popcount35_c6d4_core_215;
  assign popcount35_c6d4_core_235 = popcount35_c6d4_core_233 ^ popcount35_c6d4_core_232;
  assign popcount35_c6d4_core_236 = popcount35_c6d4_core_233 & popcount35_c6d4_core_232;
  assign popcount35_c6d4_core_238 = popcount35_c6d4_core_113 ^ popcount35_c6d4_core_216_not;
  assign popcount35_c6d4_core_239 = input_a[17] & popcount35_c6d4_core_216_not;
  assign popcount35_c6d4_core_240 = popcount35_c6d4_core_117 ^ popcount35_c6d4_core_220;
  assign popcount35_c6d4_core_241 = popcount35_c6d4_core_117 & popcount35_c6d4_core_220;
  assign popcount35_c6d4_core_242 = popcount35_c6d4_core_240 ^ popcount35_c6d4_core_239;
  assign popcount35_c6d4_core_243 = popcount35_c6d4_core_240 & popcount35_c6d4_core_239;
  assign popcount35_c6d4_core_244 = popcount35_c6d4_core_241 | popcount35_c6d4_core_243;
  assign popcount35_c6d4_core_245 = popcount35_c6d4_core_122 ^ popcount35_c6d4_core_225;
  assign popcount35_c6d4_core_246 = popcount35_c6d4_core_122 & popcount35_c6d4_core_225;
  assign popcount35_c6d4_core_247 = popcount35_c6d4_core_245 ^ popcount35_c6d4_core_244;
  assign popcount35_c6d4_core_248 = popcount35_c6d4_core_245 & popcount35_c6d4_core_244;
  assign popcount35_c6d4_core_249 = popcount35_c6d4_core_246 | popcount35_c6d4_core_248;
  assign popcount35_c6d4_core_250 = popcount35_c6d4_core_127 ^ popcount35_c6d4_core_230;
  assign popcount35_c6d4_core_251 = popcount35_c6d4_core_127 & popcount35_c6d4_core_230;
  assign popcount35_c6d4_core_252 = popcount35_c6d4_core_250 ^ popcount35_c6d4_core_249;
  assign popcount35_c6d4_core_253 = popcount35_c6d4_core_250 & popcount35_c6d4_core_249;
  assign popcount35_c6d4_core_254 = popcount35_c6d4_core_251 | popcount35_c6d4_core_253;
  assign popcount35_c6d4_core_255 = popcount35_c6d4_core_130 ^ popcount35_c6d4_core_235;
  assign popcount35_c6d4_core_256 = popcount35_c6d4_core_130 & popcount35_c6d4_core_235;
  assign popcount35_c6d4_core_257 = popcount35_c6d4_core_255 ^ popcount35_c6d4_core_254;
  assign popcount35_c6d4_core_258 = popcount35_c6d4_core_255 & popcount35_c6d4_core_254;
  assign popcount35_c6d4_core_259 = popcount35_c6d4_core_256 | popcount35_c6d4_core_258;
  assign popcount35_c6d4_core_260 = popcount35_c6d4_core_131 ^ popcount35_c6d4_core_236;
  assign popcount35_c6d4_core_262 = popcount35_c6d4_core_260 ^ popcount35_c6d4_core_259;
  assign popcount35_c6d4_core_263 = popcount35_c6d4_core_260 & input_a[27];

  assign popcount35_c6d4_out[0] = popcount35_c6d4_core_197;
  assign popcount35_c6d4_out[1] = popcount35_c6d4_core_242;
  assign popcount35_c6d4_out[2] = popcount35_c6d4_core_247;
  assign popcount35_c6d4_out[3] = popcount35_c6d4_core_252;
  assign popcount35_c6d4_out[4] = popcount35_c6d4_core_257;
  assign popcount35_c6d4_out[5] = popcount35_c6d4_core_262;
endmodule