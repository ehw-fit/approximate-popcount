// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.5492
// WCE=49.0
// EP=0.960076%
// Printed PDK parameters:
//  Area=70587676.0
//  Delay=70281536.0
//  Power=2980000.0

module popcount39_35p6(input [38:0] input_a, output [5:0] popcount39_35p6_out);
  wire popcount39_35p6_core_041;
  wire popcount39_35p6_core_042;
  wire popcount39_35p6_core_043;
  wire popcount39_35p6_core_044;
  wire popcount39_35p6_core_047;
  wire popcount39_35p6_core_048;
  wire popcount39_35p6_core_049_not;
  wire popcount39_35p6_core_052;
  wire popcount39_35p6_core_054;
  wire popcount39_35p6_core_055;
  wire popcount39_35p6_core_057;
  wire popcount39_35p6_core_058;
  wire popcount39_35p6_core_059;
  wire popcount39_35p6_core_071;
  wire popcount39_35p6_core_072;
  wire popcount39_35p6_core_073;
  wire popcount39_35p6_core_076;
  wire popcount39_35p6_core_077;
  wire popcount39_35p6_core_078;
  wire popcount39_35p6_core_084;
  wire popcount39_35p6_core_085;
  wire popcount39_35p6_core_086;
  wire popcount39_35p6_core_087;
  wire popcount39_35p6_core_088;
  wire popcount39_35p6_core_089;
  wire popcount39_35p6_core_090;
  wire popcount39_35p6_core_093;
  wire popcount39_35p6_core_094;
  wire popcount39_35p6_core_098;
  wire popcount39_35p6_core_099;
  wire popcount39_35p6_core_100;
  wire popcount39_35p6_core_101;
  wire popcount39_35p6_core_102;
  wire popcount39_35p6_core_103;
  wire popcount39_35p6_core_104;
  wire popcount39_35p6_core_105;
  wire popcount39_35p6_core_106;
  wire popcount39_35p6_core_107;
  wire popcount39_35p6_core_108;
  wire popcount39_35p6_core_109;
  wire popcount39_35p6_core_110;
  wire popcount39_35p6_core_111;
  wire popcount39_35p6_core_112;
  wire popcount39_35p6_core_113;
  wire popcount39_35p6_core_114;
  wire popcount39_35p6_core_115;
  wire popcount39_35p6_core_116;
  wire popcount39_35p6_core_117;
  wire popcount39_35p6_core_118;
  wire popcount39_35p6_core_120;
  wire popcount39_35p6_core_123;
  wire popcount39_35p6_core_124;
  wire popcount39_35p6_core_125;
  wire popcount39_35p6_core_126;
  wire popcount39_35p6_core_127;
  wire popcount39_35p6_core_128;
  wire popcount39_35p6_core_129;
  wire popcount39_35p6_core_130;
  wire popcount39_35p6_core_131;
  wire popcount39_35p6_core_132;
  wire popcount39_35p6_core_133;
  wire popcount39_35p6_core_136;
  wire popcount39_35p6_core_137;
  wire popcount39_35p6_core_141;
  wire popcount39_35p6_core_142;
  wire popcount39_35p6_core_143;
  wire popcount39_35p6_core_144;
  wire popcount39_35p6_core_145;
  wire popcount39_35p6_core_146;
  wire popcount39_35p6_core_147;
  wire popcount39_35p6_core_148;
  wire popcount39_35p6_core_149;
  wire popcount39_35p6_core_150;
  wire popcount39_35p6_core_156;
  wire popcount39_35p6_core_157;
  wire popcount39_35p6_core_158;
  wire popcount39_35p6_core_159;
  wire popcount39_35p6_core_160;
  wire popcount39_35p6_core_161;
  wire popcount39_35p6_core_162;
  wire popcount39_35p6_core_163;
  wire popcount39_35p6_core_164;
  wire popcount39_35p6_core_165;
  wire popcount39_35p6_core_166;
  wire popcount39_35p6_core_167;
  wire popcount39_35p6_core_168;
  wire popcount39_35p6_core_169;
  wire popcount39_35p6_core_170;
  wire popcount39_35p6_core_171;
  wire popcount39_35p6_core_172;
  wire popcount39_35p6_core_173;
  wire popcount39_35p6_core_174;
  wire popcount39_35p6_core_175;
  wire popcount39_35p6_core_176;
  wire popcount39_35p6_core_177;
  wire popcount39_35p6_core_178;
  wire popcount39_35p6_core_179;
  wire popcount39_35p6_core_180;
  wire popcount39_35p6_core_181;
  wire popcount39_35p6_core_183;
  wire popcount39_35p6_core_184;
  wire popcount39_35p6_core_185;
  wire popcount39_35p6_core_190;
  wire popcount39_35p6_core_192;
  wire popcount39_35p6_core_193;
  wire popcount39_35p6_core_197;
  wire popcount39_35p6_core_198;
  wire popcount39_35p6_core_199;
  wire popcount39_35p6_core_200;
  wire popcount39_35p6_core_201;
  wire popcount39_35p6_core_203;
  wire popcount39_35p6_core_204;
  wire popcount39_35p6_core_205;
  wire popcount39_35p6_core_207;
  wire popcount39_35p6_core_208;
  wire popcount39_35p6_core_209;
  wire popcount39_35p6_core_210;
  wire popcount39_35p6_core_211;
  wire popcount39_35p6_core_212;
  wire popcount39_35p6_core_213;
  wire popcount39_35p6_core_214;
  wire popcount39_35p6_core_215;
  wire popcount39_35p6_core_216;
  wire popcount39_35p6_core_217;
  wire popcount39_35p6_core_218;
  wire popcount39_35p6_core_219;
  wire popcount39_35p6_core_220;
  wire popcount39_35p6_core_221;
  wire popcount39_35p6_core_222;
  wire popcount39_35p6_core_223;
  wire popcount39_35p6_core_225;
  wire popcount39_35p6_core_226;
  wire popcount39_35p6_core_227;
  wire popcount39_35p6_core_228;
  wire popcount39_35p6_core_229;
  wire popcount39_35p6_core_230;
  wire popcount39_35p6_core_231;
  wire popcount39_35p6_core_232;
  wire popcount39_35p6_core_233;
  wire popcount39_35p6_core_234;
  wire popcount39_35p6_core_235;
  wire popcount39_35p6_core_236;
  wire popcount39_35p6_core_237;
  wire popcount39_35p6_core_238;
  wire popcount39_35p6_core_239;
  wire popcount39_35p6_core_240;
  wire popcount39_35p6_core_241;
  wire popcount39_35p6_core_242;
  wire popcount39_35p6_core_243;
  wire popcount39_35p6_core_244;
  wire popcount39_35p6_core_245;
  wire popcount39_35p6_core_246;
  wire popcount39_35p6_core_247;
  wire popcount39_35p6_core_248;
  wire popcount39_35p6_core_249;
  wire popcount39_35p6_core_250;
  wire popcount39_35p6_core_251;
  wire popcount39_35p6_core_252;
  wire popcount39_35p6_core_253;
  wire popcount39_35p6_core_254;
  wire popcount39_35p6_core_255;
  wire popcount39_35p6_core_256;
  wire popcount39_35p6_core_257;
  wire popcount39_35p6_core_258;
  wire popcount39_35p6_core_259;
  wire popcount39_35p6_core_260;
  wire popcount39_35p6_core_261;
  wire popcount39_35p6_core_262;
  wire popcount39_35p6_core_263;
  wire popcount39_35p6_core_264;
  wire popcount39_35p6_core_265;
  wire popcount39_35p6_core_266;
  wire popcount39_35p6_core_267;
  wire popcount39_35p6_core_268;
  wire popcount39_35p6_core_269;
  wire popcount39_35p6_core_270;
  wire popcount39_35p6_core_271;
  wire popcount39_35p6_core_272;
  wire popcount39_35p6_core_273;
  wire popcount39_35p6_core_274;
  wire popcount39_35p6_core_282;
  wire popcount39_35p6_core_283;
  wire popcount39_35p6_core_287;
  wire popcount39_35p6_core_288;
  wire popcount39_35p6_core_290;
  wire popcount39_35p6_core_291;
  wire popcount39_35p6_core_292;
  wire popcount39_35p6_core_293;
  wire popcount39_35p6_core_294;
  wire popcount39_35p6_core_295;
  wire popcount39_35p6_core_296;
  wire popcount39_35p6_core_297;
  wire popcount39_35p6_core_298;
  wire popcount39_35p6_core_299;
  wire popcount39_35p6_core_300;
  wire popcount39_35p6_core_301;

  assign popcount39_35p6_core_041 = input_a[0] ^ input_a[1];
  assign popcount39_35p6_core_042 = input_a[0] & input_a[1];
  assign popcount39_35p6_core_043 = input_a[2] ^ input_a[3];
  assign popcount39_35p6_core_044 = input_a[2] & input_a[3];
  assign popcount39_35p6_core_047 = popcount39_35p6_core_042 ^ input_a[38];
  assign popcount39_35p6_core_048 = popcount39_35p6_core_042 & popcount39_35p6_core_044;
  assign popcount39_35p6_core_049_not = ~popcount39_35p6_core_047;
  assign popcount39_35p6_core_052 = input_a[4] ^ input_a[5];
  assign popcount39_35p6_core_054 = input_a[7] ^ input_a[8];
  assign popcount39_35p6_core_055 = input_a[7] & input_a[8];
  assign popcount39_35p6_core_057 = input_a[6] & input_a[37];
  assign popcount39_35p6_core_058 = popcount39_35p6_core_055 ^ input_a[23];
  assign popcount39_35p6_core_059 = popcount39_35p6_core_055 & popcount39_35p6_core_057;
  assign popcount39_35p6_core_071 = ~popcount39_35p6_core_049_not;
  assign popcount39_35p6_core_072 = popcount39_35p6_core_049_not & input_a[12];
  assign popcount39_35p6_core_073 = popcount39_35p6_core_071 ^ input_a[38];
  assign popcount39_35p6_core_076 = ~(popcount39_35p6_core_048 | popcount39_35p6_core_059);
  assign popcount39_35p6_core_077 = popcount39_35p6_core_048 & popcount39_35p6_core_059;
  assign popcount39_35p6_core_078 = popcount39_35p6_core_076 ^ input_a[21];
  assign popcount39_35p6_core_084 = input_a[9] & input_a[10];
  assign popcount39_35p6_core_085 = input_a[12] ^ input_a[13];
  assign popcount39_35p6_core_086 = input_a[12] & input_a[13];
  assign popcount39_35p6_core_087 = input_a[11] ^ popcount39_35p6_core_085;
  assign popcount39_35p6_core_088 = input_a[22] & popcount39_35p6_core_085;
  assign popcount39_35p6_core_089 = popcount39_35p6_core_086 ^ popcount39_35p6_core_088;
  assign popcount39_35p6_core_090 = popcount39_35p6_core_086 & popcount39_35p6_core_088;
  assign popcount39_35p6_core_093 = popcount39_35p6_core_084 ^ popcount39_35p6_core_089;
  assign popcount39_35p6_core_094 = popcount39_35p6_core_084 & input_a[25];
  assign popcount39_35p6_core_098 = ~(popcount39_35p6_core_090 & popcount39_35p6_core_094);
  assign popcount39_35p6_core_099 = popcount39_35p6_core_090 & popcount39_35p6_core_094;
  assign popcount39_35p6_core_100 = input_a[14] ^ input_a[15];
  assign popcount39_35p6_core_101 = input_a[14] & input_a[15];
  assign popcount39_35p6_core_102 = input_a[17] ^ input_a[18];
  assign popcount39_35p6_core_103 = input_a[17] & input_a[18];
  assign popcount39_35p6_core_104 = input_a[0] | popcount39_35p6_core_102;
  assign popcount39_35p6_core_105 = input_a[16] & popcount39_35p6_core_102;
  assign popcount39_35p6_core_106 = popcount39_35p6_core_103 ^ input_a[10];
  assign popcount39_35p6_core_107 = popcount39_35p6_core_103 & popcount39_35p6_core_105;
  assign popcount39_35p6_core_108 = popcount39_35p6_core_100 ^ popcount39_35p6_core_104;
  assign popcount39_35p6_core_109 = popcount39_35p6_core_100 & input_a[24];
  assign popcount39_35p6_core_110 = input_a[38] ^ popcount39_35p6_core_106;
  assign popcount39_35p6_core_111 = popcount39_35p6_core_101 & popcount39_35p6_core_106;
  assign popcount39_35p6_core_112 = input_a[15] ^ popcount39_35p6_core_109;
  assign popcount39_35p6_core_113 = popcount39_35p6_core_110 & popcount39_35p6_core_109;
  assign popcount39_35p6_core_114 = input_a[5] | input_a[5];
  assign popcount39_35p6_core_115 = popcount39_35p6_core_107 ^ popcount39_35p6_core_114;
  assign popcount39_35p6_core_116 = popcount39_35p6_core_107 & popcount39_35p6_core_114;
  assign popcount39_35p6_core_117 = input_a[4] ^ popcount39_35p6_core_108;
  assign popcount39_35p6_core_118 = input_a[33] & popcount39_35p6_core_108;
  assign popcount39_35p6_core_120 = popcount39_35p6_core_093 & popcount39_35p6_core_112;
  assign popcount39_35p6_core_123 = popcount39_35p6_core_120 | input_a[27];
  assign popcount39_35p6_core_124 = popcount39_35p6_core_098 ^ popcount39_35p6_core_115;
  assign popcount39_35p6_core_125 = popcount39_35p6_core_098 & popcount39_35p6_core_115;
  assign popcount39_35p6_core_126 = popcount39_35p6_core_124 ^ popcount39_35p6_core_123;
  assign popcount39_35p6_core_127 = popcount39_35p6_core_124 & popcount39_35p6_core_123;
  assign popcount39_35p6_core_128 = input_a[21] | popcount39_35p6_core_127;
  assign popcount39_35p6_core_129 = popcount39_35p6_core_099 ^ input_a[26];
  assign popcount39_35p6_core_130 = popcount39_35p6_core_099 & popcount39_35p6_core_116;
  assign popcount39_35p6_core_131 = input_a[1] ^ popcount39_35p6_core_128;
  assign popcount39_35p6_core_132 = popcount39_35p6_core_129 & input_a[35];
  assign popcount39_35p6_core_133 = popcount39_35p6_core_130 | popcount39_35p6_core_132;
  assign popcount39_35p6_core_136 = popcount39_35p6_core_073 ^ popcount39_35p6_core_118;
  assign popcount39_35p6_core_137 = popcount39_35p6_core_073 & popcount39_35p6_core_118;
  assign popcount39_35p6_core_141 = input_a[2] ^ popcount39_35p6_core_126;
  assign popcount39_35p6_core_142 = input_a[10] & popcount39_35p6_core_126;
  assign popcount39_35p6_core_143 = popcount39_35p6_core_141 ^ popcount39_35p6_core_137;
  assign popcount39_35p6_core_144 = popcount39_35p6_core_141 & popcount39_35p6_core_137;
  assign popcount39_35p6_core_145 = popcount39_35p6_core_142 | popcount39_35p6_core_144;
  assign popcount39_35p6_core_146 = popcount39_35p6_core_077 ^ popcount39_35p6_core_131;
  assign popcount39_35p6_core_147 = popcount39_35p6_core_077 & popcount39_35p6_core_131;
  assign popcount39_35p6_core_148 = popcount39_35p6_core_146 ^ popcount39_35p6_core_145;
  assign popcount39_35p6_core_149 = popcount39_35p6_core_146 & popcount39_35p6_core_145;
  assign popcount39_35p6_core_150 = popcount39_35p6_core_147 | popcount39_35p6_core_149;
  assign popcount39_35p6_core_156 = input_a[19] ^ input_a[20];
  assign popcount39_35p6_core_157 = input_a[19] & input_a[20];
  assign popcount39_35p6_core_158 = input_a[22] ^ input_a[20];
  assign popcount39_35p6_core_159 = input_a[22] & input_a[23];
  assign popcount39_35p6_core_160 = input_a[21] ^ popcount39_35p6_core_158;
  assign popcount39_35p6_core_161 = input_a[21] & popcount39_35p6_core_158;
  assign popcount39_35p6_core_162 = popcount39_35p6_core_159 ^ popcount39_35p6_core_161;
  assign popcount39_35p6_core_163 = popcount39_35p6_core_159 & popcount39_35p6_core_161;
  assign popcount39_35p6_core_164 = input_a[38] ^ popcount39_35p6_core_160;
  assign popcount39_35p6_core_165 = popcount39_35p6_core_156 & popcount39_35p6_core_160;
  assign popcount39_35p6_core_166 = popcount39_35p6_core_157 ^ popcount39_35p6_core_162;
  assign popcount39_35p6_core_167 = popcount39_35p6_core_157 & popcount39_35p6_core_162;
  assign popcount39_35p6_core_168 = popcount39_35p6_core_166 ^ input_a[22];
  assign popcount39_35p6_core_169 = popcount39_35p6_core_166 & popcount39_35p6_core_165;
  assign popcount39_35p6_core_170 = popcount39_35p6_core_167 | input_a[3];
  assign popcount39_35p6_core_171 = popcount39_35p6_core_163 ^ popcount39_35p6_core_170;
  assign popcount39_35p6_core_172 = popcount39_35p6_core_163 & popcount39_35p6_core_170;
  assign popcount39_35p6_core_173 = input_a[24] ^ input_a[25];
  assign popcount39_35p6_core_174 = input_a[24] & input_a[25];
  assign popcount39_35p6_core_175 = input_a[27] ^ input_a[28];
  assign popcount39_35p6_core_176 = input_a[27] & input_a[28];
  assign popcount39_35p6_core_177 = ~(input_a[26] & popcount39_35p6_core_175);
  assign popcount39_35p6_core_178 = input_a[26] & popcount39_35p6_core_175;
  assign popcount39_35p6_core_179 = ~popcount39_35p6_core_176;
  assign popcount39_35p6_core_180 = popcount39_35p6_core_176 & popcount39_35p6_core_178;
  assign popcount39_35p6_core_181 = input_a[22] & popcount39_35p6_core_177;
  assign popcount39_35p6_core_183 = popcount39_35p6_core_174 ^ popcount39_35p6_core_179;
  assign popcount39_35p6_core_184 = popcount39_35p6_core_174 & popcount39_35p6_core_179;
  assign popcount39_35p6_core_185 = ~popcount39_35p6_core_183;
  assign popcount39_35p6_core_190 = input_a[4] | popcount39_35p6_core_181;
  assign popcount39_35p6_core_192 = popcount39_35p6_core_168 ^ popcount39_35p6_core_185;
  assign popcount39_35p6_core_193 = popcount39_35p6_core_168 & popcount39_35p6_core_185;
  assign popcount39_35p6_core_197 = popcount39_35p6_core_171 ^ input_a[24];
  assign popcount39_35p6_core_198 = popcount39_35p6_core_171 & input_a[24];
  assign popcount39_35p6_core_199 = popcount39_35p6_core_197 ^ popcount39_35p6_core_193;
  assign popcount39_35p6_core_200 = popcount39_35p6_core_197 & popcount39_35p6_core_193;
  assign popcount39_35p6_core_201 = popcount39_35p6_core_198 | input_a[14];
  assign popcount39_35p6_core_203 = popcount39_35p6_core_172 & input_a[17];
  assign popcount39_35p6_core_204 = input_a[10] ^ popcount39_35p6_core_201;
  assign popcount39_35p6_core_205 = input_a[10] & input_a[14];
  assign popcount39_35p6_core_207 = input_a[29] ^ input_a[30];
  assign popcount39_35p6_core_208 = input_a[29] & input_a[30];
  assign popcount39_35p6_core_209 = input_a[32] ^ input_a[6];
  assign popcount39_35p6_core_210 = input_a[32] & input_a[33];
  assign popcount39_35p6_core_211 = input_a[10] ^ popcount39_35p6_core_209;
  assign popcount39_35p6_core_212 = input_a[31] & popcount39_35p6_core_209;
  assign popcount39_35p6_core_213 = popcount39_35p6_core_210 ^ popcount39_35p6_core_212;
  assign popcount39_35p6_core_214 = popcount39_35p6_core_210 & popcount39_35p6_core_212;
  assign popcount39_35p6_core_215 = popcount39_35p6_core_207 ^ popcount39_35p6_core_211;
  assign popcount39_35p6_core_216 = popcount39_35p6_core_207 & popcount39_35p6_core_211;
  assign popcount39_35p6_core_217 = popcount39_35p6_core_208 ^ popcount39_35p6_core_213;
  assign popcount39_35p6_core_218 = input_a[37] & popcount39_35p6_core_213;
  assign popcount39_35p6_core_219 = popcount39_35p6_core_217 ^ popcount39_35p6_core_216;
  assign popcount39_35p6_core_220 = popcount39_35p6_core_217 & popcount39_35p6_core_216;
  assign popcount39_35p6_core_221 = popcount39_35p6_core_218 | popcount39_35p6_core_220;
  assign popcount39_35p6_core_222 = popcount39_35p6_core_214 ^ popcount39_35p6_core_221;
  assign popcount39_35p6_core_223 = popcount39_35p6_core_214 & popcount39_35p6_core_221;
  assign popcount39_35p6_core_225 = input_a[34] & input_a[8];
  assign popcount39_35p6_core_226 = ~input_a[37];
  assign popcount39_35p6_core_227 = ~(input_a[37] | input_a[6]);
  assign popcount39_35p6_core_228 = input_a[36] ^ popcount39_35p6_core_226;
  assign popcount39_35p6_core_229 = input_a[36] & popcount39_35p6_core_226;
  assign popcount39_35p6_core_230 = popcount39_35p6_core_227 ^ popcount39_35p6_core_229;
  assign popcount39_35p6_core_231 = popcount39_35p6_core_227 & popcount39_35p6_core_229;
  assign popcount39_35p6_core_232 = input_a[34] ^ popcount39_35p6_core_228;
  assign popcount39_35p6_core_233 = input_a[34] & popcount39_35p6_core_228;
  assign popcount39_35p6_core_234 = input_a[23] | popcount39_35p6_core_230;
  assign popcount39_35p6_core_235 = popcount39_35p6_core_225 & popcount39_35p6_core_230;
  assign popcount39_35p6_core_236 = popcount39_35p6_core_234 ^ popcount39_35p6_core_233;
  assign popcount39_35p6_core_237 = input_a[17] & popcount39_35p6_core_233;
  assign popcount39_35p6_core_238 = popcount39_35p6_core_235 | popcount39_35p6_core_237;
  assign popcount39_35p6_core_239 = popcount39_35p6_core_231 ^ popcount39_35p6_core_238;
  assign popcount39_35p6_core_240 = popcount39_35p6_core_231 & popcount39_35p6_core_238;
  assign popcount39_35p6_core_241 = popcount39_35p6_core_215 ^ popcount39_35p6_core_232;
  assign popcount39_35p6_core_242 = popcount39_35p6_core_215 & popcount39_35p6_core_232;
  assign popcount39_35p6_core_243 = popcount39_35p6_core_219 ^ input_a[7];
  assign popcount39_35p6_core_244 = popcount39_35p6_core_219 & popcount39_35p6_core_236;
  assign popcount39_35p6_core_245 = popcount39_35p6_core_243 ^ popcount39_35p6_core_242;
  assign popcount39_35p6_core_246 = popcount39_35p6_core_243 & popcount39_35p6_core_242;
  assign popcount39_35p6_core_247 = popcount39_35p6_core_244 | popcount39_35p6_core_246;
  assign popcount39_35p6_core_248 = popcount39_35p6_core_222 ^ popcount39_35p6_core_239;
  assign popcount39_35p6_core_249 = popcount39_35p6_core_222 & popcount39_35p6_core_239;
  assign popcount39_35p6_core_250 = popcount39_35p6_core_248 ^ popcount39_35p6_core_247;
  assign popcount39_35p6_core_251 = popcount39_35p6_core_248 & popcount39_35p6_core_247;
  assign popcount39_35p6_core_252 = popcount39_35p6_core_249 | popcount39_35p6_core_251;
  assign popcount39_35p6_core_253 = popcount39_35p6_core_223 ^ popcount39_35p6_core_240;
  assign popcount39_35p6_core_254 = popcount39_35p6_core_223 & popcount39_35p6_core_240;
  assign popcount39_35p6_core_255 = popcount39_35p6_core_253 ^ popcount39_35p6_core_252;
  assign popcount39_35p6_core_256 = popcount39_35p6_core_253 & input_a[31];
  assign popcount39_35p6_core_257 = popcount39_35p6_core_254 | popcount39_35p6_core_256;
  assign popcount39_35p6_core_258 = popcount39_35p6_core_190 ^ popcount39_35p6_core_241;
  assign popcount39_35p6_core_259 = ~(popcount39_35p6_core_190 | popcount39_35p6_core_241);
  assign popcount39_35p6_core_260 = popcount39_35p6_core_192 ^ popcount39_35p6_core_245;
  assign popcount39_35p6_core_261 = popcount39_35p6_core_192 & input_a[1];
  assign popcount39_35p6_core_262 = popcount39_35p6_core_260 ^ popcount39_35p6_core_259;
  assign popcount39_35p6_core_263 = popcount39_35p6_core_260 & popcount39_35p6_core_259;
  assign popcount39_35p6_core_264 = popcount39_35p6_core_261 | popcount39_35p6_core_263;
  assign popcount39_35p6_core_265 = popcount39_35p6_core_199 ^ input_a[18];
  assign popcount39_35p6_core_266 = popcount39_35p6_core_199 & popcount39_35p6_core_250;
  assign popcount39_35p6_core_267 = ~popcount39_35p6_core_265;
  assign popcount39_35p6_core_268 = popcount39_35p6_core_265 & input_a[7];
  assign popcount39_35p6_core_269 = input_a[16] | popcount39_35p6_core_268;
  assign popcount39_35p6_core_270 = popcount39_35p6_core_204 ^ popcount39_35p6_core_255;
  assign popcount39_35p6_core_271 = popcount39_35p6_core_204 & popcount39_35p6_core_255;
  assign popcount39_35p6_core_272 = ~popcount39_35p6_core_270;
  assign popcount39_35p6_core_273 = popcount39_35p6_core_270 & popcount39_35p6_core_269;
  assign popcount39_35p6_core_274 = popcount39_35p6_core_271 | popcount39_35p6_core_273;
  assign popcount39_35p6_core_282 = popcount39_35p6_core_136 & popcount39_35p6_core_262;
  assign popcount39_35p6_core_283 = input_a[34] & popcount39_35p6_core_262;
  assign popcount39_35p6_core_287 = popcount39_35p6_core_143 & popcount39_35p6_core_267;
  assign popcount39_35p6_core_288 = popcount39_35p6_core_143 & popcount39_35p6_core_267;
  assign popcount39_35p6_core_290 = popcount39_35p6_core_287 & popcount39_35p6_core_283;
  assign popcount39_35p6_core_291 = popcount39_35p6_core_288 | popcount39_35p6_core_290;
  assign popcount39_35p6_core_292 = popcount39_35p6_core_148 ^ popcount39_35p6_core_272;
  assign popcount39_35p6_core_293 = popcount39_35p6_core_148 & popcount39_35p6_core_272;
  assign popcount39_35p6_core_294 = popcount39_35p6_core_292 ^ popcount39_35p6_core_291;
  assign popcount39_35p6_core_295 = popcount39_35p6_core_292 & popcount39_35p6_core_291;
  assign popcount39_35p6_core_296 = popcount39_35p6_core_293 | popcount39_35p6_core_295;
  assign popcount39_35p6_core_297 = popcount39_35p6_core_150 ^ popcount39_35p6_core_274;
  assign popcount39_35p6_core_298 = popcount39_35p6_core_150 & popcount39_35p6_core_274;
  assign popcount39_35p6_core_299 = popcount39_35p6_core_297 ^ popcount39_35p6_core_296;
  assign popcount39_35p6_core_300 = popcount39_35p6_core_297 & popcount39_35p6_core_296;
  assign popcount39_35p6_core_301 = popcount39_35p6_core_298 | popcount39_35p6_core_300;

  assign popcount39_35p6_out[0] = popcount39_35p6_core_107;
  assign popcount39_35p6_out[1] = input_a[31];
  assign popcount39_35p6_out[2] = 1'b0;
  assign popcount39_35p6_out[3] = popcount39_35p6_core_294;
  assign popcount39_35p6_out[4] = popcount39_35p6_core_299;
  assign popcount39_35p6_out[5] = popcount39_35p6_core_301;
endmodule