// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.09375
// WCE=4.0
// EP=0.726562%
// Printed PDK parameters:
//  Area=42422784.0
//  Delay=73572008.0
//  Power=1807900.0

module popcount20_8y0h(input [19:0] input_a, output [4:0] popcount20_8y0h_out);
  wire popcount20_8y0h_core_022;
  wire popcount20_8y0h_core_023;
  wire popcount20_8y0h_core_024;
  wire popcount20_8y0h_core_025;
  wire popcount20_8y0h_core_026;
  wire popcount20_8y0h_core_028;
  wire popcount20_8y0h_core_029;
  wire popcount20_8y0h_core_030;
  wire popcount20_8y0h_core_031;
  wire popcount20_8y0h_core_032;
  wire popcount20_8y0h_core_033;
  wire popcount20_8y0h_core_034;
  wire popcount20_8y0h_core_035;
  wire popcount20_8y0h_core_036;
  wire popcount20_8y0h_core_037;
  wire popcount20_8y0h_core_038_not;
  wire popcount20_8y0h_core_039;
  wire popcount20_8y0h_core_040;
  wire popcount20_8y0h_core_041;
  wire popcount20_8y0h_core_042;
  wire popcount20_8y0h_core_043;
  wire popcount20_8y0h_core_044;
  wire popcount20_8y0h_core_045;
  wire popcount20_8y0h_core_047;
  wire popcount20_8y0h_core_048;
  wire popcount20_8y0h_core_049;
  wire popcount20_8y0h_core_050;
  wire popcount20_8y0h_core_051;
  wire popcount20_8y0h_core_052;
  wire popcount20_8y0h_core_053;
  wire popcount20_8y0h_core_055;
  wire popcount20_8y0h_core_056;
  wire popcount20_8y0h_core_057;
  wire popcount20_8y0h_core_058;
  wire popcount20_8y0h_core_059;
  wire popcount20_8y0h_core_060;
  wire popcount20_8y0h_core_061;
  wire popcount20_8y0h_core_062;
  wire popcount20_8y0h_core_063;
  wire popcount20_8y0h_core_064;
  wire popcount20_8y0h_core_065;
  wire popcount20_8y0h_core_066;
  wire popcount20_8y0h_core_067;
  wire popcount20_8y0h_core_071;
  wire popcount20_8y0h_core_074;
  wire popcount20_8y0h_core_075;
  wire popcount20_8y0h_core_076_not;
  wire popcount20_8y0h_core_077;
  wire popcount20_8y0h_core_078;
  wire popcount20_8y0h_core_079;
  wire popcount20_8y0h_core_081;
  wire popcount20_8y0h_core_083;
  wire popcount20_8y0h_core_084;
  wire popcount20_8y0h_core_089;
  wire popcount20_8y0h_core_090;
  wire popcount20_8y0h_core_091;
  wire popcount20_8y0h_core_092;
  wire popcount20_8y0h_core_094;
  wire popcount20_8y0h_core_095;
  wire popcount20_8y0h_core_096;
  wire popcount20_8y0h_core_097;
  wire popcount20_8y0h_core_098_not;
  wire popcount20_8y0h_core_100;
  wire popcount20_8y0h_core_102;
  wire popcount20_8y0h_core_103;
  wire popcount20_8y0h_core_104;
  wire popcount20_8y0h_core_105;
  wire popcount20_8y0h_core_106;
  wire popcount20_8y0h_core_108;
  wire popcount20_8y0h_core_109;
  wire popcount20_8y0h_core_110;
  wire popcount20_8y0h_core_111;
  wire popcount20_8y0h_core_112;
  wire popcount20_8y0h_core_113;
  wire popcount20_8y0h_core_116;
  wire popcount20_8y0h_core_117;
  wire popcount20_8y0h_core_122;
  wire popcount20_8y0h_core_123;
  wire popcount20_8y0h_core_125;
  wire popcount20_8y0h_core_126;
  wire popcount20_8y0h_core_127;
  wire popcount20_8y0h_core_128;
  wire popcount20_8y0h_core_129;
  wire popcount20_8y0h_core_130;
  wire popcount20_8y0h_core_131;
  wire popcount20_8y0h_core_132;
  wire popcount20_8y0h_core_133;
  wire popcount20_8y0h_core_134;
  wire popcount20_8y0h_core_135;
  wire popcount20_8y0h_core_136;
  wire popcount20_8y0h_core_137;
  wire popcount20_8y0h_core_138;
  wire popcount20_8y0h_core_139;
  wire popcount20_8y0h_core_140;
  wire popcount20_8y0h_core_142;

  assign popcount20_8y0h_core_022 = input_a[0] ^ input_a[1];
  assign popcount20_8y0h_core_023 = input_a[0] & input_a[1];
  assign popcount20_8y0h_core_024 = ~(input_a[12] & input_a[7]);
  assign popcount20_8y0h_core_025 = input_a[3] & input_a[4];
  assign popcount20_8y0h_core_026 = ~input_a[2];
  assign popcount20_8y0h_core_028 = popcount20_8y0h_core_025 ^ input_a[2];
  assign popcount20_8y0h_core_029 = popcount20_8y0h_core_025 & input_a[2];
  assign popcount20_8y0h_core_030 = popcount20_8y0h_core_022 ^ popcount20_8y0h_core_026;
  assign popcount20_8y0h_core_031 = popcount20_8y0h_core_022 & popcount20_8y0h_core_026;
  assign popcount20_8y0h_core_032 = popcount20_8y0h_core_023 ^ popcount20_8y0h_core_028;
  assign popcount20_8y0h_core_033 = popcount20_8y0h_core_023 & popcount20_8y0h_core_028;
  assign popcount20_8y0h_core_034 = popcount20_8y0h_core_032 ^ popcount20_8y0h_core_031;
  assign popcount20_8y0h_core_035 = popcount20_8y0h_core_032 & popcount20_8y0h_core_031;
  assign popcount20_8y0h_core_036 = popcount20_8y0h_core_033 | popcount20_8y0h_core_035;
  assign popcount20_8y0h_core_037 = popcount20_8y0h_core_029 | popcount20_8y0h_core_036;
  assign popcount20_8y0h_core_038_not = ~input_a[14];
  assign popcount20_8y0h_core_039 = input_a[5] ^ input_a[6];
  assign popcount20_8y0h_core_040 = input_a[5] & input_a[6];
  assign popcount20_8y0h_core_041 = input_a[8] ^ input_a[9];
  assign popcount20_8y0h_core_042 = input_a[8] & input_a[9];
  assign popcount20_8y0h_core_043 = input_a[7] ^ popcount20_8y0h_core_041;
  assign popcount20_8y0h_core_044 = input_a[7] & popcount20_8y0h_core_041;
  assign popcount20_8y0h_core_045 = popcount20_8y0h_core_042 | popcount20_8y0h_core_044;
  assign popcount20_8y0h_core_047 = ~(input_a[3] & input_a[11]);
  assign popcount20_8y0h_core_048 = popcount20_8y0h_core_039 & popcount20_8y0h_core_043;
  assign popcount20_8y0h_core_049 = popcount20_8y0h_core_040 ^ popcount20_8y0h_core_045;
  assign popcount20_8y0h_core_050 = popcount20_8y0h_core_040 & popcount20_8y0h_core_045;
  assign popcount20_8y0h_core_051 = popcount20_8y0h_core_049 ^ popcount20_8y0h_core_048;
  assign popcount20_8y0h_core_052 = popcount20_8y0h_core_049 & popcount20_8y0h_core_048;
  assign popcount20_8y0h_core_053 = popcount20_8y0h_core_050 | popcount20_8y0h_core_052;
  assign popcount20_8y0h_core_055 = input_a[17] ^ input_a[16];
  assign popcount20_8y0h_core_056 = input_a[0] ^ input_a[12];
  assign popcount20_8y0h_core_057 = popcount20_8y0h_core_030 & input_a[18];
  assign popcount20_8y0h_core_058 = popcount20_8y0h_core_034 ^ popcount20_8y0h_core_051;
  assign popcount20_8y0h_core_059 = popcount20_8y0h_core_034 & popcount20_8y0h_core_051;
  assign popcount20_8y0h_core_060 = popcount20_8y0h_core_058 ^ popcount20_8y0h_core_057;
  assign popcount20_8y0h_core_061 = popcount20_8y0h_core_058 & popcount20_8y0h_core_057;
  assign popcount20_8y0h_core_062 = popcount20_8y0h_core_059 | popcount20_8y0h_core_061;
  assign popcount20_8y0h_core_063 = popcount20_8y0h_core_037 ^ popcount20_8y0h_core_053;
  assign popcount20_8y0h_core_064 = popcount20_8y0h_core_037 & popcount20_8y0h_core_053;
  assign popcount20_8y0h_core_065 = popcount20_8y0h_core_063 ^ popcount20_8y0h_core_062;
  assign popcount20_8y0h_core_066 = popcount20_8y0h_core_063 & popcount20_8y0h_core_062;
  assign popcount20_8y0h_core_067 = popcount20_8y0h_core_064 | popcount20_8y0h_core_066;
  assign popcount20_8y0h_core_071 = ~(input_a[18] ^ input_a[14]);
  assign popcount20_8y0h_core_074 = input_a[10] & input_a[12];
  assign popcount20_8y0h_core_075 = ~input_a[11];
  assign popcount20_8y0h_core_076_not = ~input_a[11];
  assign popcount20_8y0h_core_077 = input_a[4] ^ input_a[8];
  assign popcount20_8y0h_core_078 = ~(input_a[3] & input_a[17]);
  assign popcount20_8y0h_core_079 = input_a[16] | input_a[19];
  assign popcount20_8y0h_core_081 = input_a[3] | input_a[8];
  assign popcount20_8y0h_core_083 = popcount20_8y0h_core_074 ^ popcount20_8y0h_core_079;
  assign popcount20_8y0h_core_084 = popcount20_8y0h_core_074 & popcount20_8y0h_core_079;
  assign popcount20_8y0h_core_089 = input_a[0] ^ input_a[19];
  assign popcount20_8y0h_core_090 = ~(input_a[6] | input_a[5]);
  assign popcount20_8y0h_core_091 = input_a[11] ^ input_a[16];
  assign popcount20_8y0h_core_092 = ~(input_a[17] ^ input_a[7]);
  assign popcount20_8y0h_core_094 = ~(input_a[8] ^ input_a[4]);
  assign popcount20_8y0h_core_095 = input_a[16] & input_a[1];
  assign popcount20_8y0h_core_096 = input_a[12] ^ input_a[5];
  assign popcount20_8y0h_core_097 = input_a[11] ^ input_a[14];
  assign popcount20_8y0h_core_098_not = ~input_a[9];
  assign popcount20_8y0h_core_100 = ~(input_a[17] & input_a[7]);
  assign popcount20_8y0h_core_102 = input_a[14] | input_a[17];
  assign popcount20_8y0h_core_103 = input_a[12] ^ input_a[9];
  assign popcount20_8y0h_core_104 = input_a[3] | input_a[13];
  assign popcount20_8y0h_core_105 = ~(input_a[10] & input_a[19]);
  assign popcount20_8y0h_core_106 = input_a[3] & input_a[0];
  assign popcount20_8y0h_core_108 = ~(input_a[7] | input_a[7]);
  assign popcount20_8y0h_core_109 = popcount20_8y0h_core_083 ^ popcount20_8y0h_core_102;
  assign popcount20_8y0h_core_110 = popcount20_8y0h_core_083 & popcount20_8y0h_core_102;
  assign popcount20_8y0h_core_111 = popcount20_8y0h_core_109 ^ input_a[11];
  assign popcount20_8y0h_core_112 = popcount20_8y0h_core_109 & input_a[11];
  assign popcount20_8y0h_core_113 = popcount20_8y0h_core_110 | popcount20_8y0h_core_112;
  assign popcount20_8y0h_core_116 = popcount20_8y0h_core_084 ^ popcount20_8y0h_core_113;
  assign popcount20_8y0h_core_117 = popcount20_8y0h_core_084 & popcount20_8y0h_core_113;
  assign popcount20_8y0h_core_122 = ~(input_a[5] ^ input_a[4]);
  assign popcount20_8y0h_core_123 = ~input_a[17];
  assign popcount20_8y0h_core_125 = input_a[13] & input_a[15];
  assign popcount20_8y0h_core_126 = popcount20_8y0h_core_060 ^ popcount20_8y0h_core_111;
  assign popcount20_8y0h_core_127 = popcount20_8y0h_core_060 & popcount20_8y0h_core_111;
  assign popcount20_8y0h_core_128 = popcount20_8y0h_core_126 ^ popcount20_8y0h_core_125;
  assign popcount20_8y0h_core_129 = popcount20_8y0h_core_126 & popcount20_8y0h_core_125;
  assign popcount20_8y0h_core_130 = popcount20_8y0h_core_127 | popcount20_8y0h_core_129;
  assign popcount20_8y0h_core_131 = popcount20_8y0h_core_065 ^ popcount20_8y0h_core_116;
  assign popcount20_8y0h_core_132 = popcount20_8y0h_core_065 & popcount20_8y0h_core_116;
  assign popcount20_8y0h_core_133 = popcount20_8y0h_core_131 ^ popcount20_8y0h_core_130;
  assign popcount20_8y0h_core_134 = popcount20_8y0h_core_131 & popcount20_8y0h_core_130;
  assign popcount20_8y0h_core_135 = popcount20_8y0h_core_132 | popcount20_8y0h_core_134;
  assign popcount20_8y0h_core_136 = popcount20_8y0h_core_067 ^ popcount20_8y0h_core_117;
  assign popcount20_8y0h_core_137 = popcount20_8y0h_core_067 & popcount20_8y0h_core_117;
  assign popcount20_8y0h_core_138 = popcount20_8y0h_core_136 ^ popcount20_8y0h_core_135;
  assign popcount20_8y0h_core_139 = popcount20_8y0h_core_136 & popcount20_8y0h_core_135;
  assign popcount20_8y0h_core_140 = popcount20_8y0h_core_137 | popcount20_8y0h_core_139;
  assign popcount20_8y0h_core_142 = ~(input_a[9] ^ input_a[14]);

  assign popcount20_8y0h_out[0] = 1'b0;
  assign popcount20_8y0h_out[1] = popcount20_8y0h_core_128;
  assign popcount20_8y0h_out[2] = popcount20_8y0h_core_133;
  assign popcount20_8y0h_out[3] = popcount20_8y0h_core_138;
  assign popcount20_8y0h_out[4] = popcount20_8y0h_core_140;
endmodule