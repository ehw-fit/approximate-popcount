// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=5.12141
// WCE=22.0
// EP=0.929557%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_vk7b(input [28:0] input_a, output [4:0] popcount29_vk7b_out);
  wire popcount29_vk7b_core_033;
  wire popcount29_vk7b_core_034;
  wire popcount29_vk7b_core_036;
  wire popcount29_vk7b_core_037;
  wire popcount29_vk7b_core_039;
  wire popcount29_vk7b_core_040;
  wire popcount29_vk7b_core_041;
  wire popcount29_vk7b_core_042;
  wire popcount29_vk7b_core_043;
  wire popcount29_vk7b_core_048;
  wire popcount29_vk7b_core_049;
  wire popcount29_vk7b_core_050;
  wire popcount29_vk7b_core_051;
  wire popcount29_vk7b_core_053;
  wire popcount29_vk7b_core_055;
  wire popcount29_vk7b_core_059;
  wire popcount29_vk7b_core_060;
  wire popcount29_vk7b_core_064;
  wire popcount29_vk7b_core_065;
  wire popcount29_vk7b_core_066;
  wire popcount29_vk7b_core_067;
  wire popcount29_vk7b_core_069;
  wire popcount29_vk7b_core_070;
  wire popcount29_vk7b_core_071;
  wire popcount29_vk7b_core_072;
  wire popcount29_vk7b_core_073;
  wire popcount29_vk7b_core_074;
  wire popcount29_vk7b_core_075;
  wire popcount29_vk7b_core_076;
  wire popcount29_vk7b_core_078;
  wire popcount29_vk7b_core_079;
  wire popcount29_vk7b_core_080;
  wire popcount29_vk7b_core_081;
  wire popcount29_vk7b_core_082;
  wire popcount29_vk7b_core_084;
  wire popcount29_vk7b_core_085;
  wire popcount29_vk7b_core_087;
  wire popcount29_vk7b_core_089;
  wire popcount29_vk7b_core_090;
  wire popcount29_vk7b_core_091;
  wire popcount29_vk7b_core_095_not;
  wire popcount29_vk7b_core_096_not;
  wire popcount29_vk7b_core_097;
  wire popcount29_vk7b_core_098;
  wire popcount29_vk7b_core_100;
  wire popcount29_vk7b_core_101;
  wire popcount29_vk7b_core_102;
  wire popcount29_vk7b_core_105;
  wire popcount29_vk7b_core_106;
  wire popcount29_vk7b_core_108;
  wire popcount29_vk7b_core_112;
  wire popcount29_vk7b_core_115;
  wire popcount29_vk7b_core_116;
  wire popcount29_vk7b_core_118;
  wire popcount29_vk7b_core_119;
  wire popcount29_vk7b_core_121;
  wire popcount29_vk7b_core_122;
  wire popcount29_vk7b_core_123;
  wire popcount29_vk7b_core_124;
  wire popcount29_vk7b_core_126;
  wire popcount29_vk7b_core_129;
  wire popcount29_vk7b_core_130;
  wire popcount29_vk7b_core_133;
  wire popcount29_vk7b_core_135;
  wire popcount29_vk7b_core_137;
  wire popcount29_vk7b_core_138;
  wire popcount29_vk7b_core_139;
  wire popcount29_vk7b_core_143;
  wire popcount29_vk7b_core_144;
  wire popcount29_vk7b_core_145;
  wire popcount29_vk7b_core_146;
  wire popcount29_vk7b_core_147;
  wire popcount29_vk7b_core_150;
  wire popcount29_vk7b_core_152;
  wire popcount29_vk7b_core_154;
  wire popcount29_vk7b_core_155;
  wire popcount29_vk7b_core_156;
  wire popcount29_vk7b_core_157;
  wire popcount29_vk7b_core_158;
  wire popcount29_vk7b_core_159;
  wire popcount29_vk7b_core_160;
  wire popcount29_vk7b_core_164;
  wire popcount29_vk7b_core_165;
  wire popcount29_vk7b_core_166;
  wire popcount29_vk7b_core_167;
  wire popcount29_vk7b_core_168;
  wire popcount29_vk7b_core_169;
  wire popcount29_vk7b_core_170;
  wire popcount29_vk7b_core_172;
  wire popcount29_vk7b_core_174;
  wire popcount29_vk7b_core_175;
  wire popcount29_vk7b_core_176;
  wire popcount29_vk7b_core_178;
  wire popcount29_vk7b_core_179;
  wire popcount29_vk7b_core_180;
  wire popcount29_vk7b_core_181;
  wire popcount29_vk7b_core_182;
  wire popcount29_vk7b_core_183;
  wire popcount29_vk7b_core_184_not;
  wire popcount29_vk7b_core_187;
  wire popcount29_vk7b_core_188;
  wire popcount29_vk7b_core_189;
  wire popcount29_vk7b_core_190;
  wire popcount29_vk7b_core_191;
  wire popcount29_vk7b_core_192;
  wire popcount29_vk7b_core_193;
  wire popcount29_vk7b_core_194;
  wire popcount29_vk7b_core_195;
  wire popcount29_vk7b_core_198;
  wire popcount29_vk7b_core_201;
  wire popcount29_vk7b_core_202;
  wire popcount29_vk7b_core_203;
  wire popcount29_vk7b_core_204_not;
  wire popcount29_vk7b_core_205;

  assign popcount29_vk7b_core_033 = ~(input_a[15] | input_a[18]);
  assign popcount29_vk7b_core_034 = ~(input_a[12] & input_a[5]);
  assign popcount29_vk7b_core_036 = ~(input_a[19] ^ input_a[11]);
  assign popcount29_vk7b_core_037 = ~(input_a[28] & input_a[13]);
  assign popcount29_vk7b_core_039 = input_a[13] | input_a[21];
  assign popcount29_vk7b_core_040 = ~input_a[8];
  assign popcount29_vk7b_core_041 = input_a[0] | input_a[22];
  assign popcount29_vk7b_core_042 = ~(input_a[3] & input_a[2]);
  assign popcount29_vk7b_core_043 = ~(input_a[4] | input_a[23]);
  assign popcount29_vk7b_core_048 = input_a[20] & input_a[3];
  assign popcount29_vk7b_core_049 = ~(input_a[25] ^ input_a[0]);
  assign popcount29_vk7b_core_050 = ~(input_a[28] | input_a[25]);
  assign popcount29_vk7b_core_051 = input_a[2] & input_a[17];
  assign popcount29_vk7b_core_053 = ~(input_a[10] & input_a[2]);
  assign popcount29_vk7b_core_055 = ~(input_a[17] ^ input_a[10]);
  assign popcount29_vk7b_core_059 = input_a[5] ^ input_a[6];
  assign popcount29_vk7b_core_060 = ~(input_a[28] | input_a[4]);
  assign popcount29_vk7b_core_064 = ~(input_a[4] ^ input_a[20]);
  assign popcount29_vk7b_core_065 = ~input_a[2];
  assign popcount29_vk7b_core_066 = ~(input_a[4] ^ input_a[7]);
  assign popcount29_vk7b_core_067 = ~(input_a[17] | input_a[19]);
  assign popcount29_vk7b_core_069 = input_a[16] | input_a[19];
  assign popcount29_vk7b_core_070 = ~input_a[15];
  assign popcount29_vk7b_core_071 = ~(input_a[21] & input_a[4]);
  assign popcount29_vk7b_core_072 = ~(input_a[28] | input_a[3]);
  assign popcount29_vk7b_core_073 = ~(input_a[17] ^ input_a[18]);
  assign popcount29_vk7b_core_074 = ~(input_a[24] & input_a[19]);
  assign popcount29_vk7b_core_075 = input_a[20] & input_a[12];
  assign popcount29_vk7b_core_076 = ~input_a[26];
  assign popcount29_vk7b_core_078 = input_a[16] & input_a[19];
  assign popcount29_vk7b_core_079 = input_a[16] | input_a[1];
  assign popcount29_vk7b_core_080 = input_a[5] & input_a[0];
  assign popcount29_vk7b_core_081 = input_a[25] & input_a[23];
  assign popcount29_vk7b_core_082 = ~(input_a[8] & input_a[9]);
  assign popcount29_vk7b_core_084 = ~(input_a[7] | input_a[12]);
  assign popcount29_vk7b_core_085 = ~(input_a[5] | input_a[21]);
  assign popcount29_vk7b_core_087 = ~(input_a[12] & input_a[26]);
  assign popcount29_vk7b_core_089 = input_a[3] ^ input_a[23];
  assign popcount29_vk7b_core_090 = input_a[17] | input_a[12];
  assign popcount29_vk7b_core_091 = ~input_a[9];
  assign popcount29_vk7b_core_095_not = ~input_a[23];
  assign popcount29_vk7b_core_096_not = ~input_a[3];
  assign popcount29_vk7b_core_097 = ~(input_a[28] & input_a[23]);
  assign popcount29_vk7b_core_098 = input_a[24] | input_a[19];
  assign popcount29_vk7b_core_100 = ~(input_a[19] | input_a[0]);
  assign popcount29_vk7b_core_101 = ~input_a[20];
  assign popcount29_vk7b_core_102 = ~(input_a[27] ^ input_a[20]);
  assign popcount29_vk7b_core_105 = ~(input_a[3] & input_a[18]);
  assign popcount29_vk7b_core_106 = input_a[4] & input_a[21];
  assign popcount29_vk7b_core_108 = input_a[28] | input_a[22];
  assign popcount29_vk7b_core_112 = input_a[24] & input_a[7];
  assign popcount29_vk7b_core_115 = ~(input_a[7] | input_a[24]);
  assign popcount29_vk7b_core_116 = ~(input_a[14] & input_a[3]);
  assign popcount29_vk7b_core_118 = ~input_a[15];
  assign popcount29_vk7b_core_119 = input_a[12] | input_a[23];
  assign popcount29_vk7b_core_121 = ~input_a[1];
  assign popcount29_vk7b_core_122 = ~input_a[1];
  assign popcount29_vk7b_core_123 = input_a[2] | input_a[23];
  assign popcount29_vk7b_core_124 = input_a[10] | input_a[20];
  assign popcount29_vk7b_core_126 = input_a[2] & input_a[15];
  assign popcount29_vk7b_core_129 = ~(input_a[12] & input_a[8]);
  assign popcount29_vk7b_core_130 = ~(input_a[20] ^ input_a[1]);
  assign popcount29_vk7b_core_133 = ~input_a[21];
  assign popcount29_vk7b_core_135 = input_a[20] ^ input_a[25];
  assign popcount29_vk7b_core_137 = ~(input_a[26] | input_a[0]);
  assign popcount29_vk7b_core_138 = input_a[21] ^ input_a[28];
  assign popcount29_vk7b_core_139 = ~(input_a[4] | input_a[12]);
  assign popcount29_vk7b_core_143 = ~(input_a[18] ^ input_a[22]);
  assign popcount29_vk7b_core_144 = input_a[6] & input_a[3];
  assign popcount29_vk7b_core_145 = ~input_a[19];
  assign popcount29_vk7b_core_146 = input_a[19] ^ input_a[28];
  assign popcount29_vk7b_core_147 = ~(input_a[7] | input_a[3]);
  assign popcount29_vk7b_core_150 = ~(input_a[9] ^ input_a[9]);
  assign popcount29_vk7b_core_152 = ~input_a[5];
  assign popcount29_vk7b_core_154 = input_a[8] | input_a[23];
  assign popcount29_vk7b_core_155 = input_a[14] ^ input_a[11];
  assign popcount29_vk7b_core_156 = input_a[3] & input_a[28];
  assign popcount29_vk7b_core_157 = ~(input_a[14] | input_a[27]);
  assign popcount29_vk7b_core_158 = ~(input_a[16] ^ input_a[18]);
  assign popcount29_vk7b_core_159 = ~(input_a[7] ^ input_a[21]);
  assign popcount29_vk7b_core_160 = ~(input_a[27] | input_a[1]);
  assign popcount29_vk7b_core_164 = ~input_a[28];
  assign popcount29_vk7b_core_165 = input_a[18] & input_a[22];
  assign popcount29_vk7b_core_166 = ~(input_a[14] & input_a[21]);
  assign popcount29_vk7b_core_167 = ~(input_a[11] ^ input_a[19]);
  assign popcount29_vk7b_core_168 = input_a[11] ^ input_a[24];
  assign popcount29_vk7b_core_169 = input_a[15] ^ input_a[19];
  assign popcount29_vk7b_core_170 = input_a[21] & input_a[26];
  assign popcount29_vk7b_core_172 = ~(input_a[25] ^ input_a[24]);
  assign popcount29_vk7b_core_174 = input_a[24] ^ input_a[14];
  assign popcount29_vk7b_core_175 = ~input_a[19];
  assign popcount29_vk7b_core_176 = ~input_a[16];
  assign popcount29_vk7b_core_178 = input_a[14] | input_a[10];
  assign popcount29_vk7b_core_179 = ~(input_a[2] & input_a[20]);
  assign popcount29_vk7b_core_180 = ~(input_a[20] ^ input_a[0]);
  assign popcount29_vk7b_core_181 = ~(input_a[26] | input_a[22]);
  assign popcount29_vk7b_core_182 = ~(input_a[17] & input_a[7]);
  assign popcount29_vk7b_core_183 = ~(input_a[14] ^ input_a[16]);
  assign popcount29_vk7b_core_184_not = ~input_a[6];
  assign popcount29_vk7b_core_187 = ~input_a[9];
  assign popcount29_vk7b_core_188 = ~(input_a[28] | input_a[19]);
  assign popcount29_vk7b_core_189 = input_a[21] & input_a[15];
  assign popcount29_vk7b_core_190 = input_a[22] | input_a[17];
  assign popcount29_vk7b_core_191 = ~(input_a[1] & input_a[16]);
  assign popcount29_vk7b_core_192 = input_a[3] ^ input_a[24];
  assign popcount29_vk7b_core_193 = ~(input_a[10] | input_a[18]);
  assign popcount29_vk7b_core_194 = ~(input_a[7] | input_a[2]);
  assign popcount29_vk7b_core_195 = input_a[22] | input_a[21];
  assign popcount29_vk7b_core_198 = input_a[11] ^ input_a[19];
  assign popcount29_vk7b_core_201 = ~(input_a[16] & input_a[17]);
  assign popcount29_vk7b_core_202 = ~(input_a[16] | input_a[10]);
  assign popcount29_vk7b_core_203 = ~(input_a[6] | input_a[20]);
  assign popcount29_vk7b_core_204_not = ~input_a[26];
  assign popcount29_vk7b_core_205 = ~(input_a[23] | input_a[8]);

  assign popcount29_vk7b_out[0] = 1'b0;
  assign popcount29_vk7b_out[1] = 1'b1;
  assign popcount29_vk7b_out[2] = 1'b1;
  assign popcount29_vk7b_out[3] = input_a[8];
  assign popcount29_vk7b_out[4] = 1'b0;
endmodule