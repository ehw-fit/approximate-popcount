// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.01475
// WCE=13.0
// EP=0.845019%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_xcpf(input [26:0] input_a, output [4:0] popcount27_xcpf_out);
  wire popcount27_xcpf_core_033;
  wire popcount27_xcpf_core_035;
  wire popcount27_xcpf_core_036;
  wire popcount27_xcpf_core_037;
  wire popcount27_xcpf_core_038;
  wire popcount27_xcpf_core_042;
  wire popcount27_xcpf_core_043;
  wire popcount27_xcpf_core_044;
  wire popcount27_xcpf_core_045;
  wire popcount27_xcpf_core_046;
  wire popcount27_xcpf_core_047;
  wire popcount27_xcpf_core_048;
  wire popcount27_xcpf_core_050;
  wire popcount27_xcpf_core_051;
  wire popcount27_xcpf_core_052;
  wire popcount27_xcpf_core_056;
  wire popcount27_xcpf_core_057;
  wire popcount27_xcpf_core_058;
  wire popcount27_xcpf_core_059;
  wire popcount27_xcpf_core_060;
  wire popcount27_xcpf_core_063;
  wire popcount27_xcpf_core_064;
  wire popcount27_xcpf_core_065;
  wire popcount27_xcpf_core_066;
  wire popcount27_xcpf_core_067;
  wire popcount27_xcpf_core_068;
  wire popcount27_xcpf_core_069;
  wire popcount27_xcpf_core_072;
  wire popcount27_xcpf_core_076;
  wire popcount27_xcpf_core_077;
  wire popcount27_xcpf_core_078;
  wire popcount27_xcpf_core_079;
  wire popcount27_xcpf_core_080;
  wire popcount27_xcpf_core_082;
  wire popcount27_xcpf_core_084;
  wire popcount27_xcpf_core_087;
  wire popcount27_xcpf_core_088;
  wire popcount27_xcpf_core_091;
  wire popcount27_xcpf_core_092;
  wire popcount27_xcpf_core_094;
  wire popcount27_xcpf_core_095_not;
  wire popcount27_xcpf_core_099;
  wire popcount27_xcpf_core_102;
  wire popcount27_xcpf_core_103;
  wire popcount27_xcpf_core_104;
  wire popcount27_xcpf_core_108;
  wire popcount27_xcpf_core_109;
  wire popcount27_xcpf_core_110;
  wire popcount27_xcpf_core_111;
  wire popcount27_xcpf_core_113;
  wire popcount27_xcpf_core_114;
  wire popcount27_xcpf_core_115;
  wire popcount27_xcpf_core_116;
  wire popcount27_xcpf_core_117;
  wire popcount27_xcpf_core_119;
  wire popcount27_xcpf_core_120;
  wire popcount27_xcpf_core_122;
  wire popcount27_xcpf_core_125;
  wire popcount27_xcpf_core_126;
  wire popcount27_xcpf_core_129;
  wire popcount27_xcpf_core_130;
  wire popcount27_xcpf_core_131;
  wire popcount27_xcpf_core_133;
  wire popcount27_xcpf_core_135;
  wire popcount27_xcpf_core_136;
  wire popcount27_xcpf_core_137;
  wire popcount27_xcpf_core_138;
  wire popcount27_xcpf_core_139;
  wire popcount27_xcpf_core_140;
  wire popcount27_xcpf_core_141;
  wire popcount27_xcpf_core_143;
  wire popcount27_xcpf_core_144;
  wire popcount27_xcpf_core_146;
  wire popcount27_xcpf_core_148;
  wire popcount27_xcpf_core_150;
  wire popcount27_xcpf_core_152;
  wire popcount27_xcpf_core_153;
  wire popcount27_xcpf_core_155;
  wire popcount27_xcpf_core_156;
  wire popcount27_xcpf_core_157;
  wire popcount27_xcpf_core_158;
  wire popcount27_xcpf_core_161;
  wire popcount27_xcpf_core_162;
  wire popcount27_xcpf_core_163;
  wire popcount27_xcpf_core_165;
  wire popcount27_xcpf_core_168;
  wire popcount27_xcpf_core_169;
  wire popcount27_xcpf_core_171;
  wire popcount27_xcpf_core_173;
  wire popcount27_xcpf_core_175;
  wire popcount27_xcpf_core_177;
  wire popcount27_xcpf_core_178;
  wire popcount27_xcpf_core_179;
  wire popcount27_xcpf_core_181;
  wire popcount27_xcpf_core_182;
  wire popcount27_xcpf_core_184;
  wire popcount27_xcpf_core_185;
  wire popcount27_xcpf_core_186;
  wire popcount27_xcpf_core_190;
  wire popcount27_xcpf_core_191;
  wire popcount27_xcpf_core_193;
  wire popcount27_xcpf_core_194;

  assign popcount27_xcpf_core_033 = ~(input_a[25] ^ input_a[9]);
  assign popcount27_xcpf_core_035 = input_a[3] | input_a[22];
  assign popcount27_xcpf_core_036 = ~(input_a[13] & input_a[15]);
  assign popcount27_xcpf_core_037 = ~(input_a[19] ^ input_a[9]);
  assign popcount27_xcpf_core_038 = ~(input_a[11] & input_a[24]);
  assign popcount27_xcpf_core_042 = input_a[20] ^ input_a[26];
  assign popcount27_xcpf_core_043 = ~input_a[12];
  assign popcount27_xcpf_core_044 = input_a[22] | input_a[11];
  assign popcount27_xcpf_core_045 = input_a[9] & input_a[0];
  assign popcount27_xcpf_core_046 = ~(input_a[23] & input_a[21]);
  assign popcount27_xcpf_core_047 = input_a[14] & input_a[17];
  assign popcount27_xcpf_core_048 = ~input_a[1];
  assign popcount27_xcpf_core_050 = input_a[16] ^ input_a[5];
  assign popcount27_xcpf_core_051 = ~(input_a[18] ^ input_a[9]);
  assign popcount27_xcpf_core_052 = ~input_a[5];
  assign popcount27_xcpf_core_056 = input_a[22] & input_a[0];
  assign popcount27_xcpf_core_057 = input_a[8] ^ input_a[14];
  assign popcount27_xcpf_core_058 = input_a[15] & input_a[16];
  assign popcount27_xcpf_core_059 = ~input_a[26];
  assign popcount27_xcpf_core_060 = ~(input_a[13] & input_a[19]);
  assign popcount27_xcpf_core_063 = ~input_a[22];
  assign popcount27_xcpf_core_064 = input_a[17] & input_a[2];
  assign popcount27_xcpf_core_065 = ~(input_a[12] ^ input_a[22]);
  assign popcount27_xcpf_core_066 = ~input_a[21];
  assign popcount27_xcpf_core_067 = ~(input_a[25] | input_a[26]);
  assign popcount27_xcpf_core_068 = input_a[9] & input_a[7];
  assign popcount27_xcpf_core_069 = ~(input_a[8] | input_a[18]);
  assign popcount27_xcpf_core_072 = ~(input_a[20] & input_a[16]);
  assign popcount27_xcpf_core_076 = ~input_a[0];
  assign popcount27_xcpf_core_077 = input_a[12] | input_a[12];
  assign popcount27_xcpf_core_078 = input_a[19] | input_a[7];
  assign popcount27_xcpf_core_079 = input_a[8] ^ input_a[13];
  assign popcount27_xcpf_core_080 = input_a[7] ^ input_a[12];
  assign popcount27_xcpf_core_082 = ~input_a[19];
  assign popcount27_xcpf_core_084 = ~(input_a[11] & input_a[24]);
  assign popcount27_xcpf_core_087 = input_a[20] ^ input_a[5];
  assign popcount27_xcpf_core_088 = ~input_a[16];
  assign popcount27_xcpf_core_091 = input_a[4] | input_a[15];
  assign popcount27_xcpf_core_092 = ~input_a[7];
  assign popcount27_xcpf_core_094 = ~(input_a[0] & input_a[7]);
  assign popcount27_xcpf_core_095_not = ~input_a[25];
  assign popcount27_xcpf_core_099 = input_a[11] | input_a[9];
  assign popcount27_xcpf_core_102 = input_a[0] & input_a[5];
  assign popcount27_xcpf_core_103 = ~(input_a[15] & input_a[2]);
  assign popcount27_xcpf_core_104 = ~(input_a[26] | input_a[16]);
  assign popcount27_xcpf_core_108 = input_a[19] ^ input_a[21];
  assign popcount27_xcpf_core_109 = input_a[24] & input_a[15];
  assign popcount27_xcpf_core_110 = ~(input_a[16] & input_a[14]);
  assign popcount27_xcpf_core_111 = input_a[5] | input_a[25];
  assign popcount27_xcpf_core_113 = ~(input_a[6] & input_a[13]);
  assign popcount27_xcpf_core_114 = input_a[2] | input_a[3];
  assign popcount27_xcpf_core_115 = ~input_a[0];
  assign popcount27_xcpf_core_116 = input_a[17] ^ input_a[17];
  assign popcount27_xcpf_core_117 = input_a[26] | input_a[6];
  assign popcount27_xcpf_core_119 = ~(input_a[26] ^ input_a[13]);
  assign popcount27_xcpf_core_120 = input_a[21] & input_a[26];
  assign popcount27_xcpf_core_122 = ~input_a[13];
  assign popcount27_xcpf_core_125 = input_a[20] ^ input_a[2];
  assign popcount27_xcpf_core_126 = ~(input_a[16] | input_a[11]);
  assign popcount27_xcpf_core_129 = ~input_a[18];
  assign popcount27_xcpf_core_130 = ~(input_a[15] | input_a[11]);
  assign popcount27_xcpf_core_131 = input_a[13] | input_a[7];
  assign popcount27_xcpf_core_133 = ~(input_a[2] & input_a[25]);
  assign popcount27_xcpf_core_135 = ~(input_a[1] | input_a[1]);
  assign popcount27_xcpf_core_136 = input_a[5] | input_a[24];
  assign popcount27_xcpf_core_137 = ~(input_a[7] | input_a[24]);
  assign popcount27_xcpf_core_138 = ~input_a[16];
  assign popcount27_xcpf_core_139 = ~(input_a[16] ^ input_a[9]);
  assign popcount27_xcpf_core_140 = ~(input_a[7] | input_a[12]);
  assign popcount27_xcpf_core_141 = input_a[25] ^ input_a[2];
  assign popcount27_xcpf_core_143 = ~input_a[25];
  assign popcount27_xcpf_core_144 = ~(input_a[11] ^ input_a[21]);
  assign popcount27_xcpf_core_146 = input_a[18] ^ input_a[19];
  assign popcount27_xcpf_core_148 = ~(input_a[26] ^ input_a[1]);
  assign popcount27_xcpf_core_150 = ~(input_a[8] & input_a[11]);
  assign popcount27_xcpf_core_152 = ~input_a[24];
  assign popcount27_xcpf_core_153 = ~(input_a[16] ^ input_a[3]);
  assign popcount27_xcpf_core_155 = input_a[14] | input_a[19];
  assign popcount27_xcpf_core_156 = ~(input_a[4] | input_a[23]);
  assign popcount27_xcpf_core_157 = ~(input_a[2] & input_a[21]);
  assign popcount27_xcpf_core_158 = ~(input_a[17] ^ input_a[5]);
  assign popcount27_xcpf_core_161 = ~(input_a[8] ^ input_a[15]);
  assign popcount27_xcpf_core_162 = ~(input_a[6] | input_a[21]);
  assign popcount27_xcpf_core_163 = input_a[18] | input_a[15];
  assign popcount27_xcpf_core_165 = input_a[20] & input_a[1];
  assign popcount27_xcpf_core_168 = ~(input_a[5] & input_a[25]);
  assign popcount27_xcpf_core_169 = input_a[20] & input_a[1];
  assign popcount27_xcpf_core_171 = input_a[9] ^ input_a[1];
  assign popcount27_xcpf_core_173 = ~(input_a[18] ^ input_a[7]);
  assign popcount27_xcpf_core_175 = input_a[25] ^ input_a[16];
  assign popcount27_xcpf_core_177 = ~(input_a[19] | input_a[1]);
  assign popcount27_xcpf_core_178 = input_a[26] & input_a[8];
  assign popcount27_xcpf_core_179 = input_a[6] & input_a[0];
  assign popcount27_xcpf_core_181 = ~(input_a[14] | input_a[23]);
  assign popcount27_xcpf_core_182 = ~(input_a[12] | input_a[23]);
  assign popcount27_xcpf_core_184 = ~(input_a[14] | input_a[21]);
  assign popcount27_xcpf_core_185 = ~(input_a[8] ^ input_a[19]);
  assign popcount27_xcpf_core_186 = ~(input_a[23] ^ input_a[18]);
  assign popcount27_xcpf_core_190 = input_a[7] ^ input_a[2];
  assign popcount27_xcpf_core_191 = input_a[20] & input_a[15];
  assign popcount27_xcpf_core_193 = ~(input_a[8] & input_a[11]);
  assign popcount27_xcpf_core_194 = ~(input_a[24] | input_a[4]);

  assign popcount27_xcpf_out[0] = input_a[1];
  assign popcount27_xcpf_out[1] = input_a[0];
  assign popcount27_xcpf_out[2] = 1'b1;
  assign popcount27_xcpf_out[3] = 1'b1;
  assign popcount27_xcpf_out[4] = 1'b0;
endmodule