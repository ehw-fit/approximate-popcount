// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.54316
// WCE=12.0
// EP=0.797723%
// Printed PDK parameters:
//  Area=42263464.0
//  Delay=53974876.0
//  Power=1863400.0

module popcount31_efxp(input [30:0] input_a, output [4:0] popcount31_efxp_out);
  wire popcount31_efxp_core_035;
  wire popcount31_efxp_core_036;
  wire popcount31_efxp_core_037;
  wire popcount31_efxp_core_039;
  wire popcount31_efxp_core_040;
  wire popcount31_efxp_core_042;
  wire popcount31_efxp_core_043;
  wire popcount31_efxp_core_044;
  wire popcount31_efxp_core_045;
  wire popcount31_efxp_core_046_not;
  wire popcount31_efxp_core_047;
  wire popcount31_efxp_core_048;
  wire popcount31_efxp_core_049;
  wire popcount31_efxp_core_051;
  wire popcount31_efxp_core_052;
  wire popcount31_efxp_core_053;
  wire popcount31_efxp_core_056;
  wire popcount31_efxp_core_057;
  wire popcount31_efxp_core_061;
  wire popcount31_efxp_core_062;
  wire popcount31_efxp_core_063;
  wire popcount31_efxp_core_064;
  wire popcount31_efxp_core_065;
  wire popcount31_efxp_core_067;
  wire popcount31_efxp_core_068;
  wire popcount31_efxp_core_069;
  wire popcount31_efxp_core_070;
  wire popcount31_efxp_core_071;
  wire popcount31_efxp_core_072;
  wire popcount31_efxp_core_073;
  wire popcount31_efxp_core_074;
  wire popcount31_efxp_core_076;
  wire popcount31_efxp_core_078;
  wire popcount31_efxp_core_079;
  wire popcount31_efxp_core_081;
  wire popcount31_efxp_core_083;
  wire popcount31_efxp_core_084;
  wire popcount31_efxp_core_085;
  wire popcount31_efxp_core_086;
  wire popcount31_efxp_core_087;
  wire popcount31_efxp_core_089;
  wire popcount31_efxp_core_092;
  wire popcount31_efxp_core_093;
  wire popcount31_efxp_core_095;
  wire popcount31_efxp_core_096;
  wire popcount31_efxp_core_098;
  wire popcount31_efxp_core_099;
  wire popcount31_efxp_core_101;
  wire popcount31_efxp_core_103;
  wire popcount31_efxp_core_104;
  wire popcount31_efxp_core_105;
  wire popcount31_efxp_core_106;
  wire popcount31_efxp_core_107;
  wire popcount31_efxp_core_109;
  wire popcount31_efxp_core_112;
  wire popcount31_efxp_core_113;
  wire popcount31_efxp_core_114;
  wire popcount31_efxp_core_116;
  wire popcount31_efxp_core_117;
  wire popcount31_efxp_core_118;
  wire popcount31_efxp_core_120;
  wire popcount31_efxp_core_121;
  wire popcount31_efxp_core_122;
  wire popcount31_efxp_core_123;
  wire popcount31_efxp_core_124;
  wire popcount31_efxp_core_125;
  wire popcount31_efxp_core_127;
  wire popcount31_efxp_core_129;
  wire popcount31_efxp_core_130;
  wire popcount31_efxp_core_131;
  wire popcount31_efxp_core_132;
  wire popcount31_efxp_core_135;
  wire popcount31_efxp_core_137;
  wire popcount31_efxp_core_138;
  wire popcount31_efxp_core_140;
  wire popcount31_efxp_core_143;
  wire popcount31_efxp_core_145;
  wire popcount31_efxp_core_147;
  wire popcount31_efxp_core_148;
  wire popcount31_efxp_core_149;
  wire popcount31_efxp_core_150;
  wire popcount31_efxp_core_151;
  wire popcount31_efxp_core_152;
  wire popcount31_efxp_core_153;
  wire popcount31_efxp_core_154;
  wire popcount31_efxp_core_155;
  wire popcount31_efxp_core_158;
  wire popcount31_efxp_core_159;
  wire popcount31_efxp_core_160;
  wire popcount31_efxp_core_161;
  wire popcount31_efxp_core_162;
  wire popcount31_efxp_core_163;
  wire popcount31_efxp_core_164;
  wire popcount31_efxp_core_165;
  wire popcount31_efxp_core_166;
  wire popcount31_efxp_core_167;
  wire popcount31_efxp_core_169;
  wire popcount31_efxp_core_170;
  wire popcount31_efxp_core_171;
  wire popcount31_efxp_core_172;
  wire popcount31_efxp_core_173;
  wire popcount31_efxp_core_174;
  wire popcount31_efxp_core_175;
  wire popcount31_efxp_core_176;
  wire popcount31_efxp_core_177;
  wire popcount31_efxp_core_178;
  wire popcount31_efxp_core_179;
  wire popcount31_efxp_core_181;
  wire popcount31_efxp_core_182;
  wire popcount31_efxp_core_183;
  wire popcount31_efxp_core_184;
  wire popcount31_efxp_core_186;
  wire popcount31_efxp_core_188;
  wire popcount31_efxp_core_189;
  wire popcount31_efxp_core_190;
  wire popcount31_efxp_core_191;
  wire popcount31_efxp_core_192;
  wire popcount31_efxp_core_197;
  wire popcount31_efxp_core_199;
  wire popcount31_efxp_core_200;
  wire popcount31_efxp_core_202;
  wire popcount31_efxp_core_204;
  wire popcount31_efxp_core_205;
  wire popcount31_efxp_core_206;
  wire popcount31_efxp_core_207;
  wire popcount31_efxp_core_208;
  wire popcount31_efxp_core_209;
  wire popcount31_efxp_core_210;
  wire popcount31_efxp_core_211;
  wire popcount31_efxp_core_212;
  wire popcount31_efxp_core_213;
  wire popcount31_efxp_core_214;
  wire popcount31_efxp_core_215;
  wire popcount31_efxp_core_216;
  wire popcount31_efxp_core_217;
  wire popcount31_efxp_core_218;
  wire popcount31_efxp_core_219;

  assign popcount31_efxp_core_035 = ~input_a[18];
  assign popcount31_efxp_core_036 = ~input_a[12];
  assign popcount31_efxp_core_037 = input_a[2] | input_a[13];
  assign popcount31_efxp_core_039 = input_a[16] ^ input_a[29];
  assign popcount31_efxp_core_040 = input_a[16] & input_a[14];
  assign popcount31_efxp_core_042 = input_a[12] & input_a[4];
  assign popcount31_efxp_core_043 = input_a[17] & input_a[30];
  assign popcount31_efxp_core_044 = ~input_a[20];
  assign popcount31_efxp_core_045 = popcount31_efxp_core_040 | popcount31_efxp_core_042;
  assign popcount31_efxp_core_046_not = ~input_a[3];
  assign popcount31_efxp_core_047 = ~(popcount31_efxp_core_045 & input_a[18]);
  assign popcount31_efxp_core_048 = popcount31_efxp_core_045 & input_a[18];
  assign popcount31_efxp_core_049 = input_a[13] | popcount31_efxp_core_048;
  assign popcount31_efxp_core_051 = input_a[15] & input_a[26];
  assign popcount31_efxp_core_052 = popcount31_efxp_core_037 ^ popcount31_efxp_core_047;
  assign popcount31_efxp_core_053 = ~(input_a[12] & input_a[1]);
  assign popcount31_efxp_core_056 = ~input_a[22];
  assign popcount31_efxp_core_057 = input_a[2] | popcount31_efxp_core_049;
  assign popcount31_efxp_core_061 = ~(input_a[6] ^ input_a[6]);
  assign popcount31_efxp_core_062 = input_a[12] & input_a[22];
  assign popcount31_efxp_core_063 = input_a[8] & input_a[5];
  assign popcount31_efxp_core_064 = input_a[9] ^ input_a[10];
  assign popcount31_efxp_core_065 = input_a[9] & input_a[10];
  assign popcount31_efxp_core_067 = input_a[7] & popcount31_efxp_core_064;
  assign popcount31_efxp_core_068 = popcount31_efxp_core_063 ^ popcount31_efxp_core_065;
  assign popcount31_efxp_core_069 = popcount31_efxp_core_063 & input_a[10];
  assign popcount31_efxp_core_070 = popcount31_efxp_core_068 ^ popcount31_efxp_core_067;
  assign popcount31_efxp_core_071 = popcount31_efxp_core_068 & popcount31_efxp_core_067;
  assign popcount31_efxp_core_072 = popcount31_efxp_core_069 | popcount31_efxp_core_071;
  assign popcount31_efxp_core_073 = input_a[18] & input_a[22];
  assign popcount31_efxp_core_074 = input_a[1] & input_a[3];
  assign popcount31_efxp_core_076 = input_a[20] & input_a[6];
  assign popcount31_efxp_core_078 = input_a[22] & input_a[21];
  assign popcount31_efxp_core_079 = popcount31_efxp_core_074 | popcount31_efxp_core_076;
  assign popcount31_efxp_core_081 = popcount31_efxp_core_079 | popcount31_efxp_core_078;
  assign popcount31_efxp_core_083 = ~(input_a[4] ^ input_a[27]);
  assign popcount31_efxp_core_084 = ~(input_a[8] | input_a[0]);
  assign popcount31_efxp_core_085 = ~input_a[15];
  assign popcount31_efxp_core_086 = popcount31_efxp_core_070 ^ popcount31_efxp_core_081;
  assign popcount31_efxp_core_087 = popcount31_efxp_core_070 & popcount31_efxp_core_081;
  assign popcount31_efxp_core_089 = input_a[2] ^ input_a[19];
  assign popcount31_efxp_core_092 = input_a[7] | input_a[9];
  assign popcount31_efxp_core_093 = popcount31_efxp_core_072 | popcount31_efxp_core_087;
  assign popcount31_efxp_core_095 = ~input_a[20];
  assign popcount31_efxp_core_096 = input_a[9] | input_a[30];
  assign popcount31_efxp_core_098 = popcount31_efxp_core_052 ^ popcount31_efxp_core_086;
  assign popcount31_efxp_core_099 = popcount31_efxp_core_052 & popcount31_efxp_core_086;
  assign popcount31_efxp_core_101 = ~input_a[15];
  assign popcount31_efxp_core_103 = popcount31_efxp_core_057 ^ popcount31_efxp_core_093;
  assign popcount31_efxp_core_104 = popcount31_efxp_core_057 & popcount31_efxp_core_093;
  assign popcount31_efxp_core_105 = popcount31_efxp_core_103 ^ popcount31_efxp_core_099;
  assign popcount31_efxp_core_106 = popcount31_efxp_core_103 & popcount31_efxp_core_099;
  assign popcount31_efxp_core_107 = popcount31_efxp_core_104 | popcount31_efxp_core_106;
  assign popcount31_efxp_core_109 = ~(input_a[2] ^ input_a[3]);
  assign popcount31_efxp_core_112 = ~(input_a[6] ^ input_a[12]);
  assign popcount31_efxp_core_113 = ~(input_a[10] & input_a[13]);
  assign popcount31_efxp_core_114 = ~(input_a[6] ^ input_a[23]);
  assign popcount31_efxp_core_116 = ~(input_a[20] & input_a[24]);
  assign popcount31_efxp_core_117 = input_a[30] & input_a[17];
  assign popcount31_efxp_core_118 = input_a[18] & input_a[19];
  assign popcount31_efxp_core_120 = ~(input_a[3] & input_a[21]);
  assign popcount31_efxp_core_121 = input_a[23] ^ input_a[19];
  assign popcount31_efxp_core_122 = ~(input_a[12] | input_a[30]);
  assign popcount31_efxp_core_123 = input_a[6] | input_a[14];
  assign popcount31_efxp_core_124 = input_a[1] ^ input_a[7];
  assign popcount31_efxp_core_125 = ~(input_a[27] ^ input_a[18]);
  assign popcount31_efxp_core_127 = input_a[29] | input_a[24];
  assign popcount31_efxp_core_129 = input_a[28] ^ input_a[22];
  assign popcount31_efxp_core_130 = ~(input_a[3] | input_a[3]);
  assign popcount31_efxp_core_131 = input_a[28] ^ input_a[12];
  assign popcount31_efxp_core_132 = input_a[29] ^ input_a[5];
  assign popcount31_efxp_core_135 = ~(input_a[23] ^ input_a[2]);
  assign popcount31_efxp_core_137 = ~(input_a[15] & input_a[17]);
  assign popcount31_efxp_core_138 = input_a[15] & input_a[17];
  assign popcount31_efxp_core_140 = input_a[4] ^ input_a[11];
  assign popcount31_efxp_core_143 = ~(input_a[30] & input_a[21]);
  assign popcount31_efxp_core_145 = input_a[20] | input_a[10];
  assign popcount31_efxp_core_147 = ~(input_a[23] & input_a[24]);
  assign popcount31_efxp_core_148 = input_a[23] & input_a[24];
  assign popcount31_efxp_core_149 = input_a[25] ^ input_a[26];
  assign popcount31_efxp_core_150 = input_a[25] & input_a[26];
  assign popcount31_efxp_core_151 = popcount31_efxp_core_147 ^ popcount31_efxp_core_149;
  assign popcount31_efxp_core_152 = popcount31_efxp_core_147 & popcount31_efxp_core_149;
  assign popcount31_efxp_core_153 = popcount31_efxp_core_148 ^ popcount31_efxp_core_150;
  assign popcount31_efxp_core_154 = input_a[25] & input_a[26];
  assign popcount31_efxp_core_155 = popcount31_efxp_core_153 | popcount31_efxp_core_152;
  assign popcount31_efxp_core_158 = ~(input_a[27] & input_a[28]);
  assign popcount31_efxp_core_159 = input_a[27] & input_a[28];
  assign popcount31_efxp_core_160 = input_a[29] ^ input_a[30];
  assign popcount31_efxp_core_161 = input_a[29] & input_a[30];
  assign popcount31_efxp_core_162 = popcount31_efxp_core_158 ^ popcount31_efxp_core_160;
  assign popcount31_efxp_core_163 = popcount31_efxp_core_158 & popcount31_efxp_core_160;
  assign popcount31_efxp_core_164 = popcount31_efxp_core_159 ^ popcount31_efxp_core_161;
  assign popcount31_efxp_core_165 = input_a[29] & input_a[30];
  assign popcount31_efxp_core_166 = popcount31_efxp_core_164 | popcount31_efxp_core_163;
  assign popcount31_efxp_core_167 = ~(input_a[10] ^ input_a[25]);
  assign popcount31_efxp_core_169 = input_a[29] & input_a[13];
  assign popcount31_efxp_core_170 = popcount31_efxp_core_151 & popcount31_efxp_core_162;
  assign popcount31_efxp_core_171 = popcount31_efxp_core_155 ^ popcount31_efxp_core_166;
  assign popcount31_efxp_core_172 = popcount31_efxp_core_155 & popcount31_efxp_core_166;
  assign popcount31_efxp_core_173 = popcount31_efxp_core_171 ^ popcount31_efxp_core_170;
  assign popcount31_efxp_core_174 = popcount31_efxp_core_171 & popcount31_efxp_core_170;
  assign popcount31_efxp_core_175 = popcount31_efxp_core_172 | popcount31_efxp_core_174;
  assign popcount31_efxp_core_176 = popcount31_efxp_core_154 | popcount31_efxp_core_165;
  assign popcount31_efxp_core_177 = ~(input_a[22] ^ input_a[4]);
  assign popcount31_efxp_core_178 = popcount31_efxp_core_176 | popcount31_efxp_core_175;
  assign popcount31_efxp_core_179 = ~(input_a[5] & input_a[23]);
  assign popcount31_efxp_core_181 = ~(input_a[18] & input_a[30]);
  assign popcount31_efxp_core_182 = ~(input_a[28] | input_a[10]);
  assign popcount31_efxp_core_183 = popcount31_efxp_core_137 ^ popcount31_efxp_core_173;
  assign popcount31_efxp_core_184 = popcount31_efxp_core_137 & popcount31_efxp_core_173;
  assign popcount31_efxp_core_186 = ~(input_a[14] | input_a[1]);
  assign popcount31_efxp_core_188 = popcount31_efxp_core_138 ^ popcount31_efxp_core_178;
  assign popcount31_efxp_core_189 = popcount31_efxp_core_138 & popcount31_efxp_core_178;
  assign popcount31_efxp_core_190 = popcount31_efxp_core_188 ^ popcount31_efxp_core_184;
  assign popcount31_efxp_core_191 = popcount31_efxp_core_188 & popcount31_efxp_core_184;
  assign popcount31_efxp_core_192 = popcount31_efxp_core_189 | popcount31_efxp_core_191;
  assign popcount31_efxp_core_197 = ~(input_a[26] ^ input_a[12]);
  assign popcount31_efxp_core_199 = ~(input_a[13] ^ input_a[8]);
  assign popcount31_efxp_core_200 = popcount31_efxp_core_098 ^ popcount31_efxp_core_183;
  assign popcount31_efxp_core_202 = ~popcount31_efxp_core_200;
  assign popcount31_efxp_core_204 = popcount31_efxp_core_098 | popcount31_efxp_core_200;
  assign popcount31_efxp_core_205 = popcount31_efxp_core_105 ^ popcount31_efxp_core_190;
  assign popcount31_efxp_core_206 = popcount31_efxp_core_105 & popcount31_efxp_core_190;
  assign popcount31_efxp_core_207 = popcount31_efxp_core_205 ^ popcount31_efxp_core_204;
  assign popcount31_efxp_core_208 = popcount31_efxp_core_205 & popcount31_efxp_core_204;
  assign popcount31_efxp_core_209 = popcount31_efxp_core_206 | popcount31_efxp_core_208;
  assign popcount31_efxp_core_210 = popcount31_efxp_core_107 ^ popcount31_efxp_core_192;
  assign popcount31_efxp_core_211 = popcount31_efxp_core_107 & popcount31_efxp_core_192;
  assign popcount31_efxp_core_212 = popcount31_efxp_core_210 ^ popcount31_efxp_core_209;
  assign popcount31_efxp_core_213 = popcount31_efxp_core_210 & popcount31_efxp_core_209;
  assign popcount31_efxp_core_214 = popcount31_efxp_core_211 | popcount31_efxp_core_213;
  assign popcount31_efxp_core_215 = input_a[22] & input_a[15];
  assign popcount31_efxp_core_216 = ~input_a[2];
  assign popcount31_efxp_core_217 = input_a[5] & input_a[7];
  assign popcount31_efxp_core_218 = ~(input_a[5] | input_a[6]);
  assign popcount31_efxp_core_219 = ~input_a[9];

  assign popcount31_efxp_out[0] = input_a[19];
  assign popcount31_efxp_out[1] = popcount31_efxp_core_202;
  assign popcount31_efxp_out[2] = popcount31_efxp_core_207;
  assign popcount31_efxp_out[3] = popcount31_efxp_core_212;
  assign popcount31_efxp_out[4] = popcount31_efxp_core_214;
endmodule