// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.02833
// WCE=27.0
// EP=0.948206%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_w9zx(input [35:0] input_a, output [5:0] popcount36_w9zx_out);
  wire popcount36_w9zx_core_038;
  wire popcount36_w9zx_core_040;
  wire popcount36_w9zx_core_042;
  wire popcount36_w9zx_core_043;
  wire popcount36_w9zx_core_044;
  wire popcount36_w9zx_core_047;
  wire popcount36_w9zx_core_048;
  wire popcount36_w9zx_core_049;
  wire popcount36_w9zx_core_050;
  wire popcount36_w9zx_core_051;
  wire popcount36_w9zx_core_052;
  wire popcount36_w9zx_core_053;
  wire popcount36_w9zx_core_056;
  wire popcount36_w9zx_core_057;
  wire popcount36_w9zx_core_058;
  wire popcount36_w9zx_core_059;
  wire popcount36_w9zx_core_060;
  wire popcount36_w9zx_core_062;
  wire popcount36_w9zx_core_063;
  wire popcount36_w9zx_core_064;
  wire popcount36_w9zx_core_066;
  wire popcount36_w9zx_core_067_not;
  wire popcount36_w9zx_core_069;
  wire popcount36_w9zx_core_070;
  wire popcount36_w9zx_core_072;
  wire popcount36_w9zx_core_073;
  wire popcount36_w9zx_core_074;
  wire popcount36_w9zx_core_076;
  wire popcount36_w9zx_core_077;
  wire popcount36_w9zx_core_078;
  wire popcount36_w9zx_core_079;
  wire popcount36_w9zx_core_082_not;
  wire popcount36_w9zx_core_083;
  wire popcount36_w9zx_core_084;
  wire popcount36_w9zx_core_086;
  wire popcount36_w9zx_core_087;
  wire popcount36_w9zx_core_088;
  wire popcount36_w9zx_core_089_not;
  wire popcount36_w9zx_core_090;
  wire popcount36_w9zx_core_093;
  wire popcount36_w9zx_core_094;
  wire popcount36_w9zx_core_095;
  wire popcount36_w9zx_core_098;
  wire popcount36_w9zx_core_100;
  wire popcount36_w9zx_core_102;
  wire popcount36_w9zx_core_103;
  wire popcount36_w9zx_core_104;
  wire popcount36_w9zx_core_106;
  wire popcount36_w9zx_core_110_not;
  wire popcount36_w9zx_core_112;
  wire popcount36_w9zx_core_113;
  wire popcount36_w9zx_core_114;
  wire popcount36_w9zx_core_118;
  wire popcount36_w9zx_core_120;
  wire popcount36_w9zx_core_121;
  wire popcount36_w9zx_core_122;
  wire popcount36_w9zx_core_123;
  wire popcount36_w9zx_core_124;
  wire popcount36_w9zx_core_126;
  wire popcount36_w9zx_core_127;
  wire popcount36_w9zx_core_128;
  wire popcount36_w9zx_core_129;
  wire popcount36_w9zx_core_130;
  wire popcount36_w9zx_core_132;
  wire popcount36_w9zx_core_133_not;
  wire popcount36_w9zx_core_134;
  wire popcount36_w9zx_core_135;
  wire popcount36_w9zx_core_136;
  wire popcount36_w9zx_core_137;
  wire popcount36_w9zx_core_138;
  wire popcount36_w9zx_core_139;
  wire popcount36_w9zx_core_140;
  wire popcount36_w9zx_core_141;
  wire popcount36_w9zx_core_142;
  wire popcount36_w9zx_core_144;
  wire popcount36_w9zx_core_146;
  wire popcount36_w9zx_core_151;
  wire popcount36_w9zx_core_152;
  wire popcount36_w9zx_core_154;
  wire popcount36_w9zx_core_155;
  wire popcount36_w9zx_core_157;
  wire popcount36_w9zx_core_159;
  wire popcount36_w9zx_core_160;
  wire popcount36_w9zx_core_161;
  wire popcount36_w9zx_core_162;
  wire popcount36_w9zx_core_163;
  wire popcount36_w9zx_core_164;
  wire popcount36_w9zx_core_165;
  wire popcount36_w9zx_core_166;
  wire popcount36_w9zx_core_167;
  wire popcount36_w9zx_core_168;
  wire popcount36_w9zx_core_169;
  wire popcount36_w9zx_core_170;
  wire popcount36_w9zx_core_172;
  wire popcount36_w9zx_core_173;
  wire popcount36_w9zx_core_174;
  wire popcount36_w9zx_core_175;
  wire popcount36_w9zx_core_178;
  wire popcount36_w9zx_core_180;
  wire popcount36_w9zx_core_181;
  wire popcount36_w9zx_core_183;
  wire popcount36_w9zx_core_185;
  wire popcount36_w9zx_core_186;
  wire popcount36_w9zx_core_187;
  wire popcount36_w9zx_core_188;
  wire popcount36_w9zx_core_189;
  wire popcount36_w9zx_core_190;
  wire popcount36_w9zx_core_191;
  wire popcount36_w9zx_core_192;
  wire popcount36_w9zx_core_193;
  wire popcount36_w9zx_core_194;
  wire popcount36_w9zx_core_196;
  wire popcount36_w9zx_core_199;
  wire popcount36_w9zx_core_201;
  wire popcount36_w9zx_core_202;
  wire popcount36_w9zx_core_203;
  wire popcount36_w9zx_core_204;
  wire popcount36_w9zx_core_205;
  wire popcount36_w9zx_core_207;
  wire popcount36_w9zx_core_209;
  wire popcount36_w9zx_core_210_not;
  wire popcount36_w9zx_core_211;
  wire popcount36_w9zx_core_213;
  wire popcount36_w9zx_core_214;
  wire popcount36_w9zx_core_215;
  wire popcount36_w9zx_core_216;
  wire popcount36_w9zx_core_218;
  wire popcount36_w9zx_core_220;
  wire popcount36_w9zx_core_222;
  wire popcount36_w9zx_core_223;
  wire popcount36_w9zx_core_224;
  wire popcount36_w9zx_core_225;
  wire popcount36_w9zx_core_227;
  wire popcount36_w9zx_core_235;
  wire popcount36_w9zx_core_236;
  wire popcount36_w9zx_core_237;
  wire popcount36_w9zx_core_238;
  wire popcount36_w9zx_core_240;
  wire popcount36_w9zx_core_242;
  wire popcount36_w9zx_core_243;
  wire popcount36_w9zx_core_244;
  wire popcount36_w9zx_core_245;
  wire popcount36_w9zx_core_246;
  wire popcount36_w9zx_core_247;
  wire popcount36_w9zx_core_248;
  wire popcount36_w9zx_core_249;
  wire popcount36_w9zx_core_251;
  wire popcount36_w9zx_core_252;
  wire popcount36_w9zx_core_254;
  wire popcount36_w9zx_core_255;
  wire popcount36_w9zx_core_258;
  wire popcount36_w9zx_core_259;
  wire popcount36_w9zx_core_260;
  wire popcount36_w9zx_core_261;
  wire popcount36_w9zx_core_262;
  wire popcount36_w9zx_core_263;
  wire popcount36_w9zx_core_264;
  wire popcount36_w9zx_core_266;
  wire popcount36_w9zx_core_267;
  wire popcount36_w9zx_core_268;
  wire popcount36_w9zx_core_269;
  wire popcount36_w9zx_core_271;
  wire popcount36_w9zx_core_272;
  wire popcount36_w9zx_core_274;
  wire popcount36_w9zx_core_275;

  assign popcount36_w9zx_core_038 = ~(input_a[4] | input_a[15]);
  assign popcount36_w9zx_core_040 = ~(input_a[30] | input_a[16]);
  assign popcount36_w9zx_core_042 = ~(input_a[6] | input_a[18]);
  assign popcount36_w9zx_core_043 = input_a[24] | input_a[5];
  assign popcount36_w9zx_core_044 = ~input_a[34];
  assign popcount36_w9zx_core_047 = ~(input_a[21] ^ input_a[8]);
  assign popcount36_w9zx_core_048 = input_a[2] & input_a[10];
  assign popcount36_w9zx_core_049 = ~(input_a[30] | input_a[17]);
  assign popcount36_w9zx_core_050 = input_a[3] & input_a[23];
  assign popcount36_w9zx_core_051 = ~(input_a[25] ^ input_a[3]);
  assign popcount36_w9zx_core_052 = input_a[15] & input_a[14];
  assign popcount36_w9zx_core_053 = input_a[19] & input_a[9];
  assign popcount36_w9zx_core_056 = ~input_a[16];
  assign popcount36_w9zx_core_057 = ~(input_a[6] | input_a[22]);
  assign popcount36_w9zx_core_058 = input_a[17] & input_a[22];
  assign popcount36_w9zx_core_059 = input_a[31] | input_a[5];
  assign popcount36_w9zx_core_060 = ~(input_a[31] | input_a[12]);
  assign popcount36_w9zx_core_062 = ~(input_a[23] ^ input_a[8]);
  assign popcount36_w9zx_core_063 = ~(input_a[9] | input_a[31]);
  assign popcount36_w9zx_core_064 = ~(input_a[31] | input_a[25]);
  assign popcount36_w9zx_core_066 = input_a[0] ^ input_a[1];
  assign popcount36_w9zx_core_067_not = ~input_a[30];
  assign popcount36_w9zx_core_069 = ~(input_a[12] & input_a[0]);
  assign popcount36_w9zx_core_070 = input_a[4] ^ input_a[31];
  assign popcount36_w9zx_core_072 = ~input_a[15];
  assign popcount36_w9zx_core_073 = input_a[25] & input_a[20];
  assign popcount36_w9zx_core_074 = input_a[21] & input_a[13];
  assign popcount36_w9zx_core_076 = input_a[6] & input_a[30];
  assign popcount36_w9zx_core_077 = ~(input_a[11] ^ input_a[4]);
  assign popcount36_w9zx_core_078 = input_a[13] ^ input_a[5];
  assign popcount36_w9zx_core_079 = ~(input_a[0] & input_a[6]);
  assign popcount36_w9zx_core_082_not = ~input_a[4];
  assign popcount36_w9zx_core_083 = ~(input_a[24] & input_a[24]);
  assign popcount36_w9zx_core_084 = input_a[0] | input_a[30];
  assign popcount36_w9zx_core_086 = input_a[0] ^ input_a[18];
  assign popcount36_w9zx_core_087 = ~input_a[34];
  assign popcount36_w9zx_core_088 = ~(input_a[16] ^ input_a[34]);
  assign popcount36_w9zx_core_089_not = ~input_a[3];
  assign popcount36_w9zx_core_090 = input_a[3] & input_a[0];
  assign popcount36_w9zx_core_093 = input_a[14] | input_a[8];
  assign popcount36_w9zx_core_094 = input_a[9] | input_a[11];
  assign popcount36_w9zx_core_095 = ~(input_a[12] | input_a[0]);
  assign popcount36_w9zx_core_098 = ~(input_a[16] & input_a[3]);
  assign popcount36_w9zx_core_100 = ~(input_a[32] | input_a[4]);
  assign popcount36_w9zx_core_102 = ~(input_a[0] | input_a[20]);
  assign popcount36_w9zx_core_103 = ~input_a[18];
  assign popcount36_w9zx_core_104 = ~input_a[3];
  assign popcount36_w9zx_core_106 = ~(input_a[18] | input_a[11]);
  assign popcount36_w9zx_core_110_not = ~input_a[31];
  assign popcount36_w9zx_core_112 = input_a[4] ^ input_a[29];
  assign popcount36_w9zx_core_113 = ~(input_a[9] & input_a[11]);
  assign popcount36_w9zx_core_114 = input_a[25] ^ input_a[3];
  assign popcount36_w9zx_core_118 = input_a[33] ^ input_a[18];
  assign popcount36_w9zx_core_120 = ~(input_a[14] ^ input_a[33]);
  assign popcount36_w9zx_core_121 = ~input_a[5];
  assign popcount36_w9zx_core_122 = input_a[31] & input_a[28];
  assign popcount36_w9zx_core_123 = ~input_a[24];
  assign popcount36_w9zx_core_124 = input_a[0] ^ input_a[7];
  assign popcount36_w9zx_core_126 = ~(input_a[25] & input_a[4]);
  assign popcount36_w9zx_core_127 = ~(input_a[18] ^ input_a[9]);
  assign popcount36_w9zx_core_128 = ~input_a[2];
  assign popcount36_w9zx_core_129 = ~(input_a[29] & input_a[2]);
  assign popcount36_w9zx_core_130 = input_a[6] ^ input_a[27];
  assign popcount36_w9zx_core_132 = ~input_a[9];
  assign popcount36_w9zx_core_133_not = ~input_a[16];
  assign popcount36_w9zx_core_134 = ~input_a[6];
  assign popcount36_w9zx_core_135 = ~input_a[25];
  assign popcount36_w9zx_core_136 = input_a[1] ^ input_a[35];
  assign popcount36_w9zx_core_137 = ~input_a[0];
  assign popcount36_w9zx_core_138 = ~(input_a[11] ^ input_a[22]);
  assign popcount36_w9zx_core_139 = input_a[18] | input_a[7];
  assign popcount36_w9zx_core_140 = ~(input_a[11] | input_a[2]);
  assign popcount36_w9zx_core_141 = input_a[8] | input_a[4];
  assign popcount36_w9zx_core_142 = input_a[16] | input_a[34];
  assign popcount36_w9zx_core_144 = ~(input_a[5] & input_a[8]);
  assign popcount36_w9zx_core_146 = input_a[22] ^ input_a[30];
  assign popcount36_w9zx_core_151 = input_a[10] & input_a[33];
  assign popcount36_w9zx_core_152 = input_a[8] | input_a[13];
  assign popcount36_w9zx_core_154 = ~(input_a[21] ^ input_a[26]);
  assign popcount36_w9zx_core_155 = ~(input_a[25] & input_a[21]);
  assign popcount36_w9zx_core_157 = ~input_a[30];
  assign popcount36_w9zx_core_159 = input_a[20] | input_a[7];
  assign popcount36_w9zx_core_160 = input_a[10] ^ input_a[28];
  assign popcount36_w9zx_core_161 = ~input_a[28];
  assign popcount36_w9zx_core_162 = ~(input_a[3] & input_a[15]);
  assign popcount36_w9zx_core_163 = input_a[6] & input_a[15];
  assign popcount36_w9zx_core_164 = ~input_a[5];
  assign popcount36_w9zx_core_165 = input_a[6] ^ input_a[17];
  assign popcount36_w9zx_core_166 = ~(input_a[11] & input_a[18]);
  assign popcount36_w9zx_core_167 = ~(input_a[31] ^ input_a[7]);
  assign popcount36_w9zx_core_168 = ~input_a[14];
  assign popcount36_w9zx_core_169 = ~(input_a[14] & input_a[19]);
  assign popcount36_w9zx_core_170 = input_a[24] | input_a[19];
  assign popcount36_w9zx_core_172 = ~(input_a[20] | input_a[21]);
  assign popcount36_w9zx_core_173 = ~input_a[22];
  assign popcount36_w9zx_core_174 = ~(input_a[28] ^ input_a[6]);
  assign popcount36_w9zx_core_175 = ~(input_a[9] ^ input_a[11]);
  assign popcount36_w9zx_core_178 = ~(input_a[6] ^ input_a[24]);
  assign popcount36_w9zx_core_180 = input_a[20] ^ input_a[35];
  assign popcount36_w9zx_core_181 = input_a[0] | input_a[4];
  assign popcount36_w9zx_core_183 = ~input_a[14];
  assign popcount36_w9zx_core_185 = input_a[10] & input_a[28];
  assign popcount36_w9zx_core_186 = input_a[35] | input_a[27];
  assign popcount36_w9zx_core_187 = ~input_a[33];
  assign popcount36_w9zx_core_188 = input_a[11] | input_a[21];
  assign popcount36_w9zx_core_189 = input_a[6] | input_a[28];
  assign popcount36_w9zx_core_190 = input_a[14] | input_a[12];
  assign popcount36_w9zx_core_191 = input_a[4] ^ input_a[34];
  assign popcount36_w9zx_core_192 = input_a[17] & input_a[20];
  assign popcount36_w9zx_core_193 = ~input_a[8];
  assign popcount36_w9zx_core_194 = input_a[35] | input_a[35];
  assign popcount36_w9zx_core_196 = input_a[28] & input_a[2];
  assign popcount36_w9zx_core_199 = input_a[7] & input_a[7];
  assign popcount36_w9zx_core_201 = input_a[19] ^ input_a[8];
  assign popcount36_w9zx_core_202 = ~(input_a[22] | input_a[21]);
  assign popcount36_w9zx_core_203 = input_a[17] | input_a[10];
  assign popcount36_w9zx_core_204 = input_a[26] | input_a[0];
  assign popcount36_w9zx_core_205 = input_a[6] & input_a[17];
  assign popcount36_w9zx_core_207 = ~(input_a[27] ^ input_a[12]);
  assign popcount36_w9zx_core_209 = ~(input_a[20] & input_a[18]);
  assign popcount36_w9zx_core_210_not = ~input_a[19];
  assign popcount36_w9zx_core_211 = ~(input_a[18] ^ input_a[16]);
  assign popcount36_w9zx_core_213 = ~(input_a[1] | input_a[18]);
  assign popcount36_w9zx_core_214 = ~(input_a[26] | input_a[30]);
  assign popcount36_w9zx_core_215 = input_a[12] & input_a[17];
  assign popcount36_w9zx_core_216 = input_a[5] & input_a[30];
  assign popcount36_w9zx_core_218 = ~input_a[13];
  assign popcount36_w9zx_core_220 = ~(input_a[5] & input_a[8]);
  assign popcount36_w9zx_core_222 = ~(input_a[21] & input_a[5]);
  assign popcount36_w9zx_core_223 = ~(input_a[34] & input_a[35]);
  assign popcount36_w9zx_core_224 = ~(input_a[12] ^ input_a[21]);
  assign popcount36_w9zx_core_225 = ~(input_a[24] & input_a[31]);
  assign popcount36_w9zx_core_227 = ~(input_a[19] ^ input_a[10]);
  assign popcount36_w9zx_core_235 = input_a[2] ^ input_a[18];
  assign popcount36_w9zx_core_236 = input_a[19] ^ input_a[32];
  assign popcount36_w9zx_core_237 = ~(input_a[18] & input_a[0]);
  assign popcount36_w9zx_core_238 = input_a[27] ^ input_a[11];
  assign popcount36_w9zx_core_240 = input_a[27] | input_a[27];
  assign popcount36_w9zx_core_242 = ~(input_a[20] & input_a[12]);
  assign popcount36_w9zx_core_243 = ~(input_a[1] & input_a[18]);
  assign popcount36_w9zx_core_244 = ~(input_a[8] & input_a[31]);
  assign popcount36_w9zx_core_245 = input_a[17] ^ input_a[30];
  assign popcount36_w9zx_core_246 = input_a[7] | input_a[9];
  assign popcount36_w9zx_core_247 = ~input_a[7];
  assign popcount36_w9zx_core_248 = input_a[15] & input_a[2];
  assign popcount36_w9zx_core_249 = input_a[22] ^ input_a[10];
  assign popcount36_w9zx_core_251 = input_a[14] | input_a[23];
  assign popcount36_w9zx_core_252 = ~(input_a[6] ^ input_a[26]);
  assign popcount36_w9zx_core_254 = ~input_a[11];
  assign popcount36_w9zx_core_255 = ~input_a[27];
  assign popcount36_w9zx_core_258 = input_a[14] ^ input_a[29];
  assign popcount36_w9zx_core_259 = input_a[32] | input_a[16];
  assign popcount36_w9zx_core_260 = input_a[19] | input_a[24];
  assign popcount36_w9zx_core_261 = input_a[28] ^ input_a[30];
  assign popcount36_w9zx_core_262 = input_a[17] & input_a[24];
  assign popcount36_w9zx_core_263 = input_a[27] | input_a[5];
  assign popcount36_w9zx_core_264 = input_a[5] ^ input_a[10];
  assign popcount36_w9zx_core_266 = ~input_a[34];
  assign popcount36_w9zx_core_267 = input_a[18] ^ input_a[9];
  assign popcount36_w9zx_core_268 = input_a[26] & input_a[32];
  assign popcount36_w9zx_core_269 = ~input_a[16];
  assign popcount36_w9zx_core_271 = input_a[15] | input_a[16];
  assign popcount36_w9zx_core_272 = ~(input_a[5] ^ input_a[7]);
  assign popcount36_w9zx_core_274 = ~(input_a[19] | input_a[12]);
  assign popcount36_w9zx_core_275 = ~(input_a[11] | input_a[23]);

  assign popcount36_w9zx_out[0] = input_a[19];
  assign popcount36_w9zx_out[1] = input_a[11];
  assign popcount36_w9zx_out[2] = input_a[20];
  assign popcount36_w9zx_out[3] = input_a[35];
  assign popcount36_w9zx_out[4] = 1'b1;
  assign popcount36_w9zx_out[5] = 1'b0;
endmodule