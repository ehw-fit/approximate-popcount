// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.67499
// WCE=13.0
// EP=0.886026%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_htwf(input [20:0] input_a, output [4:0] popcount21_htwf_out);
  wire popcount21_htwf_core_023;
  wire popcount21_htwf_core_025;
  wire popcount21_htwf_core_027;
  wire popcount21_htwf_core_029_not;
  wire popcount21_htwf_core_031;
  wire popcount21_htwf_core_033_not;
  wire popcount21_htwf_core_035;
  wire popcount21_htwf_core_036;
  wire popcount21_htwf_core_037;
  wire popcount21_htwf_core_039;
  wire popcount21_htwf_core_040;
  wire popcount21_htwf_core_041;
  wire popcount21_htwf_core_042;
  wire popcount21_htwf_core_044;
  wire popcount21_htwf_core_045;
  wire popcount21_htwf_core_048;
  wire popcount21_htwf_core_049;
  wire popcount21_htwf_core_051;
  wire popcount21_htwf_core_053;
  wire popcount21_htwf_core_054;
  wire popcount21_htwf_core_055;
  wire popcount21_htwf_core_056;
  wire popcount21_htwf_core_058;
  wire popcount21_htwf_core_059;
  wire popcount21_htwf_core_060;
  wire popcount21_htwf_core_061;
  wire popcount21_htwf_core_063;
  wire popcount21_htwf_core_064;
  wire popcount21_htwf_core_065;
  wire popcount21_htwf_core_066;
  wire popcount21_htwf_core_067;
  wire popcount21_htwf_core_069;
  wire popcount21_htwf_core_072;
  wire popcount21_htwf_core_073;
  wire popcount21_htwf_core_074;
  wire popcount21_htwf_core_076;
  wire popcount21_htwf_core_078;
  wire popcount21_htwf_core_081;
  wire popcount21_htwf_core_082;
  wire popcount21_htwf_core_088;
  wire popcount21_htwf_core_090;
  wire popcount21_htwf_core_092_not;
  wire popcount21_htwf_core_094;
  wire popcount21_htwf_core_096;
  wire popcount21_htwf_core_097;
  wire popcount21_htwf_core_098;
  wire popcount21_htwf_core_099;
  wire popcount21_htwf_core_100;
  wire popcount21_htwf_core_101;
  wire popcount21_htwf_core_102;
  wire popcount21_htwf_core_103;
  wire popcount21_htwf_core_104;
  wire popcount21_htwf_core_106;
  wire popcount21_htwf_core_107;
  wire popcount21_htwf_core_108;
  wire popcount21_htwf_core_110;
  wire popcount21_htwf_core_111;
  wire popcount21_htwf_core_112;
  wire popcount21_htwf_core_114;
  wire popcount21_htwf_core_115;
  wire popcount21_htwf_core_118;
  wire popcount21_htwf_core_120;
  wire popcount21_htwf_core_121;
  wire popcount21_htwf_core_126;
  wire popcount21_htwf_core_127;
  wire popcount21_htwf_core_128;
  wire popcount21_htwf_core_130;
  wire popcount21_htwf_core_133;
  wire popcount21_htwf_core_134;
  wire popcount21_htwf_core_135;
  wire popcount21_htwf_core_136;
  wire popcount21_htwf_core_137;
  wire popcount21_htwf_core_140;
  wire popcount21_htwf_core_141;
  wire popcount21_htwf_core_143;
  wire popcount21_htwf_core_145;
  wire popcount21_htwf_core_148;
  wire popcount21_htwf_core_149;
  wire popcount21_htwf_core_150_not;
  wire popcount21_htwf_core_152;

  assign popcount21_htwf_core_023 = input_a[6] ^ input_a[1];
  assign popcount21_htwf_core_025 = ~(input_a[8] & input_a[2]);
  assign popcount21_htwf_core_027 = ~(input_a[20] | input_a[18]);
  assign popcount21_htwf_core_029_not = ~input_a[0];
  assign popcount21_htwf_core_031 = ~input_a[12];
  assign popcount21_htwf_core_033_not = ~input_a[17];
  assign popcount21_htwf_core_035 = ~(input_a[16] & input_a[20]);
  assign popcount21_htwf_core_036 = ~(input_a[4] & input_a[13]);
  assign popcount21_htwf_core_037 = input_a[19] | input_a[20];
  assign popcount21_htwf_core_039 = ~input_a[6];
  assign popcount21_htwf_core_040 = input_a[3] ^ input_a[13];
  assign popcount21_htwf_core_041 = ~(input_a[4] ^ input_a[6]);
  assign popcount21_htwf_core_042 = input_a[0] & input_a[4];
  assign popcount21_htwf_core_044 = ~(input_a[12] | input_a[2]);
  assign popcount21_htwf_core_045 = input_a[11] | input_a[2];
  assign popcount21_htwf_core_048 = input_a[6] & input_a[10];
  assign popcount21_htwf_core_049 = input_a[6] ^ input_a[7];
  assign popcount21_htwf_core_051 = input_a[0] ^ input_a[17];
  assign popcount21_htwf_core_053 = input_a[9] | input_a[14];
  assign popcount21_htwf_core_054 = ~(input_a[0] & input_a[4]);
  assign popcount21_htwf_core_055 = input_a[9] | input_a[15];
  assign popcount21_htwf_core_056 = ~(input_a[19] | input_a[14]);
  assign popcount21_htwf_core_058 = input_a[16] ^ input_a[7];
  assign popcount21_htwf_core_059 = ~(input_a[19] ^ input_a[7]);
  assign popcount21_htwf_core_060 = input_a[12] & input_a[0];
  assign popcount21_htwf_core_061 = ~input_a[13];
  assign popcount21_htwf_core_063 = ~(input_a[4] | input_a[20]);
  assign popcount21_htwf_core_064 = ~(input_a[16] & input_a[9]);
  assign popcount21_htwf_core_065 = ~(input_a[14] ^ input_a[7]);
  assign popcount21_htwf_core_066 = ~(input_a[8] ^ input_a[3]);
  assign popcount21_htwf_core_067 = ~input_a[3];
  assign popcount21_htwf_core_069 = ~(input_a[5] | input_a[19]);
  assign popcount21_htwf_core_072 = ~(input_a[6] ^ input_a[2]);
  assign popcount21_htwf_core_073 = input_a[19] & input_a[2];
  assign popcount21_htwf_core_074 = ~(input_a[6] & input_a[19]);
  assign popcount21_htwf_core_076 = input_a[7] | input_a[13];
  assign popcount21_htwf_core_078 = ~(input_a[9] | input_a[20]);
  assign popcount21_htwf_core_081 = ~(input_a[10] ^ input_a[20]);
  assign popcount21_htwf_core_082 = input_a[13] & input_a[1];
  assign popcount21_htwf_core_088 = input_a[9] & input_a[13];
  assign popcount21_htwf_core_090 = ~(input_a[13] | input_a[3]);
  assign popcount21_htwf_core_092_not = ~input_a[17];
  assign popcount21_htwf_core_094 = input_a[4] & input_a[9];
  assign popcount21_htwf_core_096 = input_a[13] | input_a[16];
  assign popcount21_htwf_core_097 = ~(input_a[9] ^ input_a[4]);
  assign popcount21_htwf_core_098 = ~(input_a[5] | input_a[12]);
  assign popcount21_htwf_core_099 = input_a[9] | input_a[8];
  assign popcount21_htwf_core_100 = ~(input_a[8] | input_a[16]);
  assign popcount21_htwf_core_101 = ~input_a[3];
  assign popcount21_htwf_core_102 = ~(input_a[20] & input_a[17]);
  assign popcount21_htwf_core_103 = ~(input_a[7] & input_a[14]);
  assign popcount21_htwf_core_104 = input_a[15] & input_a[19];
  assign popcount21_htwf_core_106 = input_a[0] & input_a[2];
  assign popcount21_htwf_core_107 = ~(input_a[1] ^ input_a[14]);
  assign popcount21_htwf_core_108 = input_a[11] ^ input_a[17];
  assign popcount21_htwf_core_110 = input_a[8] & input_a[0];
  assign popcount21_htwf_core_111 = input_a[16] | input_a[2];
  assign popcount21_htwf_core_112 = ~(input_a[11] ^ input_a[6]);
  assign popcount21_htwf_core_114 = input_a[18] & input_a[16];
  assign popcount21_htwf_core_115 = ~(input_a[17] ^ input_a[11]);
  assign popcount21_htwf_core_118 = input_a[5] & input_a[18];
  assign popcount21_htwf_core_120 = input_a[13] ^ input_a[13];
  assign popcount21_htwf_core_121 = input_a[6] | input_a[5];
  assign popcount21_htwf_core_126 = input_a[11] | input_a[18];
  assign popcount21_htwf_core_127 = ~(input_a[16] | input_a[1]);
  assign popcount21_htwf_core_128 = ~(input_a[0] | input_a[1]);
  assign popcount21_htwf_core_130 = ~input_a[1];
  assign popcount21_htwf_core_133 = input_a[9] | input_a[3];
  assign popcount21_htwf_core_134 = ~(input_a[18] | input_a[3]);
  assign popcount21_htwf_core_135 = input_a[8] & input_a[16];
  assign popcount21_htwf_core_136 = input_a[2] ^ input_a[10];
  assign popcount21_htwf_core_137 = input_a[4] & input_a[0];
  assign popcount21_htwf_core_140 = ~(input_a[4] | input_a[19]);
  assign popcount21_htwf_core_141 = input_a[12] | input_a[3];
  assign popcount21_htwf_core_143 = ~(input_a[13] ^ input_a[0]);
  assign popcount21_htwf_core_145 = input_a[17] & input_a[2];
  assign popcount21_htwf_core_148 = ~(input_a[2] ^ input_a[5]);
  assign popcount21_htwf_core_149 = ~(input_a[6] & input_a[4]);
  assign popcount21_htwf_core_150_not = ~input_a[7];
  assign popcount21_htwf_core_152 = input_a[17] | input_a[12];

  assign popcount21_htwf_out[0] = input_a[2];
  assign popcount21_htwf_out[1] = 1'b1;
  assign popcount21_htwf_out[2] = input_a[5];
  assign popcount21_htwf_out[3] = 1'b1;
  assign popcount21_htwf_out[4] = 1'b0;
endmodule