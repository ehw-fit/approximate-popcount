// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.86159
// WCE=19.0
// EP=0.93047%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_3baw(input [29:0] input_a, output [4:0] popcount30_3baw_out);
  wire popcount30_3baw_core_033;
  wire popcount30_3baw_core_038;
  wire popcount30_3baw_core_039;
  wire popcount30_3baw_core_040;
  wire popcount30_3baw_core_041;
  wire popcount30_3baw_core_043;
  wire popcount30_3baw_core_044;
  wire popcount30_3baw_core_049;
  wire popcount30_3baw_core_050;
  wire popcount30_3baw_core_052;
  wire popcount30_3baw_core_053;
  wire popcount30_3baw_core_054;
  wire popcount30_3baw_core_058;
  wire popcount30_3baw_core_059;
  wire popcount30_3baw_core_060;
  wire popcount30_3baw_core_061;
  wire popcount30_3baw_core_062;
  wire popcount30_3baw_core_066_not;
  wire popcount30_3baw_core_067;
  wire popcount30_3baw_core_068;
  wire popcount30_3baw_core_069;
  wire popcount30_3baw_core_074;
  wire popcount30_3baw_core_075;
  wire popcount30_3baw_core_076;
  wire popcount30_3baw_core_077;
  wire popcount30_3baw_core_078;
  wire popcount30_3baw_core_081_not;
  wire popcount30_3baw_core_082;
  wire popcount30_3baw_core_083;
  wire popcount30_3baw_core_084;
  wire popcount30_3baw_core_087;
  wire popcount30_3baw_core_089;
  wire popcount30_3baw_core_090;
  wire popcount30_3baw_core_093;
  wire popcount30_3baw_core_094;
  wire popcount30_3baw_core_095;
  wire popcount30_3baw_core_096;
  wire popcount30_3baw_core_102;
  wire popcount30_3baw_core_103;
  wire popcount30_3baw_core_105;
  wire popcount30_3baw_core_106;
  wire popcount30_3baw_core_107;
  wire popcount30_3baw_core_108;
  wire popcount30_3baw_core_109;
  wire popcount30_3baw_core_112;
  wire popcount30_3baw_core_113;
  wire popcount30_3baw_core_116;
  wire popcount30_3baw_core_117;
  wire popcount30_3baw_core_119;
  wire popcount30_3baw_core_120;
  wire popcount30_3baw_core_121;
  wire popcount30_3baw_core_122;
  wire popcount30_3baw_core_123;
  wire popcount30_3baw_core_124;
  wire popcount30_3baw_core_126_not;
  wire popcount30_3baw_core_127;
  wire popcount30_3baw_core_128;
  wire popcount30_3baw_core_132;
  wire popcount30_3baw_core_135;
  wire popcount30_3baw_core_137;
  wire popcount30_3baw_core_138;
  wire popcount30_3baw_core_139;
  wire popcount30_3baw_core_140;
  wire popcount30_3baw_core_142;
  wire popcount30_3baw_core_143;
  wire popcount30_3baw_core_144;
  wire popcount30_3baw_core_153;
  wire popcount30_3baw_core_155;
  wire popcount30_3baw_core_156;
  wire popcount30_3baw_core_159_not;
  wire popcount30_3baw_core_160;
  wire popcount30_3baw_core_161;
  wire popcount30_3baw_core_162;
  wire popcount30_3baw_core_163;
  wire popcount30_3baw_core_164;
  wire popcount30_3baw_core_166;
  wire popcount30_3baw_core_168;
  wire popcount30_3baw_core_169;
  wire popcount30_3baw_core_170_not;
  wire popcount30_3baw_core_172;
  wire popcount30_3baw_core_173;
  wire popcount30_3baw_core_174;
  wire popcount30_3baw_core_176;
  wire popcount30_3baw_core_178;
  wire popcount30_3baw_core_180;
  wire popcount30_3baw_core_181;
  wire popcount30_3baw_core_182;
  wire popcount30_3baw_core_183;
  wire popcount30_3baw_core_185;
  wire popcount30_3baw_core_186;
  wire popcount30_3baw_core_187_not;
  wire popcount30_3baw_core_189;
  wire popcount30_3baw_core_190;
  wire popcount30_3baw_core_191_not;
  wire popcount30_3baw_core_193;
  wire popcount30_3baw_core_194_not;
  wire popcount30_3baw_core_195;
  wire popcount30_3baw_core_196;
  wire popcount30_3baw_core_197;
  wire popcount30_3baw_core_198;
  wire popcount30_3baw_core_200;
  wire popcount30_3baw_core_201;
  wire popcount30_3baw_core_203;
  wire popcount30_3baw_core_204;
  wire popcount30_3baw_core_205;
  wire popcount30_3baw_core_206;
  wire popcount30_3baw_core_207;
  wire popcount30_3baw_core_208;
  wire popcount30_3baw_core_209;
  wire popcount30_3baw_core_210_not;
  wire popcount30_3baw_core_211;
  wire popcount30_3baw_core_212;

  assign popcount30_3baw_core_033 = ~(input_a[15] & input_a[7]);
  assign popcount30_3baw_core_038 = input_a[28] | input_a[21];
  assign popcount30_3baw_core_039 = ~input_a[11];
  assign popcount30_3baw_core_040 = ~input_a[21];
  assign popcount30_3baw_core_041 = input_a[10] | input_a[13];
  assign popcount30_3baw_core_043 = input_a[1] & input_a[20];
  assign popcount30_3baw_core_044 = ~(input_a[11] & input_a[10]);
  assign popcount30_3baw_core_049 = ~(input_a[13] | input_a[9]);
  assign popcount30_3baw_core_050 = ~(input_a[6] ^ input_a[28]);
  assign popcount30_3baw_core_052 = input_a[9] | input_a[17];
  assign popcount30_3baw_core_053 = input_a[5] | input_a[6];
  assign popcount30_3baw_core_054 = input_a[14] & input_a[14];
  assign popcount30_3baw_core_058 = input_a[10] | input_a[19];
  assign popcount30_3baw_core_059 = input_a[22] ^ input_a[8];
  assign popcount30_3baw_core_060 = ~input_a[18];
  assign popcount30_3baw_core_061 = input_a[15] | input_a[26];
  assign popcount30_3baw_core_062 = ~input_a[9];
  assign popcount30_3baw_core_066_not = ~input_a[3];
  assign popcount30_3baw_core_067 = ~(input_a[2] | input_a[13]);
  assign popcount30_3baw_core_068 = input_a[4] | input_a[24];
  assign popcount30_3baw_core_069 = input_a[14] | input_a[25];
  assign popcount30_3baw_core_074 = input_a[10] | input_a[19];
  assign popcount30_3baw_core_075 = ~(input_a[5] & input_a[19]);
  assign popcount30_3baw_core_076 = ~(input_a[18] | input_a[21]);
  assign popcount30_3baw_core_077 = input_a[4] ^ input_a[29];
  assign popcount30_3baw_core_078 = input_a[3] & input_a[24];
  assign popcount30_3baw_core_081_not = ~input_a[23];
  assign popcount30_3baw_core_082 = ~(input_a[21] | input_a[28]);
  assign popcount30_3baw_core_083 = input_a[0] ^ input_a[25];
  assign popcount30_3baw_core_084 = input_a[29] | input_a[24];
  assign popcount30_3baw_core_087 = ~input_a[9];
  assign popcount30_3baw_core_089 = input_a[27] | input_a[17];
  assign popcount30_3baw_core_090 = input_a[23] | input_a[6];
  assign popcount30_3baw_core_093 = input_a[20] | input_a[0];
  assign popcount30_3baw_core_094 = input_a[8] | input_a[13];
  assign popcount30_3baw_core_095 = ~(input_a[29] ^ input_a[29]);
  assign popcount30_3baw_core_096 = ~(input_a[13] | input_a[7]);
  assign popcount30_3baw_core_102 = input_a[21] & input_a[0];
  assign popcount30_3baw_core_103 = ~(input_a[10] & input_a[26]);
  assign popcount30_3baw_core_105 = ~(input_a[22] & input_a[11]);
  assign popcount30_3baw_core_106 = ~input_a[3];
  assign popcount30_3baw_core_107 = input_a[13] & input_a[4];
  assign popcount30_3baw_core_108 = input_a[21] | input_a[26];
  assign popcount30_3baw_core_109 = ~(input_a[2] & input_a[22]);
  assign popcount30_3baw_core_112 = input_a[7] | input_a[25];
  assign popcount30_3baw_core_113 = ~(input_a[13] & input_a[5]);
  assign popcount30_3baw_core_116 = ~input_a[21];
  assign popcount30_3baw_core_117 = ~input_a[18];
  assign popcount30_3baw_core_119 = ~(input_a[23] & input_a[6]);
  assign popcount30_3baw_core_120 = ~(input_a[24] | input_a[12]);
  assign popcount30_3baw_core_121 = ~(input_a[28] ^ input_a[5]);
  assign popcount30_3baw_core_122 = input_a[26] & input_a[8];
  assign popcount30_3baw_core_123 = ~(input_a[29] & input_a[0]);
  assign popcount30_3baw_core_124 = ~input_a[23];
  assign popcount30_3baw_core_126_not = ~input_a[14];
  assign popcount30_3baw_core_127 = ~(input_a[3] & input_a[19]);
  assign popcount30_3baw_core_128 = ~(input_a[7] ^ input_a[9]);
  assign popcount30_3baw_core_132 = ~input_a[17];
  assign popcount30_3baw_core_135 = ~input_a[1];
  assign popcount30_3baw_core_137 = ~input_a[19];
  assign popcount30_3baw_core_138 = input_a[10] | input_a[13];
  assign popcount30_3baw_core_139 = ~input_a[20];
  assign popcount30_3baw_core_140 = ~input_a[27];
  assign popcount30_3baw_core_142 = ~input_a[29];
  assign popcount30_3baw_core_143 = input_a[11] ^ input_a[26];
  assign popcount30_3baw_core_144 = ~(input_a[18] & input_a[22]);
  assign popcount30_3baw_core_153 = input_a[19] ^ input_a[17];
  assign popcount30_3baw_core_155 = ~(input_a[7] ^ input_a[3]);
  assign popcount30_3baw_core_156 = input_a[5] & input_a[26];
  assign popcount30_3baw_core_159_not = ~input_a[17];
  assign popcount30_3baw_core_160 = input_a[21] & input_a[8];
  assign popcount30_3baw_core_161 = ~(input_a[5] | input_a[11]);
  assign popcount30_3baw_core_162 = input_a[25] ^ input_a[27];
  assign popcount30_3baw_core_163 = input_a[4] & input_a[13];
  assign popcount30_3baw_core_164 = ~(input_a[5] ^ input_a[3]);
  assign popcount30_3baw_core_166 = input_a[26] & input_a[0];
  assign popcount30_3baw_core_168 = ~(input_a[6] & input_a[6]);
  assign popcount30_3baw_core_169 = ~input_a[29];
  assign popcount30_3baw_core_170_not = ~input_a[6];
  assign popcount30_3baw_core_172 = ~input_a[7];
  assign popcount30_3baw_core_173 = input_a[4] | input_a[27];
  assign popcount30_3baw_core_174 = input_a[19] ^ input_a[11];
  assign popcount30_3baw_core_176 = ~(input_a[27] & input_a[23]);
  assign popcount30_3baw_core_178 = input_a[4] | input_a[14];
  assign popcount30_3baw_core_180 = ~(input_a[28] ^ input_a[19]);
  assign popcount30_3baw_core_181 = ~(input_a[14] | input_a[11]);
  assign popcount30_3baw_core_182 = input_a[26] | input_a[6];
  assign popcount30_3baw_core_183 = ~(input_a[21] & input_a[24]);
  assign popcount30_3baw_core_185 = input_a[18] | input_a[25];
  assign popcount30_3baw_core_186 = input_a[13] ^ input_a[20];
  assign popcount30_3baw_core_187_not = ~input_a[8];
  assign popcount30_3baw_core_189 = input_a[28] ^ input_a[24];
  assign popcount30_3baw_core_190 = ~input_a[22];
  assign popcount30_3baw_core_191_not = ~input_a[12];
  assign popcount30_3baw_core_193 = ~(input_a[21] ^ input_a[9]);
  assign popcount30_3baw_core_194_not = ~input_a[11];
  assign popcount30_3baw_core_195 = ~(input_a[24] & input_a[23]);
  assign popcount30_3baw_core_196 = input_a[12] | input_a[23];
  assign popcount30_3baw_core_197 = ~(input_a[7] ^ input_a[4]);
  assign popcount30_3baw_core_198 = ~input_a[25];
  assign popcount30_3baw_core_200 = ~(input_a[14] & input_a[7]);
  assign popcount30_3baw_core_201 = ~(input_a[21] & input_a[16]);
  assign popcount30_3baw_core_203 = ~(input_a[14] | input_a[26]);
  assign popcount30_3baw_core_204 = ~(input_a[20] & input_a[14]);
  assign popcount30_3baw_core_205 = ~input_a[0];
  assign popcount30_3baw_core_206 = input_a[19] | input_a[11];
  assign popcount30_3baw_core_207 = input_a[0] & input_a[22];
  assign popcount30_3baw_core_208 = input_a[2] | input_a[5];
  assign popcount30_3baw_core_209 = ~(input_a[25] ^ input_a[10]);
  assign popcount30_3baw_core_210_not = ~input_a[7];
  assign popcount30_3baw_core_211 = ~(input_a[24] & input_a[14]);
  assign popcount30_3baw_core_212 = ~(input_a[27] & input_a[3]);

  assign popcount30_3baw_out[0] = input_a[16];
  assign popcount30_3baw_out[1] = input_a[14];
  assign popcount30_3baw_out[2] = input_a[18];
  assign popcount30_3baw_out[3] = 1'b1;
  assign popcount30_3baw_out[4] = 1'b0;
endmodule