// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.46801
// WCE=19.0
// EP=0.918143%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_aewx(input [24:0] input_a, output [4:0] popcount25_aewx_out);
  wire popcount25_aewx_core_027;
  wire popcount25_aewx_core_028;
  wire popcount25_aewx_core_029;
  wire popcount25_aewx_core_032;
  wire popcount25_aewx_core_033;
  wire popcount25_aewx_core_036;
  wire popcount25_aewx_core_037;
  wire popcount25_aewx_core_039;
  wire popcount25_aewx_core_040;
  wire popcount25_aewx_core_045;
  wire popcount25_aewx_core_046;
  wire popcount25_aewx_core_047;
  wire popcount25_aewx_core_048;
  wire popcount25_aewx_core_050;
  wire popcount25_aewx_core_051;
  wire popcount25_aewx_core_053;
  wire popcount25_aewx_core_056;
  wire popcount25_aewx_core_057;
  wire popcount25_aewx_core_058;
  wire popcount25_aewx_core_061;
  wire popcount25_aewx_core_062;
  wire popcount25_aewx_core_063;
  wire popcount25_aewx_core_065;
  wire popcount25_aewx_core_066_not;
  wire popcount25_aewx_core_067;
  wire popcount25_aewx_core_068;
  wire popcount25_aewx_core_069;
  wire popcount25_aewx_core_070;
  wire popcount25_aewx_core_075;
  wire popcount25_aewx_core_077_not;
  wire popcount25_aewx_core_079;
  wire popcount25_aewx_core_080;
  wire popcount25_aewx_core_081;
  wire popcount25_aewx_core_082;
  wire popcount25_aewx_core_086;
  wire popcount25_aewx_core_087;
  wire popcount25_aewx_core_089;
  wire popcount25_aewx_core_090;
  wire popcount25_aewx_core_092;
  wire popcount25_aewx_core_093;
  wire popcount25_aewx_core_095;
  wire popcount25_aewx_core_096_not;
  wire popcount25_aewx_core_097;
  wire popcount25_aewx_core_099;
  wire popcount25_aewx_core_100;
  wire popcount25_aewx_core_101;
  wire popcount25_aewx_core_102;
  wire popcount25_aewx_core_105;
  wire popcount25_aewx_core_108;
  wire popcount25_aewx_core_111;
  wire popcount25_aewx_core_112_not;
  wire popcount25_aewx_core_113;
  wire popcount25_aewx_core_115;
  wire popcount25_aewx_core_116;
  wire popcount25_aewx_core_117;
  wire popcount25_aewx_core_118;
  wire popcount25_aewx_core_119;
  wire popcount25_aewx_core_122;
  wire popcount25_aewx_core_123;
  wire popcount25_aewx_core_125;
  wire popcount25_aewx_core_126;
  wire popcount25_aewx_core_127;
  wire popcount25_aewx_core_128;
  wire popcount25_aewx_core_129;
  wire popcount25_aewx_core_130;
  wire popcount25_aewx_core_133;
  wire popcount25_aewx_core_134;
  wire popcount25_aewx_core_136;
  wire popcount25_aewx_core_137;
  wire popcount25_aewx_core_147;
  wire popcount25_aewx_core_148;
  wire popcount25_aewx_core_149;
  wire popcount25_aewx_core_151;
  wire popcount25_aewx_core_157;
  wire popcount25_aewx_core_158;
  wire popcount25_aewx_core_159;
  wire popcount25_aewx_core_160;
  wire popcount25_aewx_core_166;
  wire popcount25_aewx_core_167;
  wire popcount25_aewx_core_170;
  wire popcount25_aewx_core_171;
  wire popcount25_aewx_core_175;
  wire popcount25_aewx_core_176;
  wire popcount25_aewx_core_177;
  wire popcount25_aewx_core_181;

  assign popcount25_aewx_core_027 = input_a[21] ^ input_a[5];
  assign popcount25_aewx_core_028 = ~(input_a[14] & input_a[20]);
  assign popcount25_aewx_core_029 = ~(input_a[13] ^ input_a[7]);
  assign popcount25_aewx_core_032 = ~(input_a[24] & input_a[0]);
  assign popcount25_aewx_core_033 = ~(input_a[5] & input_a[15]);
  assign popcount25_aewx_core_036 = ~(input_a[6] ^ input_a[14]);
  assign popcount25_aewx_core_037 = ~(input_a[4] | input_a[7]);
  assign popcount25_aewx_core_039 = input_a[24] & input_a[21];
  assign popcount25_aewx_core_040 = ~input_a[16];
  assign popcount25_aewx_core_045 = input_a[19] & input_a[2];
  assign popcount25_aewx_core_046 = ~(input_a[21] ^ input_a[0]);
  assign popcount25_aewx_core_047 = input_a[2] ^ input_a[7];
  assign popcount25_aewx_core_048 = ~input_a[5];
  assign popcount25_aewx_core_050 = ~(input_a[24] ^ input_a[14]);
  assign popcount25_aewx_core_051 = input_a[13] & input_a[22];
  assign popcount25_aewx_core_053 = input_a[19] ^ input_a[16];
  assign popcount25_aewx_core_056 = input_a[18] ^ input_a[6];
  assign popcount25_aewx_core_057 = ~(input_a[15] | input_a[22]);
  assign popcount25_aewx_core_058 = ~input_a[15];
  assign popcount25_aewx_core_061 = input_a[2] & input_a[20];
  assign popcount25_aewx_core_062 = ~(input_a[2] | input_a[5]);
  assign popcount25_aewx_core_063 = ~input_a[11];
  assign popcount25_aewx_core_065 = input_a[13] | input_a[24];
  assign popcount25_aewx_core_066_not = ~input_a[8];
  assign popcount25_aewx_core_067 = ~(input_a[22] | input_a[16]);
  assign popcount25_aewx_core_068 = ~(input_a[7] | input_a[19]);
  assign popcount25_aewx_core_069 = ~input_a[16];
  assign popcount25_aewx_core_070 = input_a[24] ^ input_a[18];
  assign popcount25_aewx_core_075 = ~(input_a[21] ^ input_a[24]);
  assign popcount25_aewx_core_077_not = ~input_a[12];
  assign popcount25_aewx_core_079 = ~(input_a[23] | input_a[8]);
  assign popcount25_aewx_core_080 = ~(input_a[2] | input_a[8]);
  assign popcount25_aewx_core_081 = input_a[10] | input_a[11];
  assign popcount25_aewx_core_082 = input_a[15] ^ input_a[20];
  assign popcount25_aewx_core_086 = ~(input_a[9] ^ input_a[10]);
  assign popcount25_aewx_core_087 = ~(input_a[0] ^ input_a[10]);
  assign popcount25_aewx_core_089 = ~(input_a[4] ^ input_a[2]);
  assign popcount25_aewx_core_090 = ~(input_a[20] & input_a[13]);
  assign popcount25_aewx_core_092 = ~(input_a[8] ^ input_a[0]);
  assign popcount25_aewx_core_093 = input_a[21] | input_a[3];
  assign popcount25_aewx_core_095 = ~(input_a[13] | input_a[4]);
  assign popcount25_aewx_core_096_not = ~input_a[10];
  assign popcount25_aewx_core_097 = ~(input_a[6] & input_a[21]);
  assign popcount25_aewx_core_099 = ~(input_a[10] & input_a[5]);
  assign popcount25_aewx_core_100 = ~(input_a[1] ^ input_a[12]);
  assign popcount25_aewx_core_101 = input_a[14] ^ input_a[8];
  assign popcount25_aewx_core_102 = input_a[13] ^ input_a[12];
  assign popcount25_aewx_core_105 = ~(input_a[2] | input_a[5]);
  assign popcount25_aewx_core_108 = ~(input_a[21] & input_a[3]);
  assign popcount25_aewx_core_111 = input_a[17] ^ input_a[22];
  assign popcount25_aewx_core_112_not = ~input_a[3];
  assign popcount25_aewx_core_113 = ~(input_a[8] & input_a[0]);
  assign popcount25_aewx_core_115 = ~(input_a[19] | input_a[10]);
  assign popcount25_aewx_core_116 = input_a[14] & input_a[24];
  assign popcount25_aewx_core_117 = input_a[23] | input_a[12];
  assign popcount25_aewx_core_118 = ~(input_a[3] | input_a[12]);
  assign popcount25_aewx_core_119 = input_a[14] & input_a[5];
  assign popcount25_aewx_core_122 = ~(input_a[24] & input_a[11]);
  assign popcount25_aewx_core_123 = input_a[6] & input_a[9];
  assign popcount25_aewx_core_125 = input_a[7] ^ input_a[9];
  assign popcount25_aewx_core_126 = ~(input_a[21] & input_a[17]);
  assign popcount25_aewx_core_127 = input_a[7] & input_a[9];
  assign popcount25_aewx_core_128 = ~(input_a[7] ^ input_a[17]);
  assign popcount25_aewx_core_129 = ~(input_a[12] ^ input_a[16]);
  assign popcount25_aewx_core_130 = ~(input_a[7] ^ input_a[10]);
  assign popcount25_aewx_core_133 = input_a[0] | input_a[12];
  assign popcount25_aewx_core_134 = input_a[2] & input_a[13];
  assign popcount25_aewx_core_136 = ~input_a[22];
  assign popcount25_aewx_core_137 = input_a[11] & input_a[16];
  assign popcount25_aewx_core_147 = input_a[11] & input_a[19];
  assign popcount25_aewx_core_148 = ~input_a[17];
  assign popcount25_aewx_core_149 = ~input_a[13];
  assign popcount25_aewx_core_151 = ~input_a[17];
  assign popcount25_aewx_core_157 = input_a[19] & input_a[20];
  assign popcount25_aewx_core_158 = ~(input_a[12] | input_a[9]);
  assign popcount25_aewx_core_159 = ~input_a[0];
  assign popcount25_aewx_core_160 = input_a[10] ^ input_a[13];
  assign popcount25_aewx_core_166 = ~(input_a[4] & input_a[22]);
  assign popcount25_aewx_core_167 = input_a[5] ^ input_a[17];
  assign popcount25_aewx_core_170 = input_a[17] | input_a[24];
  assign popcount25_aewx_core_171 = input_a[8] & input_a[16];
  assign popcount25_aewx_core_175 = input_a[24] ^ input_a[8];
  assign popcount25_aewx_core_176 = input_a[16] | input_a[16];
  assign popcount25_aewx_core_177 = input_a[3] & input_a[16];
  assign popcount25_aewx_core_181 = input_a[9] | input_a[8];

  assign popcount25_aewx_out[0] = 1'b0;
  assign popcount25_aewx_out[1] = input_a[0];
  assign popcount25_aewx_out[2] = 1'b1;
  assign popcount25_aewx_out[3] = input_a[13];
  assign popcount25_aewx_out[4] = 1'b0;
endmodule