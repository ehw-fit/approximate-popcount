// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.84736
// WCE=27.0
// EP=0.921989%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount45_dokv(input [44:0] input_a, output [5:0] popcount45_dokv_out);
  wire popcount45_dokv_core_049;
  wire popcount45_dokv_core_051;
  wire popcount45_dokv_core_052;
  wire popcount45_dokv_core_054;
  wire popcount45_dokv_core_055;
  wire popcount45_dokv_core_056;
  wire popcount45_dokv_core_057;
  wire popcount45_dokv_core_059;
  wire popcount45_dokv_core_061;
  wire popcount45_dokv_core_062;
  wire popcount45_dokv_core_063;
  wire popcount45_dokv_core_064;
  wire popcount45_dokv_core_065;
  wire popcount45_dokv_core_066;
  wire popcount45_dokv_core_068;
  wire popcount45_dokv_core_071;
  wire popcount45_dokv_core_072;
  wire popcount45_dokv_core_073;
  wire popcount45_dokv_core_075;
  wire popcount45_dokv_core_076;
  wire popcount45_dokv_core_077;
  wire popcount45_dokv_core_078;
  wire popcount45_dokv_core_079;
  wire popcount45_dokv_core_081;
  wire popcount45_dokv_core_083_not;
  wire popcount45_dokv_core_085;
  wire popcount45_dokv_core_086;
  wire popcount45_dokv_core_087;
  wire popcount45_dokv_core_089;
  wire popcount45_dokv_core_090;
  wire popcount45_dokv_core_092;
  wire popcount45_dokv_core_093;
  wire popcount45_dokv_core_094;
  wire popcount45_dokv_core_096;
  wire popcount45_dokv_core_098;
  wire popcount45_dokv_core_101;
  wire popcount45_dokv_core_102;
  wire popcount45_dokv_core_104;
  wire popcount45_dokv_core_105;
  wire popcount45_dokv_core_106;
  wire popcount45_dokv_core_107;
  wire popcount45_dokv_core_108;
  wire popcount45_dokv_core_113;
  wire popcount45_dokv_core_114;
  wire popcount45_dokv_core_116;
  wire popcount45_dokv_core_117;
  wire popcount45_dokv_core_118;
  wire popcount45_dokv_core_121;
  wire popcount45_dokv_core_126;
  wire popcount45_dokv_core_127;
  wire popcount45_dokv_core_128;
  wire popcount45_dokv_core_129;
  wire popcount45_dokv_core_130;
  wire popcount45_dokv_core_131_not;
  wire popcount45_dokv_core_133;
  wire popcount45_dokv_core_134;
  wire popcount45_dokv_core_135;
  wire popcount45_dokv_core_137;
  wire popcount45_dokv_core_139;
  wire popcount45_dokv_core_140;
  wire popcount45_dokv_core_143;
  wire popcount45_dokv_core_144;
  wire popcount45_dokv_core_145;
  wire popcount45_dokv_core_146;
  wire popcount45_dokv_core_148;
  wire popcount45_dokv_core_149;
  wire popcount45_dokv_core_151;
  wire popcount45_dokv_core_153;
  wire popcount45_dokv_core_154;
  wire popcount45_dokv_core_158;
  wire popcount45_dokv_core_159;
  wire popcount45_dokv_core_160;
  wire popcount45_dokv_core_162;
  wire popcount45_dokv_core_163;
  wire popcount45_dokv_core_164;
  wire popcount45_dokv_core_166;
  wire popcount45_dokv_core_167_not;
  wire popcount45_dokv_core_168;
  wire popcount45_dokv_core_170;
  wire popcount45_dokv_core_173;
  wire popcount45_dokv_core_174;
  wire popcount45_dokv_core_175;
  wire popcount45_dokv_core_176;
  wire popcount45_dokv_core_177;
  wire popcount45_dokv_core_178;
  wire popcount45_dokv_core_179;
  wire popcount45_dokv_core_181;
  wire popcount45_dokv_core_182;
  wire popcount45_dokv_core_183;
  wire popcount45_dokv_core_184;
  wire popcount45_dokv_core_185;
  wire popcount45_dokv_core_186;
  wire popcount45_dokv_core_188;
  wire popcount45_dokv_core_189;
  wire popcount45_dokv_core_190;
  wire popcount45_dokv_core_191;
  wire popcount45_dokv_core_192;
  wire popcount45_dokv_core_193;
  wire popcount45_dokv_core_196;
  wire popcount45_dokv_core_197;
  wire popcount45_dokv_core_201;
  wire popcount45_dokv_core_203;
  wire popcount45_dokv_core_206;
  wire popcount45_dokv_core_207;
  wire popcount45_dokv_core_209;
  wire popcount45_dokv_core_210;
  wire popcount45_dokv_core_214;
  wire popcount45_dokv_core_215;
  wire popcount45_dokv_core_217;
  wire popcount45_dokv_core_218;
  wire popcount45_dokv_core_221;
  wire popcount45_dokv_core_223_not;
  wire popcount45_dokv_core_224;
  wire popcount45_dokv_core_225;
  wire popcount45_dokv_core_227;
  wire popcount45_dokv_core_229;
  wire popcount45_dokv_core_231;
  wire popcount45_dokv_core_232_not;
  wire popcount45_dokv_core_235;
  wire popcount45_dokv_core_236;
  wire popcount45_dokv_core_237;
  wire popcount45_dokv_core_239;
  wire popcount45_dokv_core_240;
  wire popcount45_dokv_core_243;
  wire popcount45_dokv_core_244;
  wire popcount45_dokv_core_245;
  wire popcount45_dokv_core_246;
  wire popcount45_dokv_core_247;
  wire popcount45_dokv_core_248_not;
  wire popcount45_dokv_core_249;
  wire popcount45_dokv_core_250;
  wire popcount45_dokv_core_251;
  wire popcount45_dokv_core_253;
  wire popcount45_dokv_core_254;
  wire popcount45_dokv_core_257;
  wire popcount45_dokv_core_258;
  wire popcount45_dokv_core_259;
  wire popcount45_dokv_core_263;
  wire popcount45_dokv_core_265;
  wire popcount45_dokv_core_267;
  wire popcount45_dokv_core_269;
  wire popcount45_dokv_core_276;
  wire popcount45_dokv_core_277;
  wire popcount45_dokv_core_278;
  wire popcount45_dokv_core_280;
  wire popcount45_dokv_core_281;
  wire popcount45_dokv_core_282;
  wire popcount45_dokv_core_283;
  wire popcount45_dokv_core_286;
  wire popcount45_dokv_core_287;
  wire popcount45_dokv_core_288;
  wire popcount45_dokv_core_290;
  wire popcount45_dokv_core_291;
  wire popcount45_dokv_core_292;
  wire popcount45_dokv_core_294;
  wire popcount45_dokv_core_295;
  wire popcount45_dokv_core_296;
  wire popcount45_dokv_core_297;
  wire popcount45_dokv_core_299;
  wire popcount45_dokv_core_300;
  wire popcount45_dokv_core_302;
  wire popcount45_dokv_core_304;
  wire popcount45_dokv_core_307;
  wire popcount45_dokv_core_308;
  wire popcount45_dokv_core_310;
  wire popcount45_dokv_core_311;
  wire popcount45_dokv_core_312;
  wire popcount45_dokv_core_313;
  wire popcount45_dokv_core_315;
  wire popcount45_dokv_core_316;
  wire popcount45_dokv_core_317;
  wire popcount45_dokv_core_318;
  wire popcount45_dokv_core_319;
  wire popcount45_dokv_core_321;
  wire popcount45_dokv_core_322;
  wire popcount45_dokv_core_326;
  wire popcount45_dokv_core_328;
  wire popcount45_dokv_core_329;
  wire popcount45_dokv_core_330;
  wire popcount45_dokv_core_332;
  wire popcount45_dokv_core_333;
  wire popcount45_dokv_core_334;
  wire popcount45_dokv_core_335;
  wire popcount45_dokv_core_336;
  wire popcount45_dokv_core_337;
  wire popcount45_dokv_core_341;
  wire popcount45_dokv_core_342;
  wire popcount45_dokv_core_344;
  wire popcount45_dokv_core_346;
  wire popcount45_dokv_core_348;
  wire popcount45_dokv_core_349;
  wire popcount45_dokv_core_350;
  wire popcount45_dokv_core_351;
  wire popcount45_dokv_core_352;
  wire popcount45_dokv_core_353;
  wire popcount45_dokv_core_356;

  assign popcount45_dokv_core_049 = input_a[34] & input_a[34];
  assign popcount45_dokv_core_051 = ~input_a[23];
  assign popcount45_dokv_core_052 = input_a[36] | input_a[11];
  assign popcount45_dokv_core_054 = input_a[30] & input_a[10];
  assign popcount45_dokv_core_055 = input_a[2] | input_a[29];
  assign popcount45_dokv_core_056 = input_a[12] ^ input_a[28];
  assign popcount45_dokv_core_057 = input_a[31] & input_a[33];
  assign popcount45_dokv_core_059 = input_a[25] & input_a[19];
  assign popcount45_dokv_core_061 = ~input_a[17];
  assign popcount45_dokv_core_062 = ~(input_a[1] ^ input_a[44]);
  assign popcount45_dokv_core_063 = ~(input_a[10] | input_a[18]);
  assign popcount45_dokv_core_064 = input_a[44] | input_a[43];
  assign popcount45_dokv_core_065 = input_a[39] ^ input_a[24];
  assign popcount45_dokv_core_066 = input_a[26] & input_a[24];
  assign popcount45_dokv_core_068 = ~(input_a[18] | input_a[37]);
  assign popcount45_dokv_core_071 = ~(input_a[26] | input_a[41]);
  assign popcount45_dokv_core_072 = ~input_a[43];
  assign popcount45_dokv_core_073 = ~(input_a[36] & input_a[38]);
  assign popcount45_dokv_core_075 = input_a[4] ^ input_a[22];
  assign popcount45_dokv_core_076 = ~(input_a[7] | input_a[35]);
  assign popcount45_dokv_core_077 = input_a[38] | input_a[30];
  assign popcount45_dokv_core_078 = input_a[14] & input_a[21];
  assign popcount45_dokv_core_079 = ~(input_a[11] ^ input_a[26]);
  assign popcount45_dokv_core_081 = input_a[2] & input_a[0];
  assign popcount45_dokv_core_083_not = ~input_a[24];
  assign popcount45_dokv_core_085 = ~(input_a[33] & input_a[23]);
  assign popcount45_dokv_core_086 = input_a[33] | input_a[31];
  assign popcount45_dokv_core_087 = input_a[36] & input_a[0];
  assign popcount45_dokv_core_089 = ~(input_a[10] ^ input_a[5]);
  assign popcount45_dokv_core_090 = ~(input_a[36] & input_a[33]);
  assign popcount45_dokv_core_092 = input_a[26] & input_a[16];
  assign popcount45_dokv_core_093 = ~(input_a[34] & input_a[37]);
  assign popcount45_dokv_core_094 = input_a[9] & input_a[36];
  assign popcount45_dokv_core_096 = input_a[20] ^ input_a[14];
  assign popcount45_dokv_core_098 = ~(input_a[5] & input_a[5]);
  assign popcount45_dokv_core_101 = ~(input_a[26] ^ input_a[33]);
  assign popcount45_dokv_core_102 = ~input_a[2];
  assign popcount45_dokv_core_104 = input_a[8] & input_a[16];
  assign popcount45_dokv_core_105 = ~(input_a[43] & input_a[32]);
  assign popcount45_dokv_core_106 = ~(input_a[2] | input_a[13]);
  assign popcount45_dokv_core_107 = ~(input_a[33] | input_a[39]);
  assign popcount45_dokv_core_108 = input_a[10] & input_a[20];
  assign popcount45_dokv_core_113 = ~(input_a[5] ^ input_a[5]);
  assign popcount45_dokv_core_114 = ~(input_a[15] | input_a[38]);
  assign popcount45_dokv_core_116 = input_a[24] | input_a[5];
  assign popcount45_dokv_core_117 = input_a[13] & input_a[12];
  assign popcount45_dokv_core_118 = ~(input_a[7] | input_a[32]);
  assign popcount45_dokv_core_121 = ~(input_a[35] ^ input_a[39]);
  assign popcount45_dokv_core_126 = ~(input_a[44] ^ input_a[19]);
  assign popcount45_dokv_core_127 = input_a[32] & input_a[12];
  assign popcount45_dokv_core_128 = input_a[19] ^ input_a[7];
  assign popcount45_dokv_core_129 = input_a[19] ^ input_a[32];
  assign popcount45_dokv_core_130 = input_a[8] & input_a[32];
  assign popcount45_dokv_core_131_not = ~input_a[13];
  assign popcount45_dokv_core_133 = input_a[33] ^ input_a[7];
  assign popcount45_dokv_core_134 = input_a[3] & input_a[16];
  assign popcount45_dokv_core_135 = ~input_a[40];
  assign popcount45_dokv_core_137 = ~(input_a[0] ^ input_a[31]);
  assign popcount45_dokv_core_139 = ~(input_a[7] ^ input_a[37]);
  assign popcount45_dokv_core_140 = input_a[36] | input_a[14];
  assign popcount45_dokv_core_143 = input_a[14] ^ input_a[10];
  assign popcount45_dokv_core_144 = ~(input_a[21] & input_a[20]);
  assign popcount45_dokv_core_145 = input_a[4] | input_a[3];
  assign popcount45_dokv_core_146 = input_a[31] | input_a[44];
  assign popcount45_dokv_core_148 = input_a[26] | input_a[1];
  assign popcount45_dokv_core_149 = ~(input_a[20] | input_a[21]);
  assign popcount45_dokv_core_151 = input_a[0] ^ input_a[0];
  assign popcount45_dokv_core_153 = ~(input_a[7] | input_a[28]);
  assign popcount45_dokv_core_154 = ~input_a[9];
  assign popcount45_dokv_core_158 = ~(input_a[14] & input_a[6]);
  assign popcount45_dokv_core_159 = ~(input_a[36] ^ input_a[30]);
  assign popcount45_dokv_core_160 = ~(input_a[23] | input_a[33]);
  assign popcount45_dokv_core_162 = ~(input_a[9] | input_a[43]);
  assign popcount45_dokv_core_163 = input_a[18] | input_a[25];
  assign popcount45_dokv_core_164 = input_a[2] | input_a[0];
  assign popcount45_dokv_core_166 = input_a[4] & input_a[21];
  assign popcount45_dokv_core_167_not = ~input_a[19];
  assign popcount45_dokv_core_168 = ~(input_a[39] & input_a[39]);
  assign popcount45_dokv_core_170 = ~(input_a[10] | input_a[38]);
  assign popcount45_dokv_core_173 = input_a[21] ^ input_a[16];
  assign popcount45_dokv_core_174 = input_a[5] | input_a[42];
  assign popcount45_dokv_core_175 = input_a[11] & input_a[27];
  assign popcount45_dokv_core_176 = ~input_a[23];
  assign popcount45_dokv_core_177 = input_a[16] | input_a[8];
  assign popcount45_dokv_core_178 = ~input_a[8];
  assign popcount45_dokv_core_179 = input_a[1] ^ input_a[10];
  assign popcount45_dokv_core_181 = ~(input_a[3] ^ input_a[22]);
  assign popcount45_dokv_core_182 = ~input_a[29];
  assign popcount45_dokv_core_183 = ~(input_a[23] & input_a[18]);
  assign popcount45_dokv_core_184 = input_a[40] ^ input_a[3];
  assign popcount45_dokv_core_185 = ~(input_a[38] & input_a[15]);
  assign popcount45_dokv_core_186 = ~(input_a[8] ^ input_a[1]);
  assign popcount45_dokv_core_188 = ~(input_a[2] | input_a[42]);
  assign popcount45_dokv_core_189 = input_a[30] | input_a[26];
  assign popcount45_dokv_core_190 = ~input_a[23];
  assign popcount45_dokv_core_191 = ~(input_a[18] | input_a[44]);
  assign popcount45_dokv_core_192 = input_a[5] & input_a[28];
  assign popcount45_dokv_core_193 = ~input_a[27];
  assign popcount45_dokv_core_196 = input_a[4] | input_a[35];
  assign popcount45_dokv_core_197 = ~(input_a[30] & input_a[40]);
  assign popcount45_dokv_core_201 = input_a[8] ^ input_a[5];
  assign popcount45_dokv_core_203 = ~input_a[13];
  assign popcount45_dokv_core_206 = input_a[16] ^ input_a[11];
  assign popcount45_dokv_core_207 = ~(input_a[10] | input_a[18]);
  assign popcount45_dokv_core_209 = ~(input_a[43] ^ input_a[28]);
  assign popcount45_dokv_core_210 = input_a[24] | input_a[39];
  assign popcount45_dokv_core_214 = ~(input_a[14] & input_a[31]);
  assign popcount45_dokv_core_215 = ~input_a[30];
  assign popcount45_dokv_core_217 = ~(input_a[19] ^ input_a[36]);
  assign popcount45_dokv_core_218 = ~(input_a[30] | input_a[39]);
  assign popcount45_dokv_core_221 = ~(input_a[10] ^ input_a[26]);
  assign popcount45_dokv_core_223_not = ~input_a[32];
  assign popcount45_dokv_core_224 = input_a[30] | input_a[2];
  assign popcount45_dokv_core_225 = input_a[43] & input_a[18];
  assign popcount45_dokv_core_227 = ~(input_a[9] ^ input_a[30]);
  assign popcount45_dokv_core_229 = ~(input_a[30] & input_a[42]);
  assign popcount45_dokv_core_231 = ~(input_a[23] & input_a[16]);
  assign popcount45_dokv_core_232_not = ~input_a[7];
  assign popcount45_dokv_core_235 = ~(input_a[41] & input_a[28]);
  assign popcount45_dokv_core_236 = input_a[8] ^ input_a[34];
  assign popcount45_dokv_core_237 = ~(input_a[1] ^ input_a[34]);
  assign popcount45_dokv_core_239 = input_a[24] | input_a[42];
  assign popcount45_dokv_core_240 = ~(input_a[14] | input_a[40]);
  assign popcount45_dokv_core_243 = ~(input_a[8] ^ input_a[23]);
  assign popcount45_dokv_core_244 = input_a[11] | input_a[29];
  assign popcount45_dokv_core_245 = ~(input_a[25] & input_a[13]);
  assign popcount45_dokv_core_246 = ~input_a[21];
  assign popcount45_dokv_core_247 = ~(input_a[38] ^ input_a[5]);
  assign popcount45_dokv_core_248_not = ~input_a[44];
  assign popcount45_dokv_core_249 = ~input_a[44];
  assign popcount45_dokv_core_250 = ~input_a[5];
  assign popcount45_dokv_core_251 = ~(input_a[14] ^ input_a[1]);
  assign popcount45_dokv_core_253 = input_a[20] | input_a[7];
  assign popcount45_dokv_core_254 = ~(input_a[44] & input_a[39]);
  assign popcount45_dokv_core_257 = ~(input_a[14] ^ input_a[21]);
  assign popcount45_dokv_core_258 = input_a[6] & input_a[11];
  assign popcount45_dokv_core_259 = input_a[30] & input_a[35];
  assign popcount45_dokv_core_263 = input_a[31] ^ input_a[37];
  assign popcount45_dokv_core_265 = ~(input_a[25] ^ input_a[31]);
  assign popcount45_dokv_core_267 = input_a[28] ^ input_a[12];
  assign popcount45_dokv_core_269 = input_a[3] ^ input_a[12];
  assign popcount45_dokv_core_276 = ~(input_a[27] | input_a[36]);
  assign popcount45_dokv_core_277 = ~(input_a[37] ^ input_a[19]);
  assign popcount45_dokv_core_278 = ~input_a[19];
  assign popcount45_dokv_core_280 = ~(input_a[24] ^ input_a[13]);
  assign popcount45_dokv_core_281 = ~(input_a[22] & input_a[13]);
  assign popcount45_dokv_core_282 = ~(input_a[16] ^ input_a[25]);
  assign popcount45_dokv_core_283 = ~(input_a[17] ^ input_a[34]);
  assign popcount45_dokv_core_286 = ~(input_a[12] & input_a[22]);
  assign popcount45_dokv_core_287 = ~(input_a[14] | input_a[40]);
  assign popcount45_dokv_core_288 = input_a[32] | input_a[24];
  assign popcount45_dokv_core_290 = ~(input_a[29] | input_a[35]);
  assign popcount45_dokv_core_291 = input_a[30] & input_a[38];
  assign popcount45_dokv_core_292 = ~(input_a[38] & input_a[41]);
  assign popcount45_dokv_core_294 = input_a[10] & input_a[5];
  assign popcount45_dokv_core_295 = ~input_a[18];
  assign popcount45_dokv_core_296 = input_a[10] ^ input_a[10];
  assign popcount45_dokv_core_297 = input_a[29] | input_a[34];
  assign popcount45_dokv_core_299 = ~input_a[37];
  assign popcount45_dokv_core_300 = ~(input_a[7] ^ input_a[6]);
  assign popcount45_dokv_core_302 = ~(input_a[3] ^ input_a[19]);
  assign popcount45_dokv_core_304 = input_a[25] | input_a[37];
  assign popcount45_dokv_core_307 = ~(input_a[4] ^ input_a[5]);
  assign popcount45_dokv_core_308 = ~input_a[25];
  assign popcount45_dokv_core_310 = input_a[29] ^ input_a[43];
  assign popcount45_dokv_core_311 = ~input_a[40];
  assign popcount45_dokv_core_312 = input_a[35] | input_a[16];
  assign popcount45_dokv_core_313 = ~(input_a[43] & input_a[39]);
  assign popcount45_dokv_core_315 = input_a[27] | input_a[38];
  assign popcount45_dokv_core_316 = ~(input_a[38] & input_a[19]);
  assign popcount45_dokv_core_317 = ~input_a[37];
  assign popcount45_dokv_core_318 = ~(input_a[0] & input_a[27]);
  assign popcount45_dokv_core_319 = ~(input_a[18] | input_a[19]);
  assign popcount45_dokv_core_321 = ~(input_a[18] | input_a[29]);
  assign popcount45_dokv_core_322 = input_a[1] ^ input_a[4];
  assign popcount45_dokv_core_326 = input_a[22] | input_a[38];
  assign popcount45_dokv_core_328 = ~input_a[9];
  assign popcount45_dokv_core_329 = ~(input_a[1] & input_a[5]);
  assign popcount45_dokv_core_330 = ~(input_a[29] ^ input_a[10]);
  assign popcount45_dokv_core_332 = ~(input_a[22] | input_a[1]);
  assign popcount45_dokv_core_333 = input_a[40] & input_a[15];
  assign popcount45_dokv_core_334 = ~(input_a[3] & input_a[17]);
  assign popcount45_dokv_core_335 = input_a[41] & input_a[11];
  assign popcount45_dokv_core_336 = ~(input_a[28] & input_a[21]);
  assign popcount45_dokv_core_337 = input_a[17] ^ input_a[8];
  assign popcount45_dokv_core_341 = input_a[38] ^ input_a[18];
  assign popcount45_dokv_core_342 = input_a[30] ^ input_a[38];
  assign popcount45_dokv_core_344 = ~(input_a[19] ^ input_a[22]);
  assign popcount45_dokv_core_346 = ~input_a[2];
  assign popcount45_dokv_core_348 = input_a[42] ^ input_a[15];
  assign popcount45_dokv_core_349 = ~(input_a[15] & input_a[21]);
  assign popcount45_dokv_core_350 = ~(input_a[20] & input_a[32]);
  assign popcount45_dokv_core_351 = input_a[33] & input_a[2];
  assign popcount45_dokv_core_352 = ~(input_a[13] | input_a[33]);
  assign popcount45_dokv_core_353 = ~(input_a[10] & input_a[37]);
  assign popcount45_dokv_core_356 = ~(input_a[5] | input_a[32]);

  assign popcount45_dokv_out[0] = 1'b1;
  assign popcount45_dokv_out[1] = input_a[28];
  assign popcount45_dokv_out[2] = input_a[43];
  assign popcount45_dokv_out[3] = 1'b0;
  assign popcount45_dokv_out[4] = 1'b1;
  assign popcount45_dokv_out[5] = 1'b0;
endmodule