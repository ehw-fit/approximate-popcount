// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.6455
// WCE=14.0
// EP=0.810121%
// Printed PDK parameters:
//  Area=40907854.0
//  Delay=59913064.0
//  Power=2066300.0

module popcount33_w90i(input [32:0] input_a, output [5:0] popcount33_w90i_out);
  wire popcount33_w90i_core_036;
  wire popcount33_w90i_core_037;
  wire popcount33_w90i_core_038;
  wire popcount33_w90i_core_039;
  wire popcount33_w90i_core_040;
  wire popcount33_w90i_core_042;
  wire popcount33_w90i_core_044;
  wire popcount33_w90i_core_045;
  wire popcount33_w90i_core_046;
  wire popcount33_w90i_core_047;
  wire popcount33_w90i_core_048;
  wire popcount33_w90i_core_049;
  wire popcount33_w90i_core_050;
  wire popcount33_w90i_core_051;
  wire popcount33_w90i_core_052;
  wire popcount33_w90i_core_053;
  wire popcount33_w90i_core_055;
  wire popcount33_w90i_core_056;
  wire popcount33_w90i_core_057;
  wire popcount33_w90i_core_058;
  wire popcount33_w90i_core_059_not;
  wire popcount33_w90i_core_061;
  wire popcount33_w90i_core_062;
  wire popcount33_w90i_core_063;
  wire popcount33_w90i_core_065;
  wire popcount33_w90i_core_066;
  wire popcount33_w90i_core_067;
  wire popcount33_w90i_core_068;
  wire popcount33_w90i_core_069;
  wire popcount33_w90i_core_070;
  wire popcount33_w90i_core_071;
  wire popcount33_w90i_core_073;
  wire popcount33_w90i_core_075;
  wire popcount33_w90i_core_076;
  wire popcount33_w90i_core_077;
  wire popcount33_w90i_core_078;
  wire popcount33_w90i_core_079;
  wire popcount33_w90i_core_080;
  wire popcount33_w90i_core_081;
  wire popcount33_w90i_core_082;
  wire popcount33_w90i_core_083;
  wire popcount33_w90i_core_086;
  wire popcount33_w90i_core_088;
  wire popcount33_w90i_core_089;
  wire popcount33_w90i_core_091;
  wire popcount33_w90i_core_092;
  wire popcount33_w90i_core_093;
  wire popcount33_w90i_core_094;
  wire popcount33_w90i_core_095;
  wire popcount33_w90i_core_096;
  wire popcount33_w90i_core_097;
  wire popcount33_w90i_core_099;
  wire popcount33_w90i_core_100;
  wire popcount33_w90i_core_102;
  wire popcount33_w90i_core_104;
  wire popcount33_w90i_core_105;
  wire popcount33_w90i_core_106;
  wire popcount33_w90i_core_107;
  wire popcount33_w90i_core_108;
  wire popcount33_w90i_core_109;
  wire popcount33_w90i_core_112_not;
  wire popcount33_w90i_core_116;
  wire popcount33_w90i_core_118;
  wire popcount33_w90i_core_123;
  wire popcount33_w90i_core_124;
  wire popcount33_w90i_core_125;
  wire popcount33_w90i_core_126;
  wire popcount33_w90i_core_127;
  wire popcount33_w90i_core_129;
  wire popcount33_w90i_core_131;
  wire popcount33_w90i_core_133;
  wire popcount33_w90i_core_134;
  wire popcount33_w90i_core_135;
  wire popcount33_w90i_core_137;
  wire popcount33_w90i_core_138;
  wire popcount33_w90i_core_140;
  wire popcount33_w90i_core_142;
  wire popcount33_w90i_core_143;
  wire popcount33_w90i_core_144;
  wire popcount33_w90i_core_145;
  wire popcount33_w90i_core_146;
  wire popcount33_w90i_core_147;
  wire popcount33_w90i_core_148;
  wire popcount33_w90i_core_149;
  wire popcount33_w90i_core_150;
  wire popcount33_w90i_core_151;
  wire popcount33_w90i_core_152;
  wire popcount33_w90i_core_153;
  wire popcount33_w90i_core_154;
  wire popcount33_w90i_core_155;
  wire popcount33_w90i_core_157;
  wire popcount33_w90i_core_160;
  wire popcount33_w90i_core_161;
  wire popcount33_w90i_core_162;
  wire popcount33_w90i_core_163;
  wire popcount33_w90i_core_165;
  wire popcount33_w90i_core_166;
  wire popcount33_w90i_core_167;
  wire popcount33_w90i_core_168;
  wire popcount33_w90i_core_169;
  wire popcount33_w90i_core_172;
  wire popcount33_w90i_core_174;
  wire popcount33_w90i_core_175;
  wire popcount33_w90i_core_176;
  wire popcount33_w90i_core_179;
  wire popcount33_w90i_core_180;
  wire popcount33_w90i_core_182_not;
  wire popcount33_w90i_core_183;
  wire popcount33_w90i_core_184;
  wire popcount33_w90i_core_185;
  wire popcount33_w90i_core_186;
  wire popcount33_w90i_core_187;
  wire popcount33_w90i_core_188;
  wire popcount33_w90i_core_190_not;
  wire popcount33_w90i_core_191;
  wire popcount33_w90i_core_192_not;
  wire popcount33_w90i_core_193;
  wire popcount33_w90i_core_194;
  wire popcount33_w90i_core_198;
  wire popcount33_w90i_core_199;
  wire popcount33_w90i_core_203;
  wire popcount33_w90i_core_204;
  wire popcount33_w90i_core_205;
  wire popcount33_w90i_core_206;
  wire popcount33_w90i_core_207;
  wire popcount33_w90i_core_209;
  wire popcount33_w90i_core_210;
  wire popcount33_w90i_core_212;
  wire popcount33_w90i_core_213;
  wire popcount33_w90i_core_215;
  wire popcount33_w90i_core_216;
  wire popcount33_w90i_core_217;
  wire popcount33_w90i_core_218;
  wire popcount33_w90i_core_219;
  wire popcount33_w90i_core_220;
  wire popcount33_w90i_core_221;
  wire popcount33_w90i_core_222;
  wire popcount33_w90i_core_223;
  wire popcount33_w90i_core_224;
  wire popcount33_w90i_core_225;
  wire popcount33_w90i_core_226;
  wire popcount33_w90i_core_227;
  wire popcount33_w90i_core_228;
  wire popcount33_w90i_core_229;
  wire popcount33_w90i_core_230;
  wire popcount33_w90i_core_231;
  wire popcount33_w90i_core_233;
  wire popcount33_w90i_core_237;

  assign popcount33_w90i_core_036 = ~(input_a[15] | input_a[19]);
  assign popcount33_w90i_core_037 = ~(input_a[5] & input_a[22]);
  assign popcount33_w90i_core_038 = ~(input_a[16] & input_a[22]);
  assign popcount33_w90i_core_039 = ~(input_a[4] ^ input_a[6]);
  assign popcount33_w90i_core_040 = ~(input_a[18] & input_a[10]);
  assign popcount33_w90i_core_042 = ~(input_a[29] | input_a[27]);
  assign popcount33_w90i_core_044 = input_a[28] | input_a[23];
  assign popcount33_w90i_core_045 = ~(input_a[4] | input_a[30]);
  assign popcount33_w90i_core_046 = ~(input_a[6] & input_a[10]);
  assign popcount33_w90i_core_047 = input_a[12] ^ input_a[0];
  assign popcount33_w90i_core_048 = ~input_a[12];
  assign popcount33_w90i_core_049 = ~(input_a[23] ^ input_a[4]);
  assign popcount33_w90i_core_050 = ~(popcount33_w90i_core_046 & popcount33_w90i_core_048);
  assign popcount33_w90i_core_051 = input_a[6] ^ input_a[29];
  assign popcount33_w90i_core_052 = ~(input_a[27] & input_a[29]);
  assign popcount33_w90i_core_053 = ~(input_a[26] | input_a[7]);
  assign popcount33_w90i_core_055 = input_a[29] & input_a[20];
  assign popcount33_w90i_core_056 = ~input_a[23];
  assign popcount33_w90i_core_057 = ~(input_a[29] | input_a[17]);
  assign popcount33_w90i_core_058 = input_a[26] & popcount33_w90i_core_050;
  assign popcount33_w90i_core_059_not = ~popcount33_w90i_core_052;
  assign popcount33_w90i_core_061 = popcount33_w90i_core_059_not | popcount33_w90i_core_058;
  assign popcount33_w90i_core_062 = input_a[22] | input_a[24];
  assign popcount33_w90i_core_063 = ~(input_a[32] & input_a[20]);
  assign popcount33_w90i_core_065 = ~input_a[4];
  assign popcount33_w90i_core_066 = input_a[19] ^ input_a[18];
  assign popcount33_w90i_core_067 = input_a[9] ^ input_a[31];
  assign popcount33_w90i_core_068 = ~input_a[9];
  assign popcount33_w90i_core_069 = ~(input_a[26] | input_a[26]);
  assign popcount33_w90i_core_070 = ~(input_a[26] | input_a[27]);
  assign popcount33_w90i_core_071 = input_a[21] & input_a[19];
  assign popcount33_w90i_core_073 = input_a[24] & input_a[19];
  assign popcount33_w90i_core_075 = input_a[20] | input_a[20];
  assign popcount33_w90i_core_076 = ~input_a[8];
  assign popcount33_w90i_core_077 = input_a[22] ^ input_a[26];
  assign popcount33_w90i_core_078 = ~(input_a[23] ^ input_a[32]);
  assign popcount33_w90i_core_079 = ~(input_a[8] & input_a[20]);
  assign popcount33_w90i_core_080 = ~(input_a[25] | input_a[30]);
  assign popcount33_w90i_core_081 = input_a[20] | input_a[16];
  assign popcount33_w90i_core_082 = input_a[10] | input_a[24];
  assign popcount33_w90i_core_083 = ~(input_a[18] ^ input_a[0]);
  assign popcount33_w90i_core_086 = ~input_a[31];
  assign popcount33_w90i_core_088 = input_a[14] & input_a[22];
  assign popcount33_w90i_core_089 = ~(input_a[4] ^ input_a[29]);
  assign popcount33_w90i_core_091 = ~(input_a[4] ^ input_a[16]);
  assign popcount33_w90i_core_092 = input_a[20] & input_a[30];
  assign popcount33_w90i_core_093 = ~(input_a[4] & input_a[3]);
  assign popcount33_w90i_core_094 = ~(input_a[25] & input_a[3]);
  assign popcount33_w90i_core_095 = input_a[4] | input_a[8];
  assign popcount33_w90i_core_096 = input_a[6] & input_a[8];
  assign popcount33_w90i_core_097 = input_a[22] & input_a[1];
  assign popcount33_w90i_core_099 = input_a[24] ^ input_a[15];
  assign popcount33_w90i_core_100 = ~(input_a[5] & input_a[3]);
  assign popcount33_w90i_core_102 = ~input_a[13];
  assign popcount33_w90i_core_104 = input_a[28] | input_a[5];
  assign popcount33_w90i_core_105 = popcount33_w90i_core_061 ^ popcount33_w90i_core_095;
  assign popcount33_w90i_core_106 = popcount33_w90i_core_061 & popcount33_w90i_core_095;
  assign popcount33_w90i_core_107 = popcount33_w90i_core_105 ^ input_a[13];
  assign popcount33_w90i_core_108 = popcount33_w90i_core_105 & input_a[13];
  assign popcount33_w90i_core_109 = popcount33_w90i_core_106 | popcount33_w90i_core_108;
  assign popcount33_w90i_core_112_not = ~popcount33_w90i_core_109;
  assign popcount33_w90i_core_116 = ~(input_a[1] ^ input_a[29]);
  assign popcount33_w90i_core_118 = ~(input_a[23] & input_a[18]);
  assign popcount33_w90i_core_123 = input_a[0] & input_a[32];
  assign popcount33_w90i_core_124 = input_a[3] | input_a[14];
  assign popcount33_w90i_core_125 = input_a[31] & input_a[32];
  assign popcount33_w90i_core_126 = input_a[16] ^ popcount33_w90i_core_123;
  assign popcount33_w90i_core_127 = input_a[16] & popcount33_w90i_core_123;
  assign popcount33_w90i_core_129 = ~input_a[0];
  assign popcount33_w90i_core_131 = ~(input_a[19] | input_a[30]);
  assign popcount33_w90i_core_133 = input_a[12] & input_a[2];
  assign popcount33_w90i_core_134 = input_a[0] & input_a[16];
  assign popcount33_w90i_core_135 = ~popcount33_w90i_core_131;
  assign popcount33_w90i_core_137 = ~(input_a[23] & input_a[1]);
  assign popcount33_w90i_core_138 = input_a[23] & input_a[1];
  assign popcount33_w90i_core_140 = ~(input_a[18] & input_a[11]);
  assign popcount33_w90i_core_142 = input_a[21] ^ input_a[6];
  assign popcount33_w90i_core_143 = popcount33_w90i_core_124 & popcount33_w90i_core_135;
  assign popcount33_w90i_core_144 = popcount33_w90i_core_126 ^ popcount33_w90i_core_137;
  assign popcount33_w90i_core_145 = popcount33_w90i_core_126 & popcount33_w90i_core_137;
  assign popcount33_w90i_core_146 = popcount33_w90i_core_144 ^ popcount33_w90i_core_143;
  assign popcount33_w90i_core_147 = popcount33_w90i_core_144 & popcount33_w90i_core_143;
  assign popcount33_w90i_core_148 = popcount33_w90i_core_145 | popcount33_w90i_core_147;
  assign popcount33_w90i_core_149 = popcount33_w90i_core_127 ^ popcount33_w90i_core_138;
  assign popcount33_w90i_core_150 = popcount33_w90i_core_127 & popcount33_w90i_core_138;
  assign popcount33_w90i_core_151 = popcount33_w90i_core_149 ^ popcount33_w90i_core_148;
  assign popcount33_w90i_core_152 = popcount33_w90i_core_149 & popcount33_w90i_core_148;
  assign popcount33_w90i_core_153 = popcount33_w90i_core_150 | popcount33_w90i_core_152;
  assign popcount33_w90i_core_154 = input_a[24] ^ input_a[25];
  assign popcount33_w90i_core_155 = input_a[24] & input_a[25];
  assign popcount33_w90i_core_157 = input_a[7] & input_a[15];
  assign popcount33_w90i_core_160 = input_a[25] ^ popcount33_w90i_core_157;
  assign popcount33_w90i_core_161 = popcount33_w90i_core_155 & popcount33_w90i_core_157;
  assign popcount33_w90i_core_162 = popcount33_w90i_core_160 | popcount33_w90i_core_154;
  assign popcount33_w90i_core_163 = input_a[2] | input_a[18];
  assign popcount33_w90i_core_165 = input_a[6] | input_a[10];
  assign popcount33_w90i_core_166 = input_a[9] & input_a[28];
  assign popcount33_w90i_core_167 = input_a[11] ^ input_a[10];
  assign popcount33_w90i_core_168 = input_a[17] & input_a[20];
  assign popcount33_w90i_core_169 = ~(input_a[0] | input_a[17]);
  assign popcount33_w90i_core_172 = input_a[32] | input_a[23];
  assign popcount33_w90i_core_174 = ~(input_a[20] ^ input_a[10]);
  assign popcount33_w90i_core_175 = popcount33_w90i_core_166 | popcount33_w90i_core_168;
  assign popcount33_w90i_core_176 = ~input_a[10];
  assign popcount33_w90i_core_179 = ~(input_a[7] ^ input_a[2]);
  assign popcount33_w90i_core_180 = ~input_a[6];
  assign popcount33_w90i_core_182_not = ~input_a[13];
  assign popcount33_w90i_core_183 = input_a[18] & input_a[11];
  assign popcount33_w90i_core_184 = popcount33_w90i_core_162 ^ popcount33_w90i_core_175;
  assign popcount33_w90i_core_185 = popcount33_w90i_core_162 & popcount33_w90i_core_175;
  assign popcount33_w90i_core_186 = popcount33_w90i_core_184 ^ popcount33_w90i_core_183;
  assign popcount33_w90i_core_187 = popcount33_w90i_core_184 & popcount33_w90i_core_183;
  assign popcount33_w90i_core_188 = popcount33_w90i_core_185 | popcount33_w90i_core_187;
  assign popcount33_w90i_core_190_not = ~input_a[28];
  assign popcount33_w90i_core_191 = popcount33_w90i_core_161 | popcount33_w90i_core_188;
  assign popcount33_w90i_core_192_not = ~input_a[28];
  assign popcount33_w90i_core_193 = ~input_a[23];
  assign popcount33_w90i_core_194 = input_a[6] | input_a[14];
  assign popcount33_w90i_core_198 = popcount33_w90i_core_146 ^ popcount33_w90i_core_186;
  assign popcount33_w90i_core_199 = popcount33_w90i_core_146 & popcount33_w90i_core_186;
  assign popcount33_w90i_core_203 = popcount33_w90i_core_151 ^ popcount33_w90i_core_191;
  assign popcount33_w90i_core_204 = popcount33_w90i_core_151 & popcount33_w90i_core_191;
  assign popcount33_w90i_core_205 = popcount33_w90i_core_203 ^ popcount33_w90i_core_199;
  assign popcount33_w90i_core_206 = popcount33_w90i_core_203 & popcount33_w90i_core_199;
  assign popcount33_w90i_core_207 = popcount33_w90i_core_204 | popcount33_w90i_core_206;
  assign popcount33_w90i_core_209 = ~input_a[26];
  assign popcount33_w90i_core_210 = popcount33_w90i_core_153 | popcount33_w90i_core_207;
  assign popcount33_w90i_core_212 = ~(input_a[14] & input_a[27]);
  assign popcount33_w90i_core_213 = ~(input_a[20] ^ input_a[1]);
  assign popcount33_w90i_core_215 = input_a[28] ^ input_a[0];
  assign popcount33_w90i_core_216 = input_a[31] & input_a[2];
  assign popcount33_w90i_core_217 = popcount33_w90i_core_107 ^ popcount33_w90i_core_198;
  assign popcount33_w90i_core_218 = popcount33_w90i_core_107 & popcount33_w90i_core_198;
  assign popcount33_w90i_core_219 = popcount33_w90i_core_217 ^ popcount33_w90i_core_216;
  assign popcount33_w90i_core_220 = popcount33_w90i_core_217 & popcount33_w90i_core_216;
  assign popcount33_w90i_core_221 = popcount33_w90i_core_218 | popcount33_w90i_core_220;
  assign popcount33_w90i_core_222 = popcount33_w90i_core_112_not ^ popcount33_w90i_core_205;
  assign popcount33_w90i_core_223 = popcount33_w90i_core_112_not & popcount33_w90i_core_205;
  assign popcount33_w90i_core_224 = popcount33_w90i_core_222 ^ popcount33_w90i_core_221;
  assign popcount33_w90i_core_225 = popcount33_w90i_core_222 & popcount33_w90i_core_221;
  assign popcount33_w90i_core_226 = popcount33_w90i_core_223 | popcount33_w90i_core_225;
  assign popcount33_w90i_core_227 = popcount33_w90i_core_109 ^ popcount33_w90i_core_210;
  assign popcount33_w90i_core_228 = popcount33_w90i_core_109 & popcount33_w90i_core_210;
  assign popcount33_w90i_core_229 = popcount33_w90i_core_227 ^ popcount33_w90i_core_226;
  assign popcount33_w90i_core_230 = popcount33_w90i_core_227 & popcount33_w90i_core_226;
  assign popcount33_w90i_core_231 = popcount33_w90i_core_228 | popcount33_w90i_core_230;
  assign popcount33_w90i_core_233 = ~input_a[18];
  assign popcount33_w90i_core_237 = ~(input_a[1] | input_a[20]);

  assign popcount33_w90i_out[0] = popcount33_w90i_core_229;
  assign popcount33_w90i_out[1] = popcount33_w90i_core_219;
  assign popcount33_w90i_out[2] = popcount33_w90i_core_224;
  assign popcount33_w90i_out[3] = popcount33_w90i_core_229;
  assign popcount33_w90i_out[4] = popcount33_w90i_core_231;
  assign popcount33_w90i_out[5] = 1'b0;
endmodule