// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.76197
// WCE=10.0
// EP=0.823803%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_sqs3(input [20:0] input_a, output [4:0] popcount21_sqs3_out);
  wire popcount21_sqs3_core_024;
  wire popcount21_sqs3_core_025;
  wire popcount21_sqs3_core_029;
  wire popcount21_sqs3_core_030;
  wire popcount21_sqs3_core_032;
  wire popcount21_sqs3_core_033;
  wire popcount21_sqs3_core_034;
  wire popcount21_sqs3_core_036;
  wire popcount21_sqs3_core_037;
  wire popcount21_sqs3_core_039;
  wire popcount21_sqs3_core_040;
  wire popcount21_sqs3_core_043;
  wire popcount21_sqs3_core_044;
  wire popcount21_sqs3_core_047_not;
  wire popcount21_sqs3_core_048;
  wire popcount21_sqs3_core_051;
  wire popcount21_sqs3_core_052;
  wire popcount21_sqs3_core_055;
  wire popcount21_sqs3_core_058;
  wire popcount21_sqs3_core_059;
  wire popcount21_sqs3_core_060;
  wire popcount21_sqs3_core_063;
  wire popcount21_sqs3_core_065;
  wire popcount21_sqs3_core_067;
  wire popcount21_sqs3_core_068;
  wire popcount21_sqs3_core_070;
  wire popcount21_sqs3_core_071;
  wire popcount21_sqs3_core_072;
  wire popcount21_sqs3_core_074;
  wire popcount21_sqs3_core_075;
  wire popcount21_sqs3_core_077;
  wire popcount21_sqs3_core_078;
  wire popcount21_sqs3_core_079;
  wire popcount21_sqs3_core_083;
  wire popcount21_sqs3_core_085;
  wire popcount21_sqs3_core_087;
  wire popcount21_sqs3_core_090;
  wire popcount21_sqs3_core_091;
  wire popcount21_sqs3_core_092;
  wire popcount21_sqs3_core_094;
  wire popcount21_sqs3_core_095;
  wire popcount21_sqs3_core_096;
  wire popcount21_sqs3_core_097;
  wire popcount21_sqs3_core_100;
  wire popcount21_sqs3_core_101;
  wire popcount21_sqs3_core_102;
  wire popcount21_sqs3_core_104;
  wire popcount21_sqs3_core_105;
  wire popcount21_sqs3_core_107;
  wire popcount21_sqs3_core_109;
  wire popcount21_sqs3_core_113;
  wire popcount21_sqs3_core_116;
  wire popcount21_sqs3_core_117;
  wire popcount21_sqs3_core_118;
  wire popcount21_sqs3_core_120;
  wire popcount21_sqs3_core_121;
  wire popcount21_sqs3_core_123;
  wire popcount21_sqs3_core_124;
  wire popcount21_sqs3_core_125;
  wire popcount21_sqs3_core_127;
  wire popcount21_sqs3_core_129;
  wire popcount21_sqs3_core_130;
  wire popcount21_sqs3_core_134;
  wire popcount21_sqs3_core_136;
  wire popcount21_sqs3_core_137;
  wire popcount21_sqs3_core_138;
  wire popcount21_sqs3_core_140;
  wire popcount21_sqs3_core_141;
  wire popcount21_sqs3_core_142;
  wire popcount21_sqs3_core_144;
  wire popcount21_sqs3_core_146;
  wire popcount21_sqs3_core_148;
  wire popcount21_sqs3_core_149;
  wire popcount21_sqs3_core_150;
  wire popcount21_sqs3_core_151;
  wire popcount21_sqs3_core_152;
  wire popcount21_sqs3_core_153;

  assign popcount21_sqs3_core_024 = input_a[6] | input_a[0];
  assign popcount21_sqs3_core_025 = ~input_a[15];
  assign popcount21_sqs3_core_029 = ~(input_a[12] | input_a[17]);
  assign popcount21_sqs3_core_030 = ~(input_a[0] ^ input_a[12]);
  assign popcount21_sqs3_core_032 = input_a[1] | input_a[10];
  assign popcount21_sqs3_core_033 = ~(input_a[1] | input_a[3]);
  assign popcount21_sqs3_core_034 = ~(input_a[3] & input_a[5]);
  assign popcount21_sqs3_core_036 = ~(input_a[13] | input_a[20]);
  assign popcount21_sqs3_core_037 = ~(input_a[11] | input_a[12]);
  assign popcount21_sqs3_core_039 = ~(input_a[17] ^ input_a[13]);
  assign popcount21_sqs3_core_040 = input_a[15] ^ input_a[6];
  assign popcount21_sqs3_core_043 = input_a[18] ^ input_a[20];
  assign popcount21_sqs3_core_044 = ~(input_a[13] & input_a[16]);
  assign popcount21_sqs3_core_047_not = ~input_a[12];
  assign popcount21_sqs3_core_048 = input_a[17] & input_a[6];
  assign popcount21_sqs3_core_051 = ~input_a[1];
  assign popcount21_sqs3_core_052 = input_a[19] & input_a[6];
  assign popcount21_sqs3_core_055 = ~(input_a[10] | input_a[2]);
  assign popcount21_sqs3_core_058 = input_a[7] | input_a[2];
  assign popcount21_sqs3_core_059 = input_a[18] & input_a[2];
  assign popcount21_sqs3_core_060 = ~(input_a[1] & input_a[3]);
  assign popcount21_sqs3_core_063 = input_a[9] ^ input_a[1];
  assign popcount21_sqs3_core_065 = ~(input_a[14] ^ input_a[16]);
  assign popcount21_sqs3_core_067 = ~input_a[7];
  assign popcount21_sqs3_core_068 = input_a[2] | input_a[4];
  assign popcount21_sqs3_core_070 = ~(input_a[14] ^ input_a[10]);
  assign popcount21_sqs3_core_071 = input_a[14] & input_a[18];
  assign popcount21_sqs3_core_072 = input_a[5] & input_a[13];
  assign popcount21_sqs3_core_074 = ~(input_a[17] & input_a[4]);
  assign popcount21_sqs3_core_075 = input_a[4] | input_a[5];
  assign popcount21_sqs3_core_077 = input_a[15] ^ input_a[10];
  assign popcount21_sqs3_core_078 = input_a[8] ^ input_a[11];
  assign popcount21_sqs3_core_079 = ~(input_a[4] | input_a[4]);
  assign popcount21_sqs3_core_083 = ~input_a[14];
  assign popcount21_sqs3_core_085 = input_a[0] ^ input_a[18];
  assign popcount21_sqs3_core_087 = ~(input_a[0] & input_a[9]);
  assign popcount21_sqs3_core_090 = ~(input_a[11] & input_a[7]);
  assign popcount21_sqs3_core_091 = ~input_a[16];
  assign popcount21_sqs3_core_092 = input_a[11] & input_a[9];
  assign popcount21_sqs3_core_094 = input_a[16] ^ input_a[5];
  assign popcount21_sqs3_core_095 = ~(input_a[17] & input_a[18]);
  assign popcount21_sqs3_core_096 = ~(input_a[5] ^ input_a[18]);
  assign popcount21_sqs3_core_097 = ~(input_a[3] & input_a[8]);
  assign popcount21_sqs3_core_100 = ~(input_a[6] | input_a[18]);
  assign popcount21_sqs3_core_101 = ~(input_a[16] | input_a[11]);
  assign popcount21_sqs3_core_102 = ~(input_a[5] & input_a[17]);
  assign popcount21_sqs3_core_104 = ~(input_a[17] | input_a[13]);
  assign popcount21_sqs3_core_105 = input_a[6] ^ input_a[11];
  assign popcount21_sqs3_core_107 = input_a[20] ^ input_a[18];
  assign popcount21_sqs3_core_109 = input_a[4] & input_a[14];
  assign popcount21_sqs3_core_113 = ~(input_a[2] | input_a[0]);
  assign popcount21_sqs3_core_116 = ~input_a[6];
  assign popcount21_sqs3_core_117 = ~(input_a[20] & input_a[12]);
  assign popcount21_sqs3_core_118 = ~(input_a[16] | input_a[18]);
  assign popcount21_sqs3_core_120 = input_a[11] | input_a[19];
  assign popcount21_sqs3_core_121 = ~(input_a[15] ^ input_a[3]);
  assign popcount21_sqs3_core_123 = input_a[17] ^ input_a[11];
  assign popcount21_sqs3_core_124 = input_a[19] ^ input_a[10];
  assign popcount21_sqs3_core_125 = input_a[18] ^ input_a[3];
  assign popcount21_sqs3_core_127 = ~input_a[5];
  assign popcount21_sqs3_core_129 = ~input_a[7];
  assign popcount21_sqs3_core_130 = ~input_a[17];
  assign popcount21_sqs3_core_134 = input_a[3] | input_a[9];
  assign popcount21_sqs3_core_136 = ~(input_a[17] | input_a[4]);
  assign popcount21_sqs3_core_137 = ~input_a[9];
  assign popcount21_sqs3_core_138 = input_a[17] | input_a[4];
  assign popcount21_sqs3_core_140 = ~input_a[15];
  assign popcount21_sqs3_core_141 = ~input_a[7];
  assign popcount21_sqs3_core_142 = input_a[18] | input_a[0];
  assign popcount21_sqs3_core_144 = ~input_a[9];
  assign popcount21_sqs3_core_146 = input_a[13] | input_a[5];
  assign popcount21_sqs3_core_148 = input_a[18] ^ input_a[13];
  assign popcount21_sqs3_core_149 = ~(input_a[13] ^ input_a[12]);
  assign popcount21_sqs3_core_150 = input_a[16] ^ input_a[8];
  assign popcount21_sqs3_core_151 = ~(input_a[5] | input_a[2]);
  assign popcount21_sqs3_core_152 = input_a[16] | input_a[5];
  assign popcount21_sqs3_core_153 = ~(input_a[7] | input_a[9]);

  assign popcount21_sqs3_out[0] = input_a[17];
  assign popcount21_sqs3_out[1] = 1'b1;
  assign popcount21_sqs3_out[2] = 1'b0;
  assign popcount21_sqs3_out[3] = 1'b1;
  assign popcount21_sqs3_out[4] = 1'b0;
endmodule