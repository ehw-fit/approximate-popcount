// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.56721
// WCE=20.0
// EP=0.918543%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_sgw3(input [31:0] input_a, output [5:0] popcount32_sgw3_out);
  wire popcount32_sgw3_core_036;
  wire popcount32_sgw3_core_037;
  wire popcount32_sgw3_core_040;
  wire popcount32_sgw3_core_041;
  wire popcount32_sgw3_core_043;
  wire popcount32_sgw3_core_044;
  wire popcount32_sgw3_core_045;
  wire popcount32_sgw3_core_046;
  wire popcount32_sgw3_core_051;
  wire popcount32_sgw3_core_054;
  wire popcount32_sgw3_core_055;
  wire popcount32_sgw3_core_056;
  wire popcount32_sgw3_core_057;
  wire popcount32_sgw3_core_058;
  wire popcount32_sgw3_core_059;
  wire popcount32_sgw3_core_061;
  wire popcount32_sgw3_core_062;
  wire popcount32_sgw3_core_063;
  wire popcount32_sgw3_core_065;
  wire popcount32_sgw3_core_066_not;
  wire popcount32_sgw3_core_068;
  wire popcount32_sgw3_core_070;
  wire popcount32_sgw3_core_072;
  wire popcount32_sgw3_core_076;
  wire popcount32_sgw3_core_077;
  wire popcount32_sgw3_core_078;
  wire popcount32_sgw3_core_079;
  wire popcount32_sgw3_core_081;
  wire popcount32_sgw3_core_082;
  wire popcount32_sgw3_core_083;
  wire popcount32_sgw3_core_084;
  wire popcount32_sgw3_core_085;
  wire popcount32_sgw3_core_086;
  wire popcount32_sgw3_core_087;
  wire popcount32_sgw3_core_088;
  wire popcount32_sgw3_core_089;
  wire popcount32_sgw3_core_091;
  wire popcount32_sgw3_core_092;
  wire popcount32_sgw3_core_093;
  wire popcount32_sgw3_core_094;
  wire popcount32_sgw3_core_095;
  wire popcount32_sgw3_core_100;
  wire popcount32_sgw3_core_102;
  wire popcount32_sgw3_core_103;
  wire popcount32_sgw3_core_104;
  wire popcount32_sgw3_core_105;
  wire popcount32_sgw3_core_106;
  wire popcount32_sgw3_core_107;
  wire popcount32_sgw3_core_109;
  wire popcount32_sgw3_core_110;
  wire popcount32_sgw3_core_112;
  wire popcount32_sgw3_core_113;
  wire popcount32_sgw3_core_120;
  wire popcount32_sgw3_core_121;
  wire popcount32_sgw3_core_122;
  wire popcount32_sgw3_core_123;
  wire popcount32_sgw3_core_124;
  wire popcount32_sgw3_core_125;
  wire popcount32_sgw3_core_127_not;
  wire popcount32_sgw3_core_128;
  wire popcount32_sgw3_core_129;
  wire popcount32_sgw3_core_132;
  wire popcount32_sgw3_core_134;
  wire popcount32_sgw3_core_137;
  wire popcount32_sgw3_core_138;
  wire popcount32_sgw3_core_139;
  wire popcount32_sgw3_core_140;
  wire popcount32_sgw3_core_143;
  wire popcount32_sgw3_core_145;
  wire popcount32_sgw3_core_148;
  wire popcount32_sgw3_core_149;
  wire popcount32_sgw3_core_150;
  wire popcount32_sgw3_core_151;
  wire popcount32_sgw3_core_153;
  wire popcount32_sgw3_core_154_not;
  wire popcount32_sgw3_core_155;
  wire popcount32_sgw3_core_156;
  wire popcount32_sgw3_core_157;
  wire popcount32_sgw3_core_158;
  wire popcount32_sgw3_core_161;
  wire popcount32_sgw3_core_162;
  wire popcount32_sgw3_core_163;
  wire popcount32_sgw3_core_164;
  wire popcount32_sgw3_core_166;
  wire popcount32_sgw3_core_167;
  wire popcount32_sgw3_core_168;
  wire popcount32_sgw3_core_169;
  wire popcount32_sgw3_core_170;
  wire popcount32_sgw3_core_174;
  wire popcount32_sgw3_core_175;
  wire popcount32_sgw3_core_176;
  wire popcount32_sgw3_core_181;
  wire popcount32_sgw3_core_182;
  wire popcount32_sgw3_core_184;
  wire popcount32_sgw3_core_186;
  wire popcount32_sgw3_core_187;
  wire popcount32_sgw3_core_188;
  wire popcount32_sgw3_core_189;
  wire popcount32_sgw3_core_190;
  wire popcount32_sgw3_core_191;
  wire popcount32_sgw3_core_192;
  wire popcount32_sgw3_core_193;
  wire popcount32_sgw3_core_194;
  wire popcount32_sgw3_core_195;
  wire popcount32_sgw3_core_197;
  wire popcount32_sgw3_core_198;
  wire popcount32_sgw3_core_199;
  wire popcount32_sgw3_core_200;
  wire popcount32_sgw3_core_203;
  wire popcount32_sgw3_core_204;
  wire popcount32_sgw3_core_206;
  wire popcount32_sgw3_core_208;
  wire popcount32_sgw3_core_209;
  wire popcount32_sgw3_core_210;
  wire popcount32_sgw3_core_213;
  wire popcount32_sgw3_core_214;
  wire popcount32_sgw3_core_215;
  wire popcount32_sgw3_core_216;
  wire popcount32_sgw3_core_217;
  wire popcount32_sgw3_core_219;
  wire popcount32_sgw3_core_222;
  wire popcount32_sgw3_core_223;
  wire popcount32_sgw3_core_224;
  wire popcount32_sgw3_core_225;

  assign popcount32_sgw3_core_036 = ~(input_a[0] ^ input_a[12]);
  assign popcount32_sgw3_core_037 = input_a[25] | input_a[20];
  assign popcount32_sgw3_core_040 = ~(input_a[17] | input_a[21]);
  assign popcount32_sgw3_core_041 = ~(input_a[28] ^ input_a[9]);
  assign popcount32_sgw3_core_043 = ~(input_a[19] | input_a[26]);
  assign popcount32_sgw3_core_044 = ~input_a[28];
  assign popcount32_sgw3_core_045 = ~(input_a[19] & input_a[18]);
  assign popcount32_sgw3_core_046 = input_a[29] | input_a[23];
  assign popcount32_sgw3_core_051 = input_a[26] ^ input_a[13];
  assign popcount32_sgw3_core_054 = input_a[1] | input_a[14];
  assign popcount32_sgw3_core_055 = ~input_a[12];
  assign popcount32_sgw3_core_056 = ~(input_a[13] ^ input_a[4]);
  assign popcount32_sgw3_core_057 = ~(input_a[9] & input_a[13]);
  assign popcount32_sgw3_core_058 = ~input_a[18];
  assign popcount32_sgw3_core_059 = ~(input_a[17] & input_a[27]);
  assign popcount32_sgw3_core_061 = input_a[0] ^ input_a[25];
  assign popcount32_sgw3_core_062 = ~input_a[3];
  assign popcount32_sgw3_core_063 = input_a[29] ^ input_a[0];
  assign popcount32_sgw3_core_065 = input_a[26] | input_a[19];
  assign popcount32_sgw3_core_066_not = ~input_a[22];
  assign popcount32_sgw3_core_068 = ~(input_a[6] | input_a[10]);
  assign popcount32_sgw3_core_070 = input_a[30] & input_a[2];
  assign popcount32_sgw3_core_072 = ~(input_a[24] ^ input_a[26]);
  assign popcount32_sgw3_core_076 = input_a[4] ^ input_a[31];
  assign popcount32_sgw3_core_077 = input_a[30] ^ input_a[17];
  assign popcount32_sgw3_core_078 = ~(input_a[13] & input_a[18]);
  assign popcount32_sgw3_core_079 = ~(input_a[16] & input_a[27]);
  assign popcount32_sgw3_core_081 = input_a[1] ^ input_a[11];
  assign popcount32_sgw3_core_082 = ~(input_a[28] & input_a[17]);
  assign popcount32_sgw3_core_083 = input_a[19] ^ input_a[25];
  assign popcount32_sgw3_core_084 = ~(input_a[14] & input_a[18]);
  assign popcount32_sgw3_core_085 = ~input_a[27];
  assign popcount32_sgw3_core_086 = ~(input_a[1] | input_a[26]);
  assign popcount32_sgw3_core_087 = ~input_a[10];
  assign popcount32_sgw3_core_088 = input_a[23] & input_a[13];
  assign popcount32_sgw3_core_089 = input_a[11] | input_a[13];
  assign popcount32_sgw3_core_091 = ~(input_a[8] & input_a[21]);
  assign popcount32_sgw3_core_092 = ~(input_a[14] & input_a[12]);
  assign popcount32_sgw3_core_093 = ~input_a[28];
  assign popcount32_sgw3_core_094 = input_a[12] ^ input_a[1];
  assign popcount32_sgw3_core_095 = ~(input_a[15] ^ input_a[14]);
  assign popcount32_sgw3_core_100 = ~(input_a[25] | input_a[1]);
  assign popcount32_sgw3_core_102 = input_a[26] | input_a[23];
  assign popcount32_sgw3_core_103 = ~input_a[27];
  assign popcount32_sgw3_core_104 = ~(input_a[4] & input_a[30]);
  assign popcount32_sgw3_core_105 = ~(input_a[30] ^ input_a[1]);
  assign popcount32_sgw3_core_106 = input_a[30] & input_a[27];
  assign popcount32_sgw3_core_107 = ~input_a[13];
  assign popcount32_sgw3_core_109 = input_a[17] & input_a[27];
  assign popcount32_sgw3_core_110 = input_a[23] | input_a[31];
  assign popcount32_sgw3_core_112 = ~(input_a[16] & input_a[12]);
  assign popcount32_sgw3_core_113 = ~(input_a[12] | input_a[16]);
  assign popcount32_sgw3_core_120 = ~(input_a[2] ^ input_a[18]);
  assign popcount32_sgw3_core_121 = ~(input_a[25] | input_a[18]);
  assign popcount32_sgw3_core_122 = input_a[11] ^ input_a[15];
  assign popcount32_sgw3_core_123 = ~(input_a[30] | input_a[18]);
  assign popcount32_sgw3_core_124 = ~input_a[18];
  assign popcount32_sgw3_core_125 = ~input_a[11];
  assign popcount32_sgw3_core_127_not = ~input_a[5];
  assign popcount32_sgw3_core_128 = input_a[21] | input_a[24];
  assign popcount32_sgw3_core_129 = ~input_a[25];
  assign popcount32_sgw3_core_132 = ~input_a[20];
  assign popcount32_sgw3_core_134 = input_a[23] ^ input_a[18];
  assign popcount32_sgw3_core_137 = ~(input_a[18] | input_a[24]);
  assign popcount32_sgw3_core_138 = ~input_a[25];
  assign popcount32_sgw3_core_139 = input_a[1] & input_a[25];
  assign popcount32_sgw3_core_140 = ~(input_a[1] ^ input_a[28]);
  assign popcount32_sgw3_core_143 = ~input_a[18];
  assign popcount32_sgw3_core_145 = ~(input_a[3] | input_a[24]);
  assign popcount32_sgw3_core_148 = input_a[26] & input_a[15];
  assign popcount32_sgw3_core_149 = input_a[7] ^ input_a[11];
  assign popcount32_sgw3_core_150 = ~input_a[23];
  assign popcount32_sgw3_core_151 = input_a[22] | input_a[10];
  assign popcount32_sgw3_core_153 = ~input_a[11];
  assign popcount32_sgw3_core_154_not = ~input_a[3];
  assign popcount32_sgw3_core_155 = input_a[1] ^ input_a[21];
  assign popcount32_sgw3_core_156 = input_a[18] & input_a[27];
  assign popcount32_sgw3_core_157 = ~(input_a[2] | input_a[14]);
  assign popcount32_sgw3_core_158 = input_a[2] | input_a[8];
  assign popcount32_sgw3_core_161 = ~input_a[16];
  assign popcount32_sgw3_core_162 = input_a[3] & input_a[25];
  assign popcount32_sgw3_core_163 = input_a[16] ^ input_a[31];
  assign popcount32_sgw3_core_164 = input_a[31] | input_a[7];
  assign popcount32_sgw3_core_166 = ~(input_a[18] & input_a[29]);
  assign popcount32_sgw3_core_167 = input_a[2] & input_a[14];
  assign popcount32_sgw3_core_168 = ~(input_a[24] | input_a[5]);
  assign popcount32_sgw3_core_169 = input_a[11] ^ input_a[30];
  assign popcount32_sgw3_core_170 = ~(input_a[19] & input_a[24]);
  assign popcount32_sgw3_core_174 = input_a[13] | input_a[17];
  assign popcount32_sgw3_core_175 = ~(input_a[31] | input_a[8]);
  assign popcount32_sgw3_core_176 = input_a[31] ^ input_a[14];
  assign popcount32_sgw3_core_181 = input_a[21] & input_a[10];
  assign popcount32_sgw3_core_182 = input_a[23] & input_a[23];
  assign popcount32_sgw3_core_184 = input_a[13] ^ input_a[2];
  assign popcount32_sgw3_core_186 = ~(input_a[5] ^ input_a[1]);
  assign popcount32_sgw3_core_187 = ~(input_a[25] & input_a[27]);
  assign popcount32_sgw3_core_188 = input_a[0] ^ input_a[22];
  assign popcount32_sgw3_core_189 = ~(input_a[13] | input_a[28]);
  assign popcount32_sgw3_core_190 = ~(input_a[2] & input_a[30]);
  assign popcount32_sgw3_core_191 = input_a[9] | input_a[22];
  assign popcount32_sgw3_core_192 = input_a[16] ^ input_a[18];
  assign popcount32_sgw3_core_193 = ~(input_a[22] ^ input_a[28]);
  assign popcount32_sgw3_core_194 = ~(input_a[19] | input_a[29]);
  assign popcount32_sgw3_core_195 = ~(input_a[1] & input_a[6]);
  assign popcount32_sgw3_core_197 = input_a[25] ^ input_a[8];
  assign popcount32_sgw3_core_198 = ~(input_a[15] & input_a[31]);
  assign popcount32_sgw3_core_199 = ~(input_a[8] & input_a[7]);
  assign popcount32_sgw3_core_200 = ~(input_a[19] | input_a[26]);
  assign popcount32_sgw3_core_203 = ~(input_a[27] | input_a[29]);
  assign popcount32_sgw3_core_204 = input_a[3] & input_a[23];
  assign popcount32_sgw3_core_206 = ~(input_a[28] ^ input_a[2]);
  assign popcount32_sgw3_core_208 = input_a[19] | input_a[23];
  assign popcount32_sgw3_core_209 = ~(input_a[15] | input_a[12]);
  assign popcount32_sgw3_core_210 = input_a[15] | input_a[12];
  assign popcount32_sgw3_core_213 = ~input_a[6];
  assign popcount32_sgw3_core_214 = ~(input_a[0] & input_a[22]);
  assign popcount32_sgw3_core_215 = ~input_a[31];
  assign popcount32_sgw3_core_216 = input_a[13] ^ input_a[30];
  assign popcount32_sgw3_core_217 = ~(input_a[30] & input_a[7]);
  assign popcount32_sgw3_core_219 = input_a[24] ^ input_a[7];
  assign popcount32_sgw3_core_222 = input_a[23] | input_a[1];
  assign popcount32_sgw3_core_223 = ~input_a[20];
  assign popcount32_sgw3_core_224 = ~(input_a[10] | input_a[24]);
  assign popcount32_sgw3_core_225 = ~(input_a[10] | input_a[28]);

  assign popcount32_sgw3_out[0] = 1'b0;
  assign popcount32_sgw3_out[1] = input_a[21];
  assign popcount32_sgw3_out[2] = input_a[2];
  assign popcount32_sgw3_out[3] = 1'b0;
  assign popcount32_sgw3_out[4] = 1'b1;
  assign popcount32_sgw3_out[5] = 1'b0;
endmodule