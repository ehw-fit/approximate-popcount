// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.2392
// WCE=16.0
// EP=0.86005%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_j5tm(input [30:0] input_a, output [4:0] popcount31_j5tm_out);
  wire popcount31_j5tm_core_033;
  wire popcount31_j5tm_core_035;
  wire popcount31_j5tm_core_036;
  wire popcount31_j5tm_core_037;
  wire popcount31_j5tm_core_038;
  wire popcount31_j5tm_core_039;
  wire popcount31_j5tm_core_042;
  wire popcount31_j5tm_core_043;
  wire popcount31_j5tm_core_045;
  wire popcount31_j5tm_core_046;
  wire popcount31_j5tm_core_049;
  wire popcount31_j5tm_core_051;
  wire popcount31_j5tm_core_052;
  wire popcount31_j5tm_core_053;
  wire popcount31_j5tm_core_055_not;
  wire popcount31_j5tm_core_056;
  wire popcount31_j5tm_core_059;
  wire popcount31_j5tm_core_061;
  wire popcount31_j5tm_core_062;
  wire popcount31_j5tm_core_064;
  wire popcount31_j5tm_core_065;
  wire popcount31_j5tm_core_067;
  wire popcount31_j5tm_core_070;
  wire popcount31_j5tm_core_071;
  wire popcount31_j5tm_core_073;
  wire popcount31_j5tm_core_075;
  wire popcount31_j5tm_core_076;
  wire popcount31_j5tm_core_077;
  wire popcount31_j5tm_core_078;
  wire popcount31_j5tm_core_080;
  wire popcount31_j5tm_core_082;
  wire popcount31_j5tm_core_084;
  wire popcount31_j5tm_core_087;
  wire popcount31_j5tm_core_089;
  wire popcount31_j5tm_core_090;
  wire popcount31_j5tm_core_092;
  wire popcount31_j5tm_core_094;
  wire popcount31_j5tm_core_100;
  wire popcount31_j5tm_core_104;
  wire popcount31_j5tm_core_105;
  wire popcount31_j5tm_core_106;
  wire popcount31_j5tm_core_110;
  wire popcount31_j5tm_core_113;
  wire popcount31_j5tm_core_114;
  wire popcount31_j5tm_core_115;
  wire popcount31_j5tm_core_119;
  wire popcount31_j5tm_core_121;
  wire popcount31_j5tm_core_123;
  wire popcount31_j5tm_core_124;
  wire popcount31_j5tm_core_125;
  wire popcount31_j5tm_core_126;
  wire popcount31_j5tm_core_130;
  wire popcount31_j5tm_core_131;
  wire popcount31_j5tm_core_133;
  wire popcount31_j5tm_core_134;
  wire popcount31_j5tm_core_136;
  wire popcount31_j5tm_core_138;
  wire popcount31_j5tm_core_140;
  wire popcount31_j5tm_core_141;
  wire popcount31_j5tm_core_143;
  wire popcount31_j5tm_core_145;
  wire popcount31_j5tm_core_147;
  wire popcount31_j5tm_core_149;
  wire popcount31_j5tm_core_151;
  wire popcount31_j5tm_core_152;
  wire popcount31_j5tm_core_154;
  wire popcount31_j5tm_core_155;
  wire popcount31_j5tm_core_156;
  wire popcount31_j5tm_core_157;
  wire popcount31_j5tm_core_158;
  wire popcount31_j5tm_core_159;
  wire popcount31_j5tm_core_161;
  wire popcount31_j5tm_core_163;
  wire popcount31_j5tm_core_165;
  wire popcount31_j5tm_core_171;
  wire popcount31_j5tm_core_173;
  wire popcount31_j5tm_core_174;
  wire popcount31_j5tm_core_175;
  wire popcount31_j5tm_core_176;
  wire popcount31_j5tm_core_177;
  wire popcount31_j5tm_core_178;
  wire popcount31_j5tm_core_179;
  wire popcount31_j5tm_core_182;
  wire popcount31_j5tm_core_184;
  wire popcount31_j5tm_core_186;
  wire popcount31_j5tm_core_187;
  wire popcount31_j5tm_core_188;
  wire popcount31_j5tm_core_189;
  wire popcount31_j5tm_core_190;
  wire popcount31_j5tm_core_191;
  wire popcount31_j5tm_core_192;
  wire popcount31_j5tm_core_194;
  wire popcount31_j5tm_core_195;
  wire popcount31_j5tm_core_197;
  wire popcount31_j5tm_core_199;
  wire popcount31_j5tm_core_200;
  wire popcount31_j5tm_core_202;
  wire popcount31_j5tm_core_205;
  wire popcount31_j5tm_core_206;
  wire popcount31_j5tm_core_208;
  wire popcount31_j5tm_core_209;
  wire popcount31_j5tm_core_211;
  wire popcount31_j5tm_core_213;
  wire popcount31_j5tm_core_214;
  wire popcount31_j5tm_core_215;
  wire popcount31_j5tm_core_216;

  assign popcount31_j5tm_core_033 = ~(input_a[15] & input_a[26]);
  assign popcount31_j5tm_core_035 = input_a[14] ^ input_a[21];
  assign popcount31_j5tm_core_036 = ~input_a[15];
  assign popcount31_j5tm_core_037 = input_a[10] ^ input_a[2];
  assign popcount31_j5tm_core_038 = input_a[16] ^ input_a[17];
  assign popcount31_j5tm_core_039 = input_a[23] ^ input_a[24];
  assign popcount31_j5tm_core_042 = ~(input_a[11] ^ input_a[14]);
  assign popcount31_j5tm_core_043 = ~(input_a[4] & input_a[18]);
  assign popcount31_j5tm_core_045 = ~(input_a[23] | input_a[1]);
  assign popcount31_j5tm_core_046 = input_a[25] ^ input_a[8];
  assign popcount31_j5tm_core_049 = ~input_a[14];
  assign popcount31_j5tm_core_051 = input_a[29] & input_a[30];
  assign popcount31_j5tm_core_052 = input_a[7] ^ input_a[26];
  assign popcount31_j5tm_core_053 = input_a[20] ^ input_a[22];
  assign popcount31_j5tm_core_055_not = ~input_a[5];
  assign popcount31_j5tm_core_056 = ~(input_a[22] | input_a[19]);
  assign popcount31_j5tm_core_059 = ~input_a[0];
  assign popcount31_j5tm_core_061 = input_a[8] | input_a[17];
  assign popcount31_j5tm_core_062 = input_a[29] | input_a[6];
  assign popcount31_j5tm_core_064 = input_a[29] & input_a[20];
  assign popcount31_j5tm_core_065 = ~(input_a[15] ^ input_a[11]);
  assign popcount31_j5tm_core_067 = input_a[8] & input_a[29];
  assign popcount31_j5tm_core_070 = input_a[13] | input_a[9];
  assign popcount31_j5tm_core_071 = input_a[16] | input_a[0];
  assign popcount31_j5tm_core_073 = ~(input_a[30] ^ input_a[15]);
  assign popcount31_j5tm_core_075 = ~(input_a[5] ^ input_a[17]);
  assign popcount31_j5tm_core_076 = ~(input_a[18] & input_a[4]);
  assign popcount31_j5tm_core_077 = input_a[23] | input_a[18];
  assign popcount31_j5tm_core_078 = input_a[25] ^ input_a[16];
  assign popcount31_j5tm_core_080 = ~input_a[16];
  assign popcount31_j5tm_core_082 = input_a[10] | input_a[4];
  assign popcount31_j5tm_core_084 = input_a[10] & input_a[24];
  assign popcount31_j5tm_core_087 = input_a[28] | input_a[28];
  assign popcount31_j5tm_core_089 = ~(input_a[7] ^ input_a[23]);
  assign popcount31_j5tm_core_090 = ~(input_a[12] ^ input_a[0]);
  assign popcount31_j5tm_core_092 = input_a[27] & input_a[17];
  assign popcount31_j5tm_core_094 = input_a[4] ^ input_a[14];
  assign popcount31_j5tm_core_100 = ~(input_a[7] | input_a[2]);
  assign popcount31_j5tm_core_104 = ~(input_a[16] ^ input_a[6]);
  assign popcount31_j5tm_core_105 = input_a[16] | input_a[15];
  assign popcount31_j5tm_core_106 = ~(input_a[24] ^ input_a[25]);
  assign popcount31_j5tm_core_110 = input_a[11] ^ input_a[7];
  assign popcount31_j5tm_core_113 = ~(input_a[18] | input_a[15]);
  assign popcount31_j5tm_core_114 = ~(input_a[2] | input_a[24]);
  assign popcount31_j5tm_core_115 = input_a[19] & input_a[24];
  assign popcount31_j5tm_core_119 = ~input_a[15];
  assign popcount31_j5tm_core_121 = input_a[9] & input_a[20];
  assign popcount31_j5tm_core_123 = ~input_a[1];
  assign popcount31_j5tm_core_124 = input_a[2] ^ input_a[4];
  assign popcount31_j5tm_core_125 = ~(input_a[23] ^ input_a[5]);
  assign popcount31_j5tm_core_126 = input_a[10] & input_a[17];
  assign popcount31_j5tm_core_130 = ~(input_a[7] ^ input_a[24]);
  assign popcount31_j5tm_core_131 = ~(input_a[6] ^ input_a[20]);
  assign popcount31_j5tm_core_133 = ~input_a[23];
  assign popcount31_j5tm_core_134 = input_a[19] | input_a[11];
  assign popcount31_j5tm_core_136 = input_a[10] & input_a[20];
  assign popcount31_j5tm_core_138 = ~(input_a[1] | input_a[29]);
  assign popcount31_j5tm_core_140 = ~(input_a[6] | input_a[29]);
  assign popcount31_j5tm_core_141 = input_a[13] & input_a[23];
  assign popcount31_j5tm_core_143 = ~(input_a[27] | input_a[11]);
  assign popcount31_j5tm_core_145 = input_a[12] & input_a[17];
  assign popcount31_j5tm_core_147 = input_a[20] & input_a[14];
  assign popcount31_j5tm_core_149 = input_a[26] ^ input_a[21];
  assign popcount31_j5tm_core_151 = ~(input_a[23] ^ input_a[5]);
  assign popcount31_j5tm_core_152 = ~(input_a[5] & input_a[8]);
  assign popcount31_j5tm_core_154 = ~(input_a[7] & input_a[0]);
  assign popcount31_j5tm_core_155 = ~(input_a[17] & input_a[7]);
  assign popcount31_j5tm_core_156 = input_a[6] ^ input_a[23];
  assign popcount31_j5tm_core_157 = ~(input_a[17] & input_a[2]);
  assign popcount31_j5tm_core_158 = ~(input_a[17] | input_a[9]);
  assign popcount31_j5tm_core_159 = ~input_a[9];
  assign popcount31_j5tm_core_161 = input_a[18] ^ input_a[3];
  assign popcount31_j5tm_core_163 = ~(input_a[10] ^ input_a[17]);
  assign popcount31_j5tm_core_165 = ~(input_a[5] ^ input_a[8]);
  assign popcount31_j5tm_core_171 = input_a[18] | input_a[10];
  assign popcount31_j5tm_core_173 = ~(input_a[24] & input_a[16]);
  assign popcount31_j5tm_core_174 = input_a[5] & input_a[16];
  assign popcount31_j5tm_core_175 = input_a[23] ^ input_a[11];
  assign popcount31_j5tm_core_176 = ~input_a[7];
  assign popcount31_j5tm_core_177 = ~(input_a[23] & input_a[3]);
  assign popcount31_j5tm_core_178 = ~(input_a[16] ^ input_a[10]);
  assign popcount31_j5tm_core_179 = ~(input_a[2] & input_a[6]);
  assign popcount31_j5tm_core_182 = ~input_a[18];
  assign popcount31_j5tm_core_184 = input_a[28] & input_a[16];
  assign popcount31_j5tm_core_186 = ~input_a[29];
  assign popcount31_j5tm_core_187 = ~(input_a[13] ^ input_a[29]);
  assign popcount31_j5tm_core_188 = ~(input_a[6] | input_a[18]);
  assign popcount31_j5tm_core_189 = ~(input_a[27] | input_a[28]);
  assign popcount31_j5tm_core_190 = ~(input_a[4] ^ input_a[13]);
  assign popcount31_j5tm_core_191 = ~(input_a[9] | input_a[30]);
  assign popcount31_j5tm_core_192 = input_a[23] ^ input_a[5];
  assign popcount31_j5tm_core_194 = input_a[27] | input_a[21];
  assign popcount31_j5tm_core_195 = input_a[12] ^ input_a[0];
  assign popcount31_j5tm_core_197 = input_a[13] | input_a[6];
  assign popcount31_j5tm_core_199 = input_a[24] | input_a[28];
  assign popcount31_j5tm_core_200 = input_a[30] | input_a[11];
  assign popcount31_j5tm_core_202 = input_a[23] ^ input_a[19];
  assign popcount31_j5tm_core_205 = ~(input_a[11] & input_a[22]);
  assign popcount31_j5tm_core_206 = ~(input_a[5] ^ input_a[23]);
  assign popcount31_j5tm_core_208 = input_a[0] & input_a[14];
  assign popcount31_j5tm_core_209 = ~input_a[4];
  assign popcount31_j5tm_core_211 = input_a[2] ^ input_a[5];
  assign popcount31_j5tm_core_213 = ~(input_a[2] ^ input_a[26]);
  assign popcount31_j5tm_core_214 = ~(input_a[2] ^ input_a[1]);
  assign popcount31_j5tm_core_215 = ~(input_a[29] ^ input_a[2]);
  assign popcount31_j5tm_core_216 = input_a[30] & input_a[17];

  assign popcount31_j5tm_out[0] = 1'b1;
  assign popcount31_j5tm_out[1] = 1'b1;
  assign popcount31_j5tm_out[2] = 1'b1;
  assign popcount31_j5tm_out[3] = 1'b1;
  assign popcount31_j5tm_out[4] = 1'b0;
endmodule