// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.64747
// WCE=27.0
// EP=0.970683%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount31_1hjn(input [30:0] input_a, output [4:0] popcount31_1hjn_out);
  wire popcount31_1hjn_core_035;
  wire popcount31_1hjn_core_037;
  wire popcount31_1hjn_core_038;
  wire popcount31_1hjn_core_039;
  wire popcount31_1hjn_core_040;
  wire popcount31_1hjn_core_041;
  wire popcount31_1hjn_core_042;
  wire popcount31_1hjn_core_043;
  wire popcount31_1hjn_core_044;
  wire popcount31_1hjn_core_047;
  wire popcount31_1hjn_core_050;
  wire popcount31_1hjn_core_051;
  wire popcount31_1hjn_core_052;
  wire popcount31_1hjn_core_053;
  wire popcount31_1hjn_core_055;
  wire popcount31_1hjn_core_056;
  wire popcount31_1hjn_core_057;
  wire popcount31_1hjn_core_058;
  wire popcount31_1hjn_core_060;
  wire popcount31_1hjn_core_061;
  wire popcount31_1hjn_core_062;
  wire popcount31_1hjn_core_064;
  wire popcount31_1hjn_core_065;
  wire popcount31_1hjn_core_066;
  wire popcount31_1hjn_core_067;
  wire popcount31_1hjn_core_068;
  wire popcount31_1hjn_core_071;
  wire popcount31_1hjn_core_072;
  wire popcount31_1hjn_core_073;
  wire popcount31_1hjn_core_074;
  wire popcount31_1hjn_core_075;
  wire popcount31_1hjn_core_076;
  wire popcount31_1hjn_core_079;
  wire popcount31_1hjn_core_080;
  wire popcount31_1hjn_core_082_not;
  wire popcount31_1hjn_core_083;
  wire popcount31_1hjn_core_084;
  wire popcount31_1hjn_core_085;
  wire popcount31_1hjn_core_088;
  wire popcount31_1hjn_core_092;
  wire popcount31_1hjn_core_093;
  wire popcount31_1hjn_core_094;
  wire popcount31_1hjn_core_095;
  wire popcount31_1hjn_core_097;
  wire popcount31_1hjn_core_099;
  wire popcount31_1hjn_core_100;
  wire popcount31_1hjn_core_103;
  wire popcount31_1hjn_core_104;
  wire popcount31_1hjn_core_106;
  wire popcount31_1hjn_core_108;
  wire popcount31_1hjn_core_110;
  wire popcount31_1hjn_core_111;
  wire popcount31_1hjn_core_113;
  wire popcount31_1hjn_core_117;
  wire popcount31_1hjn_core_119;
  wire popcount31_1hjn_core_121;
  wire popcount31_1hjn_core_122;
  wire popcount31_1hjn_core_123;
  wire popcount31_1hjn_core_124;
  wire popcount31_1hjn_core_125_not;
  wire popcount31_1hjn_core_126;
  wire popcount31_1hjn_core_130;
  wire popcount31_1hjn_core_132;
  wire popcount31_1hjn_core_135_not;
  wire popcount31_1hjn_core_139;
  wire popcount31_1hjn_core_140;
  wire popcount31_1hjn_core_143;
  wire popcount31_1hjn_core_145;
  wire popcount31_1hjn_core_146;
  wire popcount31_1hjn_core_147;
  wire popcount31_1hjn_core_148;
  wire popcount31_1hjn_core_149;
  wire popcount31_1hjn_core_150_not;
  wire popcount31_1hjn_core_151;
  wire popcount31_1hjn_core_152;
  wire popcount31_1hjn_core_154;
  wire popcount31_1hjn_core_155;
  wire popcount31_1hjn_core_156;
  wire popcount31_1hjn_core_158;
  wire popcount31_1hjn_core_160;
  wire popcount31_1hjn_core_162;
  wire popcount31_1hjn_core_163;
  wire popcount31_1hjn_core_166;
  wire popcount31_1hjn_core_168;
  wire popcount31_1hjn_core_169;
  wire popcount31_1hjn_core_170;
  wire popcount31_1hjn_core_171;
  wire popcount31_1hjn_core_173;
  wire popcount31_1hjn_core_174;
  wire popcount31_1hjn_core_175;
  wire popcount31_1hjn_core_176;
  wire popcount31_1hjn_core_177;
  wire popcount31_1hjn_core_178;
  wire popcount31_1hjn_core_179;
  wire popcount31_1hjn_core_180;
  wire popcount31_1hjn_core_181;
  wire popcount31_1hjn_core_182;
  wire popcount31_1hjn_core_183;
  wire popcount31_1hjn_core_185;
  wire popcount31_1hjn_core_186;
  wire popcount31_1hjn_core_189;
  wire popcount31_1hjn_core_190;
  wire popcount31_1hjn_core_191;
  wire popcount31_1hjn_core_192;
  wire popcount31_1hjn_core_193;
  wire popcount31_1hjn_core_197;
  wire popcount31_1hjn_core_198;
  wire popcount31_1hjn_core_199;
  wire popcount31_1hjn_core_201;
  wire popcount31_1hjn_core_202;
  wire popcount31_1hjn_core_203;
  wire popcount31_1hjn_core_206;
  wire popcount31_1hjn_core_207;
  wire popcount31_1hjn_core_208;
  wire popcount31_1hjn_core_209;
  wire popcount31_1hjn_core_211;
  wire popcount31_1hjn_core_212;
  wire popcount31_1hjn_core_214;
  wire popcount31_1hjn_core_215;
  wire popcount31_1hjn_core_217;

  assign popcount31_1hjn_core_035 = ~input_a[10];
  assign popcount31_1hjn_core_037 = ~(input_a[28] | input_a[26]);
  assign popcount31_1hjn_core_038 = ~input_a[3];
  assign popcount31_1hjn_core_039 = ~(input_a[23] | input_a[11]);
  assign popcount31_1hjn_core_040 = input_a[18] ^ input_a[5];
  assign popcount31_1hjn_core_041 = input_a[26] ^ input_a[23];
  assign popcount31_1hjn_core_042 = ~(input_a[25] | input_a[25]);
  assign popcount31_1hjn_core_043 = ~(input_a[11] ^ input_a[21]);
  assign popcount31_1hjn_core_044 = ~(input_a[23] & input_a[0]);
  assign popcount31_1hjn_core_047 = input_a[21] ^ input_a[30];
  assign popcount31_1hjn_core_050 = ~input_a[0];
  assign popcount31_1hjn_core_051 = input_a[23] ^ input_a[30];
  assign popcount31_1hjn_core_052 = ~(input_a[8] ^ input_a[0]);
  assign popcount31_1hjn_core_053 = ~input_a[8];
  assign popcount31_1hjn_core_055 = ~(input_a[27] ^ input_a[17]);
  assign popcount31_1hjn_core_056 = input_a[8] ^ input_a[29];
  assign popcount31_1hjn_core_057 = ~input_a[11];
  assign popcount31_1hjn_core_058 = ~(input_a[28] ^ input_a[16]);
  assign popcount31_1hjn_core_060 = ~(input_a[6] & input_a[12]);
  assign popcount31_1hjn_core_061 = ~(input_a[8] ^ input_a[3]);
  assign popcount31_1hjn_core_062 = ~(input_a[1] ^ input_a[0]);
  assign popcount31_1hjn_core_064 = ~(input_a[13] & input_a[7]);
  assign popcount31_1hjn_core_065 = input_a[0] ^ input_a[15];
  assign popcount31_1hjn_core_066 = ~(input_a[0] & input_a[28]);
  assign popcount31_1hjn_core_067 = ~input_a[9];
  assign popcount31_1hjn_core_068 = ~input_a[29];
  assign popcount31_1hjn_core_071 = ~(input_a[1] | input_a[23]);
  assign popcount31_1hjn_core_072 = input_a[25] & input_a[13];
  assign popcount31_1hjn_core_073 = ~(input_a[14] | input_a[8]);
  assign popcount31_1hjn_core_074 = ~(input_a[22] | input_a[8]);
  assign popcount31_1hjn_core_075 = ~input_a[24];
  assign popcount31_1hjn_core_076 = ~(input_a[6] | input_a[11]);
  assign popcount31_1hjn_core_079 = input_a[29] | input_a[29];
  assign popcount31_1hjn_core_080 = input_a[9] ^ input_a[2];
  assign popcount31_1hjn_core_082_not = ~input_a[0];
  assign popcount31_1hjn_core_083 = input_a[21] & input_a[24];
  assign popcount31_1hjn_core_084 = input_a[20] | input_a[27];
  assign popcount31_1hjn_core_085 = ~input_a[2];
  assign popcount31_1hjn_core_088 = input_a[2] | input_a[15];
  assign popcount31_1hjn_core_092 = input_a[4] & input_a[19];
  assign popcount31_1hjn_core_093 = ~input_a[13];
  assign popcount31_1hjn_core_094 = ~(input_a[25] | input_a[14]);
  assign popcount31_1hjn_core_095 = ~input_a[1];
  assign popcount31_1hjn_core_097 = ~(input_a[24] & input_a[27]);
  assign popcount31_1hjn_core_099 = input_a[8] ^ input_a[14];
  assign popcount31_1hjn_core_100 = input_a[11] | input_a[18];
  assign popcount31_1hjn_core_103 = ~(input_a[13] ^ input_a[0]);
  assign popcount31_1hjn_core_104 = input_a[9] ^ input_a[10];
  assign popcount31_1hjn_core_106 = ~(input_a[3] & input_a[11]);
  assign popcount31_1hjn_core_108 = input_a[6] & input_a[7];
  assign popcount31_1hjn_core_110 = input_a[17] ^ input_a[9];
  assign popcount31_1hjn_core_111 = ~(input_a[12] | input_a[5]);
  assign popcount31_1hjn_core_113 = ~(input_a[1] ^ input_a[10]);
  assign popcount31_1hjn_core_117 = input_a[8] & input_a[11];
  assign popcount31_1hjn_core_119 = ~(input_a[11] & input_a[27]);
  assign popcount31_1hjn_core_121 = ~input_a[5];
  assign popcount31_1hjn_core_122 = input_a[1] | input_a[7];
  assign popcount31_1hjn_core_123 = ~(input_a[20] ^ input_a[20]);
  assign popcount31_1hjn_core_124 = input_a[15] ^ input_a[20];
  assign popcount31_1hjn_core_125_not = ~input_a[24];
  assign popcount31_1hjn_core_126 = ~(input_a[23] ^ input_a[0]);
  assign popcount31_1hjn_core_130 = input_a[8] | input_a[3];
  assign popcount31_1hjn_core_132 = ~(input_a[27] | input_a[6]);
  assign popcount31_1hjn_core_135_not = ~input_a[8];
  assign popcount31_1hjn_core_139 = ~(input_a[18] & input_a[21]);
  assign popcount31_1hjn_core_140 = input_a[21] | input_a[26];
  assign popcount31_1hjn_core_143 = input_a[10] ^ input_a[14];
  assign popcount31_1hjn_core_145 = input_a[16] & input_a[3];
  assign popcount31_1hjn_core_146 = input_a[5] ^ input_a[10];
  assign popcount31_1hjn_core_147 = ~input_a[14];
  assign popcount31_1hjn_core_148 = ~(input_a[25] ^ input_a[17]);
  assign popcount31_1hjn_core_149 = input_a[0] & input_a[22];
  assign popcount31_1hjn_core_150_not = ~input_a[12];
  assign popcount31_1hjn_core_151 = ~(input_a[1] & input_a[28]);
  assign popcount31_1hjn_core_152 = ~(input_a[21] & input_a[8]);
  assign popcount31_1hjn_core_154 = ~(input_a[24] | input_a[2]);
  assign popcount31_1hjn_core_155 = input_a[4] ^ input_a[30];
  assign popcount31_1hjn_core_156 = ~(input_a[20] | input_a[14]);
  assign popcount31_1hjn_core_158 = ~(input_a[5] & input_a[17]);
  assign popcount31_1hjn_core_160 = ~(input_a[6] | input_a[19]);
  assign popcount31_1hjn_core_162 = ~(input_a[20] | input_a[22]);
  assign popcount31_1hjn_core_163 = ~(input_a[28] ^ input_a[5]);
  assign popcount31_1hjn_core_166 = ~(input_a[22] | input_a[18]);
  assign popcount31_1hjn_core_168 = input_a[21] | input_a[0];
  assign popcount31_1hjn_core_169 = ~input_a[22];
  assign popcount31_1hjn_core_170 = input_a[25] & input_a[11];
  assign popcount31_1hjn_core_171 = input_a[30] & input_a[27];
  assign popcount31_1hjn_core_173 = input_a[9] ^ input_a[14];
  assign popcount31_1hjn_core_174 = input_a[22] ^ input_a[3];
  assign popcount31_1hjn_core_175 = ~input_a[30];
  assign popcount31_1hjn_core_176 = input_a[5] ^ input_a[15];
  assign popcount31_1hjn_core_177 = ~(input_a[24] & input_a[2]);
  assign popcount31_1hjn_core_178 = ~input_a[16];
  assign popcount31_1hjn_core_179 = ~(input_a[21] | input_a[24]);
  assign popcount31_1hjn_core_180 = ~(input_a[23] ^ input_a[19]);
  assign popcount31_1hjn_core_181 = ~input_a[5];
  assign popcount31_1hjn_core_182 = input_a[25] | input_a[11];
  assign popcount31_1hjn_core_183 = ~(input_a[30] & input_a[24]);
  assign popcount31_1hjn_core_185 = input_a[4] & input_a[30];
  assign popcount31_1hjn_core_186 = ~(input_a[1] | input_a[30]);
  assign popcount31_1hjn_core_189 = ~(input_a[25] & input_a[5]);
  assign popcount31_1hjn_core_190 = input_a[17] ^ input_a[17];
  assign popcount31_1hjn_core_191 = ~(input_a[12] & input_a[8]);
  assign popcount31_1hjn_core_192 = ~input_a[1];
  assign popcount31_1hjn_core_193 = ~(input_a[23] ^ input_a[0]);
  assign popcount31_1hjn_core_197 = input_a[12] | input_a[29];
  assign popcount31_1hjn_core_198 = input_a[1] | input_a[17];
  assign popcount31_1hjn_core_199 = input_a[3] | input_a[11];
  assign popcount31_1hjn_core_201 = ~(input_a[5] | input_a[10]);
  assign popcount31_1hjn_core_202 = input_a[11] | input_a[0];
  assign popcount31_1hjn_core_203 = input_a[3] ^ input_a[4];
  assign popcount31_1hjn_core_206 = ~(input_a[11] | input_a[15]);
  assign popcount31_1hjn_core_207 = input_a[19] & input_a[9];
  assign popcount31_1hjn_core_208 = ~(input_a[2] | input_a[18]);
  assign popcount31_1hjn_core_209 = ~input_a[7];
  assign popcount31_1hjn_core_211 = input_a[18] & input_a[24];
  assign popcount31_1hjn_core_212 = ~(input_a[27] | input_a[3]);
  assign popcount31_1hjn_core_214 = ~(input_a[22] ^ input_a[4]);
  assign popcount31_1hjn_core_215 = input_a[8] ^ input_a[3];
  assign popcount31_1hjn_core_217 = input_a[14] | input_a[14];

  assign popcount31_1hjn_out[0] = input_a[3];
  assign popcount31_1hjn_out[1] = 1'b0;
  assign popcount31_1hjn_out[2] = input_a[28];
  assign popcount31_1hjn_out[3] = input_a[26];
  assign popcount31_1hjn_out[4] = input_a[1];
endmodule