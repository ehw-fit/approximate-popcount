// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.61873
// WCE=25.0
// EP=0.971465%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_exvj(input [26:0] input_a, output [4:0] popcount27_exvj_out);
  wire popcount27_exvj_core_032;
  wire popcount27_exvj_core_033;
  wire popcount27_exvj_core_035;
  wire popcount27_exvj_core_037;
  wire popcount27_exvj_core_039;
  wire popcount27_exvj_core_041;
  wire popcount27_exvj_core_044;
  wire popcount27_exvj_core_045;
  wire popcount27_exvj_core_046;
  wire popcount27_exvj_core_048;
  wire popcount27_exvj_core_050;
  wire popcount27_exvj_core_053;
  wire popcount27_exvj_core_054;
  wire popcount27_exvj_core_055;
  wire popcount27_exvj_core_057;
  wire popcount27_exvj_core_058;
  wire popcount27_exvj_core_059_not;
  wire popcount27_exvj_core_060;
  wire popcount27_exvj_core_062;
  wire popcount27_exvj_core_064;
  wire popcount27_exvj_core_065;
  wire popcount27_exvj_core_066;
  wire popcount27_exvj_core_067;
  wire popcount27_exvj_core_068;
  wire popcount27_exvj_core_071;
  wire popcount27_exvj_core_073;
  wire popcount27_exvj_core_076;
  wire popcount27_exvj_core_079_not;
  wire popcount27_exvj_core_081;
  wire popcount27_exvj_core_083;
  wire popcount27_exvj_core_084;
  wire popcount27_exvj_core_085;
  wire popcount27_exvj_core_087;
  wire popcount27_exvj_core_088;
  wire popcount27_exvj_core_090;
  wire popcount27_exvj_core_092;
  wire popcount27_exvj_core_094;
  wire popcount27_exvj_core_095;
  wire popcount27_exvj_core_096;
  wire popcount27_exvj_core_097;
  wire popcount27_exvj_core_100;
  wire popcount27_exvj_core_101;
  wire popcount27_exvj_core_103;
  wire popcount27_exvj_core_105;
  wire popcount27_exvj_core_106;
  wire popcount27_exvj_core_107;
  wire popcount27_exvj_core_108;
  wire popcount27_exvj_core_109;
  wire popcount27_exvj_core_111;
  wire popcount27_exvj_core_112;
  wire popcount27_exvj_core_113;
  wire popcount27_exvj_core_114;
  wire popcount27_exvj_core_116;
  wire popcount27_exvj_core_117;
  wire popcount27_exvj_core_119;
  wire popcount27_exvj_core_120;
  wire popcount27_exvj_core_121;
  wire popcount27_exvj_core_122;
  wire popcount27_exvj_core_123;
  wire popcount27_exvj_core_124;
  wire popcount27_exvj_core_125;
  wire popcount27_exvj_core_128;
  wire popcount27_exvj_core_129;
  wire popcount27_exvj_core_130;
  wire popcount27_exvj_core_131;
  wire popcount27_exvj_core_132;
  wire popcount27_exvj_core_134;
  wire popcount27_exvj_core_136;
  wire popcount27_exvj_core_137;
  wire popcount27_exvj_core_140;
  wire popcount27_exvj_core_141;
  wire popcount27_exvj_core_143;
  wire popcount27_exvj_core_144_not;
  wire popcount27_exvj_core_147_not;
  wire popcount27_exvj_core_148;
  wire popcount27_exvj_core_149;
  wire popcount27_exvj_core_151;
  wire popcount27_exvj_core_152_not;
  wire popcount27_exvj_core_153;
  wire popcount27_exvj_core_154;
  wire popcount27_exvj_core_157;
  wire popcount27_exvj_core_159;
  wire popcount27_exvj_core_160;
  wire popcount27_exvj_core_161;
  wire popcount27_exvj_core_162;
  wire popcount27_exvj_core_163;
  wire popcount27_exvj_core_164;
  wire popcount27_exvj_core_167;
  wire popcount27_exvj_core_168;
  wire popcount27_exvj_core_170;
  wire popcount27_exvj_core_172;
  wire popcount27_exvj_core_173;
  wire popcount27_exvj_core_174;
  wire popcount27_exvj_core_175;
  wire popcount27_exvj_core_177;
  wire popcount27_exvj_core_179;
  wire popcount27_exvj_core_180;
  wire popcount27_exvj_core_181;
  wire popcount27_exvj_core_182;
  wire popcount27_exvj_core_183;
  wire popcount27_exvj_core_185;
  wire popcount27_exvj_core_186;
  wire popcount27_exvj_core_187;
  wire popcount27_exvj_core_188;
  wire popcount27_exvj_core_189;
  wire popcount27_exvj_core_190;
  wire popcount27_exvj_core_195;

  assign popcount27_exvj_core_032 = ~(input_a[20] | input_a[21]);
  assign popcount27_exvj_core_033 = ~(input_a[15] ^ input_a[11]);
  assign popcount27_exvj_core_035 = ~(input_a[15] & input_a[8]);
  assign popcount27_exvj_core_037 = input_a[13] & input_a[22];
  assign popcount27_exvj_core_039 = input_a[26] & input_a[20];
  assign popcount27_exvj_core_041 = input_a[25] ^ input_a[26];
  assign popcount27_exvj_core_044 = ~(input_a[10] | input_a[7]);
  assign popcount27_exvj_core_045 = input_a[2] ^ input_a[1];
  assign popcount27_exvj_core_046 = ~input_a[1];
  assign popcount27_exvj_core_048 = ~(input_a[8] & input_a[26]);
  assign popcount27_exvj_core_050 = ~(input_a[8] & input_a[18]);
  assign popcount27_exvj_core_053 = ~input_a[12];
  assign popcount27_exvj_core_054 = input_a[14] & input_a[2];
  assign popcount27_exvj_core_055 = input_a[8] ^ input_a[5];
  assign popcount27_exvj_core_057 = ~(input_a[6] | input_a[12]);
  assign popcount27_exvj_core_058 = ~(input_a[2] ^ input_a[16]);
  assign popcount27_exvj_core_059_not = ~input_a[20];
  assign popcount27_exvj_core_060 = input_a[15] | input_a[26];
  assign popcount27_exvj_core_062 = ~(input_a[0] ^ input_a[8]);
  assign popcount27_exvj_core_064 = ~input_a[4];
  assign popcount27_exvj_core_065 = ~(input_a[16] | input_a[10]);
  assign popcount27_exvj_core_066 = ~input_a[10];
  assign popcount27_exvj_core_067 = ~(input_a[2] ^ input_a[13]);
  assign popcount27_exvj_core_068 = input_a[0] | input_a[9];
  assign popcount27_exvj_core_071 = input_a[23] ^ input_a[16];
  assign popcount27_exvj_core_073 = input_a[22] | input_a[25];
  assign popcount27_exvj_core_076 = input_a[12] | input_a[25];
  assign popcount27_exvj_core_079_not = ~input_a[12];
  assign popcount27_exvj_core_081 = ~(input_a[25] & input_a[7]);
  assign popcount27_exvj_core_083 = ~(input_a[15] & input_a[2]);
  assign popcount27_exvj_core_084 = ~input_a[16];
  assign popcount27_exvj_core_085 = input_a[22] ^ input_a[22];
  assign popcount27_exvj_core_087 = ~(input_a[6] ^ input_a[16]);
  assign popcount27_exvj_core_088 = input_a[20] & input_a[15];
  assign popcount27_exvj_core_090 = ~(input_a[13] | input_a[18]);
  assign popcount27_exvj_core_092 = ~(input_a[0] ^ input_a[16]);
  assign popcount27_exvj_core_094 = ~(input_a[16] & input_a[22]);
  assign popcount27_exvj_core_095 = input_a[21] ^ input_a[26];
  assign popcount27_exvj_core_096 = ~(input_a[4] | input_a[10]);
  assign popcount27_exvj_core_097 = ~(input_a[8] ^ input_a[19]);
  assign popcount27_exvj_core_100 = input_a[9] | input_a[4];
  assign popcount27_exvj_core_101 = input_a[22] & input_a[14];
  assign popcount27_exvj_core_103 = ~(input_a[19] | input_a[11]);
  assign popcount27_exvj_core_105 = input_a[4] & input_a[3];
  assign popcount27_exvj_core_106 = input_a[9] | input_a[15];
  assign popcount27_exvj_core_107 = ~(input_a[26] ^ input_a[10]);
  assign popcount27_exvj_core_108 = ~input_a[5];
  assign popcount27_exvj_core_109 = ~(input_a[2] ^ input_a[26]);
  assign popcount27_exvj_core_111 = ~input_a[2];
  assign popcount27_exvj_core_112 = ~(input_a[11] | input_a[2]);
  assign popcount27_exvj_core_113 = ~(input_a[24] ^ input_a[19]);
  assign popcount27_exvj_core_114 = ~(input_a[20] | input_a[7]);
  assign popcount27_exvj_core_116 = input_a[14] ^ input_a[14];
  assign popcount27_exvj_core_117 = ~input_a[20];
  assign popcount27_exvj_core_119 = ~(input_a[22] | input_a[21]);
  assign popcount27_exvj_core_120 = input_a[1] | input_a[6];
  assign popcount27_exvj_core_121 = ~(input_a[15] ^ input_a[11]);
  assign popcount27_exvj_core_122 = input_a[19] ^ input_a[7];
  assign popcount27_exvj_core_123 = input_a[3] & input_a[24];
  assign popcount27_exvj_core_124 = ~(input_a[1] & input_a[0]);
  assign popcount27_exvj_core_125 = input_a[24] | input_a[1];
  assign popcount27_exvj_core_128 = ~input_a[5];
  assign popcount27_exvj_core_129 = ~(input_a[9] | input_a[3]);
  assign popcount27_exvj_core_130 = ~(input_a[1] | input_a[10]);
  assign popcount27_exvj_core_131 = ~(input_a[0] | input_a[12]);
  assign popcount27_exvj_core_132 = ~(input_a[15] ^ input_a[19]);
  assign popcount27_exvj_core_134 = input_a[22] & input_a[20];
  assign popcount27_exvj_core_136 = ~(input_a[24] | input_a[25]);
  assign popcount27_exvj_core_137 = ~(input_a[24] & input_a[9]);
  assign popcount27_exvj_core_140 = input_a[20] | input_a[14];
  assign popcount27_exvj_core_141 = input_a[22] | input_a[15];
  assign popcount27_exvj_core_143 = ~input_a[24];
  assign popcount27_exvj_core_144_not = ~input_a[11];
  assign popcount27_exvj_core_147_not = ~input_a[13];
  assign popcount27_exvj_core_148 = input_a[26] | input_a[13];
  assign popcount27_exvj_core_149 = input_a[23] | input_a[14];
  assign popcount27_exvj_core_151 = input_a[24] ^ input_a[2];
  assign popcount27_exvj_core_152_not = ~input_a[19];
  assign popcount27_exvj_core_153 = input_a[4] | input_a[10];
  assign popcount27_exvj_core_154 = ~(input_a[24] | input_a[16]);
  assign popcount27_exvj_core_157 = ~(input_a[22] & input_a[4]);
  assign popcount27_exvj_core_159 = ~input_a[25];
  assign popcount27_exvj_core_160 = input_a[17] ^ input_a[14];
  assign popcount27_exvj_core_161 = ~(input_a[15] | input_a[12]);
  assign popcount27_exvj_core_162 = ~(input_a[25] & input_a[11]);
  assign popcount27_exvj_core_163 = input_a[3] | input_a[10];
  assign popcount27_exvj_core_164 = ~(input_a[23] ^ input_a[1]);
  assign popcount27_exvj_core_167 = input_a[0] & input_a[17];
  assign popcount27_exvj_core_168 = ~(input_a[6] ^ input_a[17]);
  assign popcount27_exvj_core_170 = ~input_a[5];
  assign popcount27_exvj_core_172 = input_a[26] ^ input_a[22];
  assign popcount27_exvj_core_173 = ~input_a[14];
  assign popcount27_exvj_core_174 = ~(input_a[6] | input_a[9]);
  assign popcount27_exvj_core_175 = ~(input_a[20] ^ input_a[13]);
  assign popcount27_exvj_core_177 = input_a[2] ^ input_a[23];
  assign popcount27_exvj_core_179 = ~(input_a[18] & input_a[10]);
  assign popcount27_exvj_core_180 = ~(input_a[1] & input_a[19]);
  assign popcount27_exvj_core_181 = input_a[11] ^ input_a[23];
  assign popcount27_exvj_core_182 = ~input_a[19];
  assign popcount27_exvj_core_183 = ~(input_a[1] ^ input_a[18]);
  assign popcount27_exvj_core_185 = ~input_a[21];
  assign popcount27_exvj_core_186 = ~input_a[12];
  assign popcount27_exvj_core_187 = ~(input_a[24] ^ input_a[18]);
  assign popcount27_exvj_core_188 = ~(input_a[17] & input_a[18]);
  assign popcount27_exvj_core_189 = input_a[2] | input_a[9];
  assign popcount27_exvj_core_190 = ~input_a[4];
  assign popcount27_exvj_core_195 = input_a[13] & input_a[26];

  assign popcount27_exvj_out[0] = input_a[22];
  assign popcount27_exvj_out[1] = 1'b0;
  assign popcount27_exvj_out[2] = input_a[10];
  assign popcount27_exvj_out[3] = input_a[2];
  assign popcount27_exvj_out[4] = input_a[25];
endmodule