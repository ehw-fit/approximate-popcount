// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5794
// WCE=44.0
// EP=0.980625%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_xcpb(input [34:0] input_a, output [5:0] popcount35_xcpb_out);
  wire popcount35_xcpb_core_037;
  wire popcount35_xcpb_core_038;
  wire popcount35_xcpb_core_039;
  wire popcount35_xcpb_core_040;
  wire popcount35_xcpb_core_041;
  wire popcount35_xcpb_core_043;
  wire popcount35_xcpb_core_044;
  wire popcount35_xcpb_core_045;
  wire popcount35_xcpb_core_046;
  wire popcount35_xcpb_core_048;
  wire popcount35_xcpb_core_050;
  wire popcount35_xcpb_core_051;
  wire popcount35_xcpb_core_054;
  wire popcount35_xcpb_core_055;
  wire popcount35_xcpb_core_058;
  wire popcount35_xcpb_core_059;
  wire popcount35_xcpb_core_060;
  wire popcount35_xcpb_core_061;
  wire popcount35_xcpb_core_063;
  wire popcount35_xcpb_core_064;
  wire popcount35_xcpb_core_065;
  wire popcount35_xcpb_core_066;
  wire popcount35_xcpb_core_067;
  wire popcount35_xcpb_core_068;
  wire popcount35_xcpb_core_069;
  wire popcount35_xcpb_core_070;
  wire popcount35_xcpb_core_073;
  wire popcount35_xcpb_core_074;
  wire popcount35_xcpb_core_076;
  wire popcount35_xcpb_core_078;
  wire popcount35_xcpb_core_079;
  wire popcount35_xcpb_core_081;
  wire popcount35_xcpb_core_083;
  wire popcount35_xcpb_core_084;
  wire popcount35_xcpb_core_086;
  wire popcount35_xcpb_core_090;
  wire popcount35_xcpb_core_091;
  wire popcount35_xcpb_core_092;
  wire popcount35_xcpb_core_094;
  wire popcount35_xcpb_core_096;
  wire popcount35_xcpb_core_098;
  wire popcount35_xcpb_core_100;
  wire popcount35_xcpb_core_101;
  wire popcount35_xcpb_core_102;
  wire popcount35_xcpb_core_104;
  wire popcount35_xcpb_core_105;
  wire popcount35_xcpb_core_106;
  wire popcount35_xcpb_core_107;
  wire popcount35_xcpb_core_108_not;
  wire popcount35_xcpb_core_109;
  wire popcount35_xcpb_core_112;
  wire popcount35_xcpb_core_113;
  wire popcount35_xcpb_core_115;
  wire popcount35_xcpb_core_116;
  wire popcount35_xcpb_core_117;
  wire popcount35_xcpb_core_118;
  wire popcount35_xcpb_core_120;
  wire popcount35_xcpb_core_123;
  wire popcount35_xcpb_core_124;
  wire popcount35_xcpb_core_126;
  wire popcount35_xcpb_core_127;
  wire popcount35_xcpb_core_128;
  wire popcount35_xcpb_core_129;
  wire popcount35_xcpb_core_131_not;
  wire popcount35_xcpb_core_132;
  wire popcount35_xcpb_core_133;
  wire popcount35_xcpb_core_134;
  wire popcount35_xcpb_core_136;
  wire popcount35_xcpb_core_139;
  wire popcount35_xcpb_core_140;
  wire popcount35_xcpb_core_141;
  wire popcount35_xcpb_core_144;
  wire popcount35_xcpb_core_145;
  wire popcount35_xcpb_core_146;
  wire popcount35_xcpb_core_147;
  wire popcount35_xcpb_core_148;
  wire popcount35_xcpb_core_150;
  wire popcount35_xcpb_core_151;
  wire popcount35_xcpb_core_152;
  wire popcount35_xcpb_core_153;
  wire popcount35_xcpb_core_156;
  wire popcount35_xcpb_core_158;
  wire popcount35_xcpb_core_160;
  wire popcount35_xcpb_core_163;
  wire popcount35_xcpb_core_164;
  wire popcount35_xcpb_core_165;
  wire popcount35_xcpb_core_166;
  wire popcount35_xcpb_core_167;
  wire popcount35_xcpb_core_168;
  wire popcount35_xcpb_core_170;
  wire popcount35_xcpb_core_171;
  wire popcount35_xcpb_core_172;
  wire popcount35_xcpb_core_173;
  wire popcount35_xcpb_core_174;
  wire popcount35_xcpb_core_177;
  wire popcount35_xcpb_core_179;
  wire popcount35_xcpb_core_180;
  wire popcount35_xcpb_core_181;
  wire popcount35_xcpb_core_182;
  wire popcount35_xcpb_core_183;
  wire popcount35_xcpb_core_185;
  wire popcount35_xcpb_core_186;
  wire popcount35_xcpb_core_187;
  wire popcount35_xcpb_core_188;
  wire popcount35_xcpb_core_189;
  wire popcount35_xcpb_core_191;
  wire popcount35_xcpb_core_192;
  wire popcount35_xcpb_core_193;
  wire popcount35_xcpb_core_194;
  wire popcount35_xcpb_core_195;
  wire popcount35_xcpb_core_196;
  wire popcount35_xcpb_core_197;
  wire popcount35_xcpb_core_199;
  wire popcount35_xcpb_core_206;
  wire popcount35_xcpb_core_207;
  wire popcount35_xcpb_core_212;
  wire popcount35_xcpb_core_213;
  wire popcount35_xcpb_core_214;
  wire popcount35_xcpb_core_215;
  wire popcount35_xcpb_core_217;
  wire popcount35_xcpb_core_220;
  wire popcount35_xcpb_core_221;
  wire popcount35_xcpb_core_222;
  wire popcount35_xcpb_core_223;
  wire popcount35_xcpb_core_224;
  wire popcount35_xcpb_core_225;
  wire popcount35_xcpb_core_226;
  wire popcount35_xcpb_core_227;
  wire popcount35_xcpb_core_230;
  wire popcount35_xcpb_core_231;
  wire popcount35_xcpb_core_239;
  wire popcount35_xcpb_core_240;
  wire popcount35_xcpb_core_241;
  wire popcount35_xcpb_core_242;
  wire popcount35_xcpb_core_244;
  wire popcount35_xcpb_core_245;
  wire popcount35_xcpb_core_246;
  wire popcount35_xcpb_core_247;
  wire popcount35_xcpb_core_249;
  wire popcount35_xcpb_core_250;
  wire popcount35_xcpb_core_253;
  wire popcount35_xcpb_core_254;
  wire popcount35_xcpb_core_255;
  wire popcount35_xcpb_core_258;
  wire popcount35_xcpb_core_260;
  wire popcount35_xcpb_core_262;
  wire popcount35_xcpb_core_263;
  wire popcount35_xcpb_core_264;

  assign popcount35_xcpb_core_037 = ~(input_a[7] ^ input_a[4]);
  assign popcount35_xcpb_core_038 = input_a[20] | input_a[3];
  assign popcount35_xcpb_core_039 = input_a[31] & input_a[21];
  assign popcount35_xcpb_core_040 = ~input_a[14];
  assign popcount35_xcpb_core_041 = ~(input_a[24] | input_a[32]);
  assign popcount35_xcpb_core_043 = input_a[4] ^ input_a[1];
  assign popcount35_xcpb_core_044 = input_a[22] ^ input_a[29];
  assign popcount35_xcpb_core_045 = input_a[2] ^ input_a[3];
  assign popcount35_xcpb_core_046 = ~input_a[28];
  assign popcount35_xcpb_core_048 = ~(input_a[21] | input_a[19]);
  assign popcount35_xcpb_core_050 = ~input_a[25];
  assign popcount35_xcpb_core_051 = ~(input_a[32] | input_a[16]);
  assign popcount35_xcpb_core_054 = input_a[0] ^ input_a[0];
  assign popcount35_xcpb_core_055 = ~(input_a[11] ^ input_a[30]);
  assign popcount35_xcpb_core_058 = ~input_a[12];
  assign popcount35_xcpb_core_059 = ~input_a[11];
  assign popcount35_xcpb_core_060 = input_a[11] & input_a[27];
  assign popcount35_xcpb_core_061 = ~(input_a[0] | input_a[4]);
  assign popcount35_xcpb_core_063 = ~input_a[16];
  assign popcount35_xcpb_core_064 = input_a[17] | input_a[3];
  assign popcount35_xcpb_core_065 = input_a[2] | input_a[34];
  assign popcount35_xcpb_core_066 = ~(input_a[15] ^ input_a[9]);
  assign popcount35_xcpb_core_067 = ~input_a[34];
  assign popcount35_xcpb_core_068 = input_a[34] | input_a[30];
  assign popcount35_xcpb_core_069 = input_a[7] | input_a[1];
  assign popcount35_xcpb_core_070 = ~input_a[34];
  assign popcount35_xcpb_core_073 = input_a[2] & input_a[19];
  assign popcount35_xcpb_core_074 = ~input_a[0];
  assign popcount35_xcpb_core_076 = input_a[30] ^ input_a[26];
  assign popcount35_xcpb_core_078 = ~input_a[25];
  assign popcount35_xcpb_core_079 = input_a[23] & input_a[17];
  assign popcount35_xcpb_core_081 = input_a[19] & input_a[13];
  assign popcount35_xcpb_core_083 = ~(input_a[3] & input_a[18]);
  assign popcount35_xcpb_core_084 = ~(input_a[27] | input_a[20]);
  assign popcount35_xcpb_core_086 = input_a[15] | input_a[10];
  assign popcount35_xcpb_core_090 = ~(input_a[20] & input_a[0]);
  assign popcount35_xcpb_core_091 = ~input_a[1];
  assign popcount35_xcpb_core_092 = ~input_a[0];
  assign popcount35_xcpb_core_094 = input_a[34] & input_a[28];
  assign popcount35_xcpb_core_096 = input_a[0] ^ input_a[26];
  assign popcount35_xcpb_core_098 = ~(input_a[20] & input_a[33]);
  assign popcount35_xcpb_core_100 = input_a[12] | input_a[11];
  assign popcount35_xcpb_core_101 = ~(input_a[9] & input_a[33]);
  assign popcount35_xcpb_core_102 = ~(input_a[32] ^ input_a[29]);
  assign popcount35_xcpb_core_104 = ~input_a[10];
  assign popcount35_xcpb_core_105 = ~input_a[15];
  assign popcount35_xcpb_core_106 = ~(input_a[28] & input_a[10]);
  assign popcount35_xcpb_core_107 = input_a[31] ^ input_a[31];
  assign popcount35_xcpb_core_108_not = ~input_a[16];
  assign popcount35_xcpb_core_109 = ~(input_a[4] & input_a[9]);
  assign popcount35_xcpb_core_112 = ~(input_a[34] | input_a[22]);
  assign popcount35_xcpb_core_113 = input_a[6] | input_a[8];
  assign popcount35_xcpb_core_115 = input_a[21] | input_a[2];
  assign popcount35_xcpb_core_116 = input_a[28] | input_a[9];
  assign popcount35_xcpb_core_117 = ~(input_a[7] | input_a[3]);
  assign popcount35_xcpb_core_118 = input_a[3] & input_a[21];
  assign popcount35_xcpb_core_120 = ~input_a[23];
  assign popcount35_xcpb_core_123 = input_a[26] & input_a[11];
  assign popcount35_xcpb_core_124 = ~(input_a[14] ^ input_a[23]);
  assign popcount35_xcpb_core_126 = input_a[2] | input_a[1];
  assign popcount35_xcpb_core_127 = input_a[7] | input_a[31];
  assign popcount35_xcpb_core_128 = ~(input_a[33] & input_a[34]);
  assign popcount35_xcpb_core_129 = ~(input_a[16] & input_a[19]);
  assign popcount35_xcpb_core_131_not = ~input_a[4];
  assign popcount35_xcpb_core_132 = ~(input_a[10] | input_a[30]);
  assign popcount35_xcpb_core_133 = ~(input_a[19] ^ input_a[2]);
  assign popcount35_xcpb_core_134 = input_a[11] | input_a[5];
  assign popcount35_xcpb_core_136 = input_a[5] & input_a[29];
  assign popcount35_xcpb_core_139 = ~(input_a[3] & input_a[33]);
  assign popcount35_xcpb_core_140 = ~input_a[22];
  assign popcount35_xcpb_core_141 = input_a[11] | input_a[24];
  assign popcount35_xcpb_core_144 = input_a[11] ^ input_a[7];
  assign popcount35_xcpb_core_145 = ~(input_a[14] | input_a[3]);
  assign popcount35_xcpb_core_146 = ~(input_a[5] ^ input_a[10]);
  assign popcount35_xcpb_core_147 = input_a[28] ^ input_a[0];
  assign popcount35_xcpb_core_148 = ~(input_a[7] & input_a[23]);
  assign popcount35_xcpb_core_150 = input_a[8] ^ input_a[16];
  assign popcount35_xcpb_core_151 = ~(input_a[26] & input_a[10]);
  assign popcount35_xcpb_core_152 = ~(input_a[10] ^ input_a[12]);
  assign popcount35_xcpb_core_153 = ~(input_a[4] & input_a[6]);
  assign popcount35_xcpb_core_156 = input_a[16] ^ input_a[21];
  assign popcount35_xcpb_core_158 = ~(input_a[14] | input_a[4]);
  assign popcount35_xcpb_core_160 = ~input_a[27];
  assign popcount35_xcpb_core_163 = input_a[9] & input_a[30];
  assign popcount35_xcpb_core_164 = input_a[27] ^ input_a[1];
  assign popcount35_xcpb_core_165 = input_a[0] & input_a[6];
  assign popcount35_xcpb_core_166 = ~(input_a[11] | input_a[19]);
  assign popcount35_xcpb_core_167 = input_a[16] | input_a[2];
  assign popcount35_xcpb_core_168 = ~(input_a[32] ^ input_a[27]);
  assign popcount35_xcpb_core_170 = ~input_a[2];
  assign popcount35_xcpb_core_171 = ~input_a[24];
  assign popcount35_xcpb_core_172 = input_a[13] ^ input_a[8];
  assign popcount35_xcpb_core_173 = ~(input_a[20] & input_a[26]);
  assign popcount35_xcpb_core_174 = ~(input_a[24] ^ input_a[19]);
  assign popcount35_xcpb_core_177 = ~(input_a[10] ^ input_a[16]);
  assign popcount35_xcpb_core_179 = ~input_a[16];
  assign popcount35_xcpb_core_180 = ~(input_a[28] | input_a[19]);
  assign popcount35_xcpb_core_181 = ~(input_a[7] | input_a[8]);
  assign popcount35_xcpb_core_182 = input_a[31] | input_a[16];
  assign popcount35_xcpb_core_183 = input_a[18] | input_a[27];
  assign popcount35_xcpb_core_185 = ~(input_a[3] & input_a[4]);
  assign popcount35_xcpb_core_186 = input_a[5] ^ input_a[34];
  assign popcount35_xcpb_core_187 = ~(input_a[14] ^ input_a[18]);
  assign popcount35_xcpb_core_188 = ~(input_a[15] ^ input_a[1]);
  assign popcount35_xcpb_core_189 = ~(input_a[18] | input_a[33]);
  assign popcount35_xcpb_core_191 = ~(input_a[10] ^ input_a[32]);
  assign popcount35_xcpb_core_192 = ~(input_a[9] ^ input_a[23]);
  assign popcount35_xcpb_core_193 = ~input_a[22];
  assign popcount35_xcpb_core_194 = ~(input_a[15] ^ input_a[28]);
  assign popcount35_xcpb_core_195 = ~(input_a[32] & input_a[21]);
  assign popcount35_xcpb_core_196 = input_a[10] & input_a[14];
  assign popcount35_xcpb_core_197 = ~(input_a[2] & input_a[10]);
  assign popcount35_xcpb_core_199 = input_a[21] & input_a[27];
  assign popcount35_xcpb_core_206 = input_a[24] | input_a[26];
  assign popcount35_xcpb_core_207 = ~(input_a[11] ^ input_a[5]);
  assign popcount35_xcpb_core_212 = ~(input_a[27] | input_a[34]);
  assign popcount35_xcpb_core_213 = ~(input_a[0] ^ input_a[7]);
  assign popcount35_xcpb_core_214 = ~(input_a[25] ^ input_a[19]);
  assign popcount35_xcpb_core_215 = input_a[14] | input_a[13];
  assign popcount35_xcpb_core_217 = ~input_a[10];
  assign popcount35_xcpb_core_220 = ~input_a[21];
  assign popcount35_xcpb_core_221 = input_a[33] | input_a[32];
  assign popcount35_xcpb_core_222 = ~(input_a[3] ^ input_a[33]);
  assign popcount35_xcpb_core_223 = input_a[24] | input_a[17];
  assign popcount35_xcpb_core_224 = input_a[6] & input_a[0];
  assign popcount35_xcpb_core_225 = input_a[17] | input_a[7];
  assign popcount35_xcpb_core_226 = input_a[18] ^ input_a[26];
  assign popcount35_xcpb_core_227 = ~(input_a[27] & input_a[31]);
  assign popcount35_xcpb_core_230 = ~(input_a[19] & input_a[21]);
  assign popcount35_xcpb_core_231 = ~(input_a[7] & input_a[34]);
  assign popcount35_xcpb_core_239 = input_a[12] & input_a[22];
  assign popcount35_xcpb_core_240 = ~input_a[16];
  assign popcount35_xcpb_core_241 = input_a[8] & input_a[27];
  assign popcount35_xcpb_core_242 = input_a[11] | input_a[24];
  assign popcount35_xcpb_core_244 = ~(input_a[7] | input_a[5]);
  assign popcount35_xcpb_core_245 = ~(input_a[29] ^ input_a[12]);
  assign popcount35_xcpb_core_246 = input_a[21] | input_a[8];
  assign popcount35_xcpb_core_247 = ~(input_a[34] & input_a[5]);
  assign popcount35_xcpb_core_249 = ~(input_a[14] & input_a[19]);
  assign popcount35_xcpb_core_250 = ~input_a[6];
  assign popcount35_xcpb_core_253 = ~(input_a[33] ^ input_a[15]);
  assign popcount35_xcpb_core_254 = input_a[32] | input_a[0];
  assign popcount35_xcpb_core_255 = input_a[23] ^ input_a[2];
  assign popcount35_xcpb_core_258 = ~(input_a[11] ^ input_a[28]);
  assign popcount35_xcpb_core_260 = input_a[17] | input_a[0];
  assign popcount35_xcpb_core_262 = ~(input_a[11] & input_a[17]);
  assign popcount35_xcpb_core_263 = input_a[13] & input_a[3];
  assign popcount35_xcpb_core_264 = ~(input_a[6] & input_a[15]);

  assign popcount35_xcpb_out[0] = 1'b1;
  assign popcount35_xcpb_out[1] = input_a[9];
  assign popcount35_xcpb_out[2] = input_a[2];
  assign popcount35_xcpb_out[3] = 1'b1;
  assign popcount35_xcpb_out[4] = 1'b0;
  assign popcount35_xcpb_out[5] = input_a[26];
endmodule