// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.89143
// WCE=20.0
// EP=0.893656%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_ab6g(input [35:0] input_a, output [5:0] popcount36_ab6g_out);
  wire popcount36_ab6g_core_038;
  wire popcount36_ab6g_core_039;
  wire popcount36_ab6g_core_040;
  wire popcount36_ab6g_core_041;
  wire popcount36_ab6g_core_043;
  wire popcount36_ab6g_core_044;
  wire popcount36_ab6g_core_045;
  wire popcount36_ab6g_core_046;
  wire popcount36_ab6g_core_047;
  wire popcount36_ab6g_core_048;
  wire popcount36_ab6g_core_050;
  wire popcount36_ab6g_core_051;
  wire popcount36_ab6g_core_052;
  wire popcount36_ab6g_core_055;
  wire popcount36_ab6g_core_056;
  wire popcount36_ab6g_core_057;
  wire popcount36_ab6g_core_058;
  wire popcount36_ab6g_core_059;
  wire popcount36_ab6g_core_061;
  wire popcount36_ab6g_core_062;
  wire popcount36_ab6g_core_063;
  wire popcount36_ab6g_core_065;
  wire popcount36_ab6g_core_068;
  wire popcount36_ab6g_core_069;
  wire popcount36_ab6g_core_070;
  wire popcount36_ab6g_core_071;
  wire popcount36_ab6g_core_072;
  wire popcount36_ab6g_core_073;
  wire popcount36_ab6g_core_074;
  wire popcount36_ab6g_core_075;
  wire popcount36_ab6g_core_078;
  wire popcount36_ab6g_core_082;
  wire popcount36_ab6g_core_083;
  wire popcount36_ab6g_core_085;
  wire popcount36_ab6g_core_090;
  wire popcount36_ab6g_core_091;
  wire popcount36_ab6g_core_092;
  wire popcount36_ab6g_core_093;
  wire popcount36_ab6g_core_095;
  wire popcount36_ab6g_core_097;
  wire popcount36_ab6g_core_098;
  wire popcount36_ab6g_core_099;
  wire popcount36_ab6g_core_100;
  wire popcount36_ab6g_core_102;
  wire popcount36_ab6g_core_104;
  wire popcount36_ab6g_core_105;
  wire popcount36_ab6g_core_107;
  wire popcount36_ab6g_core_109;
  wire popcount36_ab6g_core_111;
  wire popcount36_ab6g_core_113;
  wire popcount36_ab6g_core_115;
  wire popcount36_ab6g_core_116;
  wire popcount36_ab6g_core_117;
  wire popcount36_ab6g_core_118;
  wire popcount36_ab6g_core_119;
  wire popcount36_ab6g_core_120;
  wire popcount36_ab6g_core_122;
  wire popcount36_ab6g_core_123;
  wire popcount36_ab6g_core_124;
  wire popcount36_ab6g_core_125;
  wire popcount36_ab6g_core_126;
  wire popcount36_ab6g_core_130;
  wire popcount36_ab6g_core_133;
  wire popcount36_ab6g_core_134;
  wire popcount36_ab6g_core_135;
  wire popcount36_ab6g_core_136;
  wire popcount36_ab6g_core_139;
  wire popcount36_ab6g_core_140;
  wire popcount36_ab6g_core_141;
  wire popcount36_ab6g_core_146;
  wire popcount36_ab6g_core_147;
  wire popcount36_ab6g_core_148_not;
  wire popcount36_ab6g_core_149;
  wire popcount36_ab6g_core_151;
  wire popcount36_ab6g_core_152;
  wire popcount36_ab6g_core_154;
  wire popcount36_ab6g_core_155;
  wire popcount36_ab6g_core_156;
  wire popcount36_ab6g_core_158;
  wire popcount36_ab6g_core_160_not;
  wire popcount36_ab6g_core_161;
  wire popcount36_ab6g_core_162;
  wire popcount36_ab6g_core_164;
  wire popcount36_ab6g_core_165;
  wire popcount36_ab6g_core_167_not;
  wire popcount36_ab6g_core_168;
  wire popcount36_ab6g_core_169;
  wire popcount36_ab6g_core_171;
  wire popcount36_ab6g_core_172;
  wire popcount36_ab6g_core_174;
  wire popcount36_ab6g_core_175;
  wire popcount36_ab6g_core_177;
  wire popcount36_ab6g_core_179;
  wire popcount36_ab6g_core_181;
  wire popcount36_ab6g_core_184;
  wire popcount36_ab6g_core_185;
  wire popcount36_ab6g_core_186_not;
  wire popcount36_ab6g_core_187;
  wire popcount36_ab6g_core_191;
  wire popcount36_ab6g_core_192;
  wire popcount36_ab6g_core_194;
  wire popcount36_ab6g_core_195;
  wire popcount36_ab6g_core_196;
  wire popcount36_ab6g_core_198;
  wire popcount36_ab6g_core_199;
  wire popcount36_ab6g_core_202;
  wire popcount36_ab6g_core_203;
  wire popcount36_ab6g_core_207;
  wire popcount36_ab6g_core_208;
  wire popcount36_ab6g_core_210;
  wire popcount36_ab6g_core_211;
  wire popcount36_ab6g_core_212;
  wire popcount36_ab6g_core_213;
  wire popcount36_ab6g_core_214;
  wire popcount36_ab6g_core_215;
  wire popcount36_ab6g_core_216;
  wire popcount36_ab6g_core_217;
  wire popcount36_ab6g_core_220;
  wire popcount36_ab6g_core_222;
  wire popcount36_ab6g_core_224;
  wire popcount36_ab6g_core_227;
  wire popcount36_ab6g_core_228;
  wire popcount36_ab6g_core_229;
  wire popcount36_ab6g_core_230;
  wire popcount36_ab6g_core_231;
  wire popcount36_ab6g_core_233;
  wire popcount36_ab6g_core_235;
  wire popcount36_ab6g_core_236;
  wire popcount36_ab6g_core_237;
  wire popcount36_ab6g_core_239;
  wire popcount36_ab6g_core_241;
  wire popcount36_ab6g_core_242;
  wire popcount36_ab6g_core_244;
  wire popcount36_ab6g_core_247;
  wire popcount36_ab6g_core_250;
  wire popcount36_ab6g_core_251;
  wire popcount36_ab6g_core_252;
  wire popcount36_ab6g_core_253;
  wire popcount36_ab6g_core_254;
  wire popcount36_ab6g_core_255;
  wire popcount36_ab6g_core_257;
  wire popcount36_ab6g_core_258;
  wire popcount36_ab6g_core_260;
  wire popcount36_ab6g_core_261;
  wire popcount36_ab6g_core_262;
  wire popcount36_ab6g_core_263;
  wire popcount36_ab6g_core_264_not;
  wire popcount36_ab6g_core_266;
  wire popcount36_ab6g_core_268;
  wire popcount36_ab6g_core_270;
  wire popcount36_ab6g_core_271;
  wire popcount36_ab6g_core_272;
  wire popcount36_ab6g_core_273;
  wire popcount36_ab6g_core_274;
  wire popcount36_ab6g_core_275;
  wire popcount36_ab6g_core_276;

  assign popcount36_ab6g_core_038 = ~(input_a[11] & input_a[24]);
  assign popcount36_ab6g_core_039 = ~(input_a[2] & input_a[35]);
  assign popcount36_ab6g_core_040 = input_a[23] ^ input_a[21];
  assign popcount36_ab6g_core_041 = ~input_a[24];
  assign popcount36_ab6g_core_043 = ~(input_a[30] | input_a[27]);
  assign popcount36_ab6g_core_044 = input_a[11] | input_a[16];
  assign popcount36_ab6g_core_045 = input_a[31] ^ input_a[1];
  assign popcount36_ab6g_core_046 = input_a[23] & input_a[17];
  assign popcount36_ab6g_core_047 = input_a[23] ^ input_a[28];
  assign popcount36_ab6g_core_048 = ~(input_a[4] | input_a[4]);
  assign popcount36_ab6g_core_050 = ~(input_a[5] & input_a[10]);
  assign popcount36_ab6g_core_051 = input_a[23] ^ input_a[14];
  assign popcount36_ab6g_core_052 = ~(input_a[24] ^ input_a[12]);
  assign popcount36_ab6g_core_055 = input_a[14] & input_a[27];
  assign popcount36_ab6g_core_056 = ~(input_a[35] ^ input_a[8]);
  assign popcount36_ab6g_core_057 = ~input_a[0];
  assign popcount36_ab6g_core_058 = input_a[19] | input_a[11];
  assign popcount36_ab6g_core_059 = ~(input_a[11] | input_a[33]);
  assign popcount36_ab6g_core_061 = input_a[35] ^ input_a[33];
  assign popcount36_ab6g_core_062 = input_a[7] | input_a[30];
  assign popcount36_ab6g_core_063 = ~input_a[7];
  assign popcount36_ab6g_core_065 = input_a[15] & input_a[8];
  assign popcount36_ab6g_core_068 = input_a[29] | input_a[23];
  assign popcount36_ab6g_core_069 = input_a[35] ^ input_a[8];
  assign popcount36_ab6g_core_070 = input_a[17] | input_a[5];
  assign popcount36_ab6g_core_071 = input_a[16] | input_a[4];
  assign popcount36_ab6g_core_072 = ~(input_a[32] ^ input_a[8]);
  assign popcount36_ab6g_core_073 = input_a[31] ^ input_a[21];
  assign popcount36_ab6g_core_074 = input_a[26] | input_a[19];
  assign popcount36_ab6g_core_075 = input_a[12] ^ input_a[19];
  assign popcount36_ab6g_core_078 = ~(input_a[16] ^ input_a[27]);
  assign popcount36_ab6g_core_082 = input_a[13] ^ input_a[24];
  assign popcount36_ab6g_core_083 = ~input_a[11];
  assign popcount36_ab6g_core_085 = ~input_a[12];
  assign popcount36_ab6g_core_090 = ~(input_a[0] & input_a[23]);
  assign popcount36_ab6g_core_091 = ~(input_a[13] & input_a[20]);
  assign popcount36_ab6g_core_092 = input_a[0] & input_a[31];
  assign popcount36_ab6g_core_093 = ~(input_a[29] & input_a[8]);
  assign popcount36_ab6g_core_095 = ~(input_a[10] | input_a[7]);
  assign popcount36_ab6g_core_097 = ~(input_a[32] ^ input_a[9]);
  assign popcount36_ab6g_core_098 = ~(input_a[34] & input_a[3]);
  assign popcount36_ab6g_core_099 = input_a[13] & input_a[18];
  assign popcount36_ab6g_core_100 = input_a[12] ^ input_a[33];
  assign popcount36_ab6g_core_102 = input_a[12] | input_a[17];
  assign popcount36_ab6g_core_104 = input_a[22] & input_a[3];
  assign popcount36_ab6g_core_105 = ~input_a[6];
  assign popcount36_ab6g_core_107 = input_a[9] ^ input_a[2];
  assign popcount36_ab6g_core_109 = input_a[10] ^ input_a[9];
  assign popcount36_ab6g_core_111 = input_a[19] ^ input_a[18];
  assign popcount36_ab6g_core_113 = input_a[30] & input_a[19];
  assign popcount36_ab6g_core_115 = ~(input_a[28] | input_a[22]);
  assign popcount36_ab6g_core_116 = ~(input_a[0] ^ input_a[22]);
  assign popcount36_ab6g_core_117 = ~input_a[2];
  assign popcount36_ab6g_core_118 = input_a[31] ^ input_a[15];
  assign popcount36_ab6g_core_119 = ~input_a[20];
  assign popcount36_ab6g_core_120 = input_a[16] & input_a[15];
  assign popcount36_ab6g_core_122 = ~input_a[25];
  assign popcount36_ab6g_core_123 = ~(input_a[25] ^ input_a[32]);
  assign popcount36_ab6g_core_124 = input_a[30] | input_a[4];
  assign popcount36_ab6g_core_125 = ~input_a[24];
  assign popcount36_ab6g_core_126 = ~input_a[27];
  assign popcount36_ab6g_core_130 = input_a[27] ^ input_a[11];
  assign popcount36_ab6g_core_133 = input_a[31] | input_a[5];
  assign popcount36_ab6g_core_134 = ~input_a[6];
  assign popcount36_ab6g_core_135 = input_a[25] ^ input_a[34];
  assign popcount36_ab6g_core_136 = ~(input_a[32] & input_a[34]);
  assign popcount36_ab6g_core_139 = input_a[6] | input_a[2];
  assign popcount36_ab6g_core_140 = input_a[2] ^ input_a[31];
  assign popcount36_ab6g_core_141 = ~(input_a[11] & input_a[11]);
  assign popcount36_ab6g_core_146 = input_a[16] & input_a[5];
  assign popcount36_ab6g_core_147 = input_a[1] ^ input_a[19];
  assign popcount36_ab6g_core_148_not = ~input_a[31];
  assign popcount36_ab6g_core_149 = input_a[35] | input_a[28];
  assign popcount36_ab6g_core_151 = ~(input_a[6] & input_a[5]);
  assign popcount36_ab6g_core_152 = ~input_a[11];
  assign popcount36_ab6g_core_154 = input_a[30] & input_a[0];
  assign popcount36_ab6g_core_155 = ~(input_a[30] & input_a[5]);
  assign popcount36_ab6g_core_156 = ~(input_a[23] ^ input_a[35]);
  assign popcount36_ab6g_core_158 = ~(input_a[9] & input_a[17]);
  assign popcount36_ab6g_core_160_not = ~input_a[2];
  assign popcount36_ab6g_core_161 = input_a[1] | input_a[32];
  assign popcount36_ab6g_core_162 = input_a[15] & input_a[19];
  assign popcount36_ab6g_core_164 = ~input_a[2];
  assign popcount36_ab6g_core_165 = ~input_a[3];
  assign popcount36_ab6g_core_167_not = ~input_a[2];
  assign popcount36_ab6g_core_168 = input_a[4] & input_a[34];
  assign popcount36_ab6g_core_169 = ~(input_a[13] & input_a[12]);
  assign popcount36_ab6g_core_171 = ~(input_a[34] | input_a[25]);
  assign popcount36_ab6g_core_172 = input_a[3] | input_a[11];
  assign popcount36_ab6g_core_174 = ~(input_a[0] & input_a[2]);
  assign popcount36_ab6g_core_175 = ~input_a[12];
  assign popcount36_ab6g_core_177 = ~input_a[15];
  assign popcount36_ab6g_core_179 = ~(input_a[29] | input_a[2]);
  assign popcount36_ab6g_core_181 = ~(input_a[23] ^ input_a[13]);
  assign popcount36_ab6g_core_184 = ~input_a[25];
  assign popcount36_ab6g_core_185 = ~input_a[20];
  assign popcount36_ab6g_core_186_not = ~input_a[24];
  assign popcount36_ab6g_core_187 = input_a[14] ^ input_a[16];
  assign popcount36_ab6g_core_191 = input_a[2] & input_a[12];
  assign popcount36_ab6g_core_192 = input_a[17] & input_a[5];
  assign popcount36_ab6g_core_194 = ~(input_a[22] & input_a[23]);
  assign popcount36_ab6g_core_195 = input_a[8] & input_a[5];
  assign popcount36_ab6g_core_196 = ~(input_a[0] & input_a[33]);
  assign popcount36_ab6g_core_198 = ~(input_a[25] | input_a[23]);
  assign popcount36_ab6g_core_199 = input_a[27] | input_a[12];
  assign popcount36_ab6g_core_202 = input_a[30] | input_a[23];
  assign popcount36_ab6g_core_203 = input_a[7] & input_a[31];
  assign popcount36_ab6g_core_207 = ~(input_a[31] ^ input_a[21]);
  assign popcount36_ab6g_core_208 = ~(input_a[29] ^ input_a[29]);
  assign popcount36_ab6g_core_210 = input_a[13] ^ input_a[30];
  assign popcount36_ab6g_core_211 = input_a[22] ^ input_a[16];
  assign popcount36_ab6g_core_212 = input_a[14] ^ input_a[29];
  assign popcount36_ab6g_core_213 = ~input_a[18];
  assign popcount36_ab6g_core_214 = input_a[8] | input_a[23];
  assign popcount36_ab6g_core_215 = ~input_a[27];
  assign popcount36_ab6g_core_216 = input_a[34] | input_a[17];
  assign popcount36_ab6g_core_217 = ~(input_a[15] & input_a[25]);
  assign popcount36_ab6g_core_220 = ~(input_a[22] ^ input_a[29]);
  assign popcount36_ab6g_core_222 = input_a[12] ^ input_a[5];
  assign popcount36_ab6g_core_224 = ~(input_a[30] & input_a[17]);
  assign popcount36_ab6g_core_227 = input_a[14] | input_a[34];
  assign popcount36_ab6g_core_228 = input_a[33] ^ input_a[34];
  assign popcount36_ab6g_core_229 = ~input_a[17];
  assign popcount36_ab6g_core_230 = ~(input_a[2] ^ input_a[30]);
  assign popcount36_ab6g_core_231 = ~input_a[27];
  assign popcount36_ab6g_core_233 = input_a[8] | input_a[35];
  assign popcount36_ab6g_core_235 = input_a[35] ^ input_a[32];
  assign popcount36_ab6g_core_236 = ~(input_a[16] & input_a[30]);
  assign popcount36_ab6g_core_237 = input_a[6] ^ input_a[25];
  assign popcount36_ab6g_core_239 = input_a[30] | input_a[6];
  assign popcount36_ab6g_core_241 = ~(input_a[2] ^ input_a[12]);
  assign popcount36_ab6g_core_242 = input_a[19] ^ input_a[25];
  assign popcount36_ab6g_core_244 = input_a[22] ^ input_a[1];
  assign popcount36_ab6g_core_247 = ~input_a[27];
  assign popcount36_ab6g_core_250 = ~(input_a[12] & input_a[13]);
  assign popcount36_ab6g_core_251 = ~(input_a[35] ^ input_a[1]);
  assign popcount36_ab6g_core_252 = ~(input_a[33] | input_a[1]);
  assign popcount36_ab6g_core_253 = input_a[3] ^ input_a[17];
  assign popcount36_ab6g_core_254 = input_a[30] | input_a[30];
  assign popcount36_ab6g_core_255 = ~(input_a[18] | input_a[8]);
  assign popcount36_ab6g_core_257 = input_a[1] | input_a[6];
  assign popcount36_ab6g_core_258 = input_a[10] | input_a[7];
  assign popcount36_ab6g_core_260 = ~(input_a[22] ^ input_a[26]);
  assign popcount36_ab6g_core_261 = ~input_a[26];
  assign popcount36_ab6g_core_262 = input_a[26] & input_a[5];
  assign popcount36_ab6g_core_263 = ~(input_a[19] ^ input_a[2]);
  assign popcount36_ab6g_core_264_not = ~input_a[11];
  assign popcount36_ab6g_core_266 = ~input_a[27];
  assign popcount36_ab6g_core_268 = input_a[18] | input_a[25];
  assign popcount36_ab6g_core_270 = ~(input_a[16] | input_a[11]);
  assign popcount36_ab6g_core_271 = ~(input_a[4] | input_a[23]);
  assign popcount36_ab6g_core_272 = input_a[0] ^ input_a[7];
  assign popcount36_ab6g_core_273 = ~(input_a[15] ^ input_a[7]);
  assign popcount36_ab6g_core_274 = ~(input_a[28] | input_a[0]);
  assign popcount36_ab6g_core_275 = input_a[20] & input_a[11];
  assign popcount36_ab6g_core_276 = input_a[26] ^ input_a[34];

  assign popcount36_ab6g_out[0] = input_a[14];
  assign popcount36_ab6g_out[1] = 1'b0;
  assign popcount36_ab6g_out[2] = 1'b1;
  assign popcount36_ab6g_out[3] = 1'b0;
  assign popcount36_ab6g_out[4] = 1'b1;
  assign popcount36_ab6g_out[5] = 1'b0;
endmodule