// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=10.5
// WCE=24.0
// EP=0.999978%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_6bx8(input [27:0] input_a, output [4:0] popcount28_6bx8_out);
  wire popcount28_6bx8_core_030;
  wire popcount28_6bx8_core_032;
  wire popcount28_6bx8_core_033;
  wire popcount28_6bx8_core_035;
  wire popcount28_6bx8_core_037;
  wire popcount28_6bx8_core_038;
  wire popcount28_6bx8_core_039;
  wire popcount28_6bx8_core_040;
  wire popcount28_6bx8_core_041;
  wire popcount28_6bx8_core_042;
  wire popcount28_6bx8_core_045;
  wire popcount28_6bx8_core_046;
  wire popcount28_6bx8_core_047;
  wire popcount28_6bx8_core_049;
  wire popcount28_6bx8_core_052;
  wire popcount28_6bx8_core_053;
  wire popcount28_6bx8_core_055;
  wire popcount28_6bx8_core_058;
  wire popcount28_6bx8_core_059_not;
  wire popcount28_6bx8_core_062;
  wire popcount28_6bx8_core_063;
  wire popcount28_6bx8_core_064;
  wire popcount28_6bx8_core_065;
  wire popcount28_6bx8_core_066;
  wire popcount28_6bx8_core_068;
  wire popcount28_6bx8_core_070;
  wire popcount28_6bx8_core_071;
  wire popcount28_6bx8_core_072;
  wire popcount28_6bx8_core_074;
  wire popcount28_6bx8_core_075;
  wire popcount28_6bx8_core_080;
  wire popcount28_6bx8_core_082;
  wire popcount28_6bx8_core_084;
  wire popcount28_6bx8_core_085;
  wire popcount28_6bx8_core_088;
  wire popcount28_6bx8_core_089;
  wire popcount28_6bx8_core_090;
  wire popcount28_6bx8_core_091;
  wire popcount28_6bx8_core_092;
  wire popcount28_6bx8_core_093;
  wire popcount28_6bx8_core_094;
  wire popcount28_6bx8_core_098;
  wire popcount28_6bx8_core_099;
  wire popcount28_6bx8_core_100;
  wire popcount28_6bx8_core_102;
  wire popcount28_6bx8_core_103;
  wire popcount28_6bx8_core_105;
  wire popcount28_6bx8_core_108;
  wire popcount28_6bx8_core_111;
  wire popcount28_6bx8_core_116;
  wire popcount28_6bx8_core_117;
  wire popcount28_6bx8_core_118;
  wire popcount28_6bx8_core_120;
  wire popcount28_6bx8_core_123;
  wire popcount28_6bx8_core_124;
  wire popcount28_6bx8_core_125;
  wire popcount28_6bx8_core_126;
  wire popcount28_6bx8_core_127;
  wire popcount28_6bx8_core_128;
  wire popcount28_6bx8_core_130;
  wire popcount28_6bx8_core_131;
  wire popcount28_6bx8_core_132;
  wire popcount28_6bx8_core_135;
  wire popcount28_6bx8_core_136;
  wire popcount28_6bx8_core_137;
  wire popcount28_6bx8_core_138;
  wire popcount28_6bx8_core_141;
  wire popcount28_6bx8_core_142;
  wire popcount28_6bx8_core_143;
  wire popcount28_6bx8_core_144;
  wire popcount28_6bx8_core_145;
  wire popcount28_6bx8_core_146;
  wire popcount28_6bx8_core_147;
  wire popcount28_6bx8_core_148;
  wire popcount28_6bx8_core_150;
  wire popcount28_6bx8_core_152;
  wire popcount28_6bx8_core_156;
  wire popcount28_6bx8_core_159;
  wire popcount28_6bx8_core_160;
  wire popcount28_6bx8_core_165;
  wire popcount28_6bx8_core_166;
  wire popcount28_6bx8_core_167_not;
  wire popcount28_6bx8_core_169;
  wire popcount28_6bx8_core_170_not;
  wire popcount28_6bx8_core_171;
  wire popcount28_6bx8_core_172;
  wire popcount28_6bx8_core_173;
  wire popcount28_6bx8_core_175;
  wire popcount28_6bx8_core_177;
  wire popcount28_6bx8_core_179;
  wire popcount28_6bx8_core_180;
  wire popcount28_6bx8_core_181;
  wire popcount28_6bx8_core_182;
  wire popcount28_6bx8_core_183;
  wire popcount28_6bx8_core_184;
  wire popcount28_6bx8_core_185;
  wire popcount28_6bx8_core_186;
  wire popcount28_6bx8_core_187;
  wire popcount28_6bx8_core_188_not;
  wire popcount28_6bx8_core_191;
  wire popcount28_6bx8_core_193;
  wire popcount28_6bx8_core_195;
  wire popcount28_6bx8_core_198;
  wire popcount28_6bx8_core_200;

  assign popcount28_6bx8_core_030 = ~(input_a[10] | input_a[13]);
  assign popcount28_6bx8_core_032 = input_a[25] ^ input_a[0];
  assign popcount28_6bx8_core_033 = input_a[2] ^ input_a[22];
  assign popcount28_6bx8_core_035 = ~input_a[15];
  assign popcount28_6bx8_core_037 = ~(input_a[23] ^ input_a[2]);
  assign popcount28_6bx8_core_038 = ~(input_a[6] | input_a[20]);
  assign popcount28_6bx8_core_039 = input_a[17] ^ input_a[5];
  assign popcount28_6bx8_core_040 = ~(input_a[11] ^ input_a[6]);
  assign popcount28_6bx8_core_041 = input_a[2] & input_a[3];
  assign popcount28_6bx8_core_042 = ~(input_a[0] | input_a[12]);
  assign popcount28_6bx8_core_045 = ~input_a[2];
  assign popcount28_6bx8_core_046 = ~input_a[0];
  assign popcount28_6bx8_core_047 = input_a[10] ^ input_a[1];
  assign popcount28_6bx8_core_049 = ~(input_a[26] & input_a[16]);
  assign popcount28_6bx8_core_052 = input_a[20] | input_a[13];
  assign popcount28_6bx8_core_053 = ~input_a[3];
  assign popcount28_6bx8_core_055 = ~(input_a[11] ^ input_a[10]);
  assign popcount28_6bx8_core_058 = input_a[5] & input_a[17];
  assign popcount28_6bx8_core_059_not = ~input_a[9];
  assign popcount28_6bx8_core_062 = ~(input_a[17] & input_a[11]);
  assign popcount28_6bx8_core_063 = input_a[20] & input_a[21];
  assign popcount28_6bx8_core_064 = ~(input_a[14] & input_a[20]);
  assign popcount28_6bx8_core_065 = input_a[20] & input_a[24];
  assign popcount28_6bx8_core_066 = input_a[12] | input_a[5];
  assign popcount28_6bx8_core_068 = input_a[13] ^ input_a[25];
  assign popcount28_6bx8_core_070 = ~(input_a[9] & input_a[25]);
  assign popcount28_6bx8_core_071 = input_a[14] | input_a[22];
  assign popcount28_6bx8_core_072 = ~(input_a[0] & input_a[16]);
  assign popcount28_6bx8_core_074 = ~(input_a[18] ^ input_a[15]);
  assign popcount28_6bx8_core_075 = ~(input_a[21] | input_a[15]);
  assign popcount28_6bx8_core_080 = ~input_a[16];
  assign popcount28_6bx8_core_082 = input_a[25] ^ input_a[20];
  assign popcount28_6bx8_core_084 = input_a[23] | input_a[21];
  assign popcount28_6bx8_core_085 = ~(input_a[1] & input_a[6]);
  assign popcount28_6bx8_core_088 = ~(input_a[20] ^ input_a[0]);
  assign popcount28_6bx8_core_089 = ~input_a[23];
  assign popcount28_6bx8_core_090 = input_a[24] ^ input_a[16];
  assign popcount28_6bx8_core_091 = input_a[16] & input_a[0];
  assign popcount28_6bx8_core_092 = ~(input_a[24] ^ input_a[27]);
  assign popcount28_6bx8_core_093 = input_a[10] ^ input_a[20];
  assign popcount28_6bx8_core_094 = input_a[25] | input_a[0];
  assign popcount28_6bx8_core_098 = input_a[5] & input_a[25];
  assign popcount28_6bx8_core_099 = input_a[27] | input_a[21];
  assign popcount28_6bx8_core_100 = ~(input_a[16] | input_a[14]);
  assign popcount28_6bx8_core_102 = input_a[22] | input_a[19];
  assign popcount28_6bx8_core_103 = ~(input_a[7] ^ input_a[15]);
  assign popcount28_6bx8_core_105 = ~(input_a[8] | input_a[1]);
  assign popcount28_6bx8_core_108 = input_a[2] | input_a[3];
  assign popcount28_6bx8_core_111 = ~input_a[14];
  assign popcount28_6bx8_core_116 = input_a[11] ^ input_a[27];
  assign popcount28_6bx8_core_117 = ~input_a[5];
  assign popcount28_6bx8_core_118 = ~(input_a[21] ^ input_a[13]);
  assign popcount28_6bx8_core_120 = ~(input_a[27] ^ input_a[15]);
  assign popcount28_6bx8_core_123 = ~(input_a[25] ^ input_a[17]);
  assign popcount28_6bx8_core_124 = input_a[11] | input_a[25];
  assign popcount28_6bx8_core_125 = input_a[0] ^ input_a[17];
  assign popcount28_6bx8_core_126 = input_a[25] & input_a[23];
  assign popcount28_6bx8_core_127 = ~(input_a[27] & input_a[22]);
  assign popcount28_6bx8_core_128 = ~input_a[1];
  assign popcount28_6bx8_core_130 = input_a[10] & input_a[19];
  assign popcount28_6bx8_core_131 = ~(input_a[25] & input_a[7]);
  assign popcount28_6bx8_core_132 = ~(input_a[5] & input_a[13]);
  assign popcount28_6bx8_core_135 = ~(input_a[13] ^ input_a[19]);
  assign popcount28_6bx8_core_136 = ~(input_a[11] ^ input_a[21]);
  assign popcount28_6bx8_core_137 = input_a[5] | input_a[0];
  assign popcount28_6bx8_core_138 = input_a[13] ^ input_a[1];
  assign popcount28_6bx8_core_141 = input_a[13] & input_a[9];
  assign popcount28_6bx8_core_142 = ~input_a[20];
  assign popcount28_6bx8_core_143 = input_a[5] | input_a[22];
  assign popcount28_6bx8_core_144 = ~(input_a[26] | input_a[22]);
  assign popcount28_6bx8_core_145 = ~(input_a[26] | input_a[14]);
  assign popcount28_6bx8_core_146 = ~(input_a[1] ^ input_a[24]);
  assign popcount28_6bx8_core_147 = input_a[15] & input_a[4];
  assign popcount28_6bx8_core_148 = input_a[3] ^ input_a[18];
  assign popcount28_6bx8_core_150 = input_a[17] | input_a[23];
  assign popcount28_6bx8_core_152 = input_a[2] | input_a[3];
  assign popcount28_6bx8_core_156 = ~(input_a[5] ^ input_a[25]);
  assign popcount28_6bx8_core_159 = ~input_a[0];
  assign popcount28_6bx8_core_160 = ~(input_a[4] & input_a[15]);
  assign popcount28_6bx8_core_165 = input_a[7] ^ input_a[8];
  assign popcount28_6bx8_core_166 = input_a[9] & input_a[0];
  assign popcount28_6bx8_core_167_not = ~input_a[21];
  assign popcount28_6bx8_core_169 = ~(input_a[13] ^ input_a[6]);
  assign popcount28_6bx8_core_170_not = ~input_a[18];
  assign popcount28_6bx8_core_171 = input_a[3] | input_a[1];
  assign popcount28_6bx8_core_172 = input_a[16] | input_a[10];
  assign popcount28_6bx8_core_173 = input_a[24] & input_a[9];
  assign popcount28_6bx8_core_175 = ~(input_a[25] & input_a[3]);
  assign popcount28_6bx8_core_177 = input_a[27] | input_a[6];
  assign popcount28_6bx8_core_179 = ~(input_a[5] & input_a[0]);
  assign popcount28_6bx8_core_180 = input_a[15] | input_a[22];
  assign popcount28_6bx8_core_181 = input_a[17] & input_a[17];
  assign popcount28_6bx8_core_182 = ~(input_a[4] ^ input_a[3]);
  assign popcount28_6bx8_core_183 = ~(input_a[18] & input_a[15]);
  assign popcount28_6bx8_core_184 = ~(input_a[16] ^ input_a[1]);
  assign popcount28_6bx8_core_185 = input_a[17] ^ input_a[11];
  assign popcount28_6bx8_core_186 = ~(input_a[25] ^ input_a[9]);
  assign popcount28_6bx8_core_187 = input_a[16] & input_a[14];
  assign popcount28_6bx8_core_188_not = ~input_a[3];
  assign popcount28_6bx8_core_191 = ~input_a[13];
  assign popcount28_6bx8_core_193 = input_a[0] ^ input_a[1];
  assign popcount28_6bx8_core_195 = input_a[18] & input_a[26];
  assign popcount28_6bx8_core_198 = ~input_a[22];
  assign popcount28_6bx8_core_200 = ~(input_a[7] & input_a[27]);

  assign popcount28_6bx8_out[0] = input_a[18];
  assign popcount28_6bx8_out[1] = 1'b0;
  assign popcount28_6bx8_out[2] = 1'b0;
  assign popcount28_6bx8_out[3] = 1'b1;
  assign popcount28_6bx8_out[4] = 1'b1;
endmodule