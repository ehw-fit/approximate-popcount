// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.39291
// WCE=14.0
// EP=0.870702%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount24_3wel(input [23:0] input_a, output [4:0] popcount24_3wel_out);
  wire popcount24_3wel_core_026;
  wire popcount24_3wel_core_027;
  wire popcount24_3wel_core_028;
  wire popcount24_3wel_core_029;
  wire popcount24_3wel_core_030;
  wire popcount24_3wel_core_031;
  wire popcount24_3wel_core_032;
  wire popcount24_3wel_core_034;
  wire popcount24_3wel_core_035;
  wire popcount24_3wel_core_036;
  wire popcount24_3wel_core_037;
  wire popcount24_3wel_core_038;
  wire popcount24_3wel_core_040;
  wire popcount24_3wel_core_042;
  wire popcount24_3wel_core_046;
  wire popcount24_3wel_core_047;
  wire popcount24_3wel_core_051;
  wire popcount24_3wel_core_053;
  wire popcount24_3wel_core_054;
  wire popcount24_3wel_core_055;
  wire popcount24_3wel_core_056;
  wire popcount24_3wel_core_058;
  wire popcount24_3wel_core_060;
  wire popcount24_3wel_core_064;
  wire popcount24_3wel_core_065;
  wire popcount24_3wel_core_066;
  wire popcount24_3wel_core_068;
  wire popcount24_3wel_core_069;
  wire popcount24_3wel_core_075;
  wire popcount24_3wel_core_076;
  wire popcount24_3wel_core_077;
  wire popcount24_3wel_core_079;
  wire popcount24_3wel_core_081;
  wire popcount24_3wel_core_082;
  wire popcount24_3wel_core_088;
  wire popcount24_3wel_core_089;
  wire popcount24_3wel_core_090;
  wire popcount24_3wel_core_091;
  wire popcount24_3wel_core_092;
  wire popcount24_3wel_core_093;
  wire popcount24_3wel_core_095_not;
  wire popcount24_3wel_core_096;
  wire popcount24_3wel_core_097;
  wire popcount24_3wel_core_098;
  wire popcount24_3wel_core_100;
  wire popcount24_3wel_core_101_not;
  wire popcount24_3wel_core_102;
  wire popcount24_3wel_core_103;
  wire popcount24_3wel_core_105;
  wire popcount24_3wel_core_106;
  wire popcount24_3wel_core_107;
  wire popcount24_3wel_core_109;
  wire popcount24_3wel_core_112;
  wire popcount24_3wel_core_113_not;
  wire popcount24_3wel_core_115;
  wire popcount24_3wel_core_117;
  wire popcount24_3wel_core_119;
  wire popcount24_3wel_core_125;
  wire popcount24_3wel_core_126;
  wire popcount24_3wel_core_128;
  wire popcount24_3wel_core_129;
  wire popcount24_3wel_core_131;
  wire popcount24_3wel_core_133;
  wire popcount24_3wel_core_136;
  wire popcount24_3wel_core_139_not;
  wire popcount24_3wel_core_140;
  wire popcount24_3wel_core_142;
  wire popcount24_3wel_core_143;
  wire popcount24_3wel_core_144;
  wire popcount24_3wel_core_146;
  wire popcount24_3wel_core_147;
  wire popcount24_3wel_core_149;
  wire popcount24_3wel_core_150;
  wire popcount24_3wel_core_151;
  wire popcount24_3wel_core_153;
  wire popcount24_3wel_core_155;
  wire popcount24_3wel_core_156;
  wire popcount24_3wel_core_157_not;
  wire popcount24_3wel_core_160;
  wire popcount24_3wel_core_161;
  wire popcount24_3wel_core_164;
  wire popcount24_3wel_core_165_not;
  wire popcount24_3wel_core_166;
  wire popcount24_3wel_core_167_not;
  wire popcount24_3wel_core_171;
  wire popcount24_3wel_core_172;
  wire popcount24_3wel_core_175;
  wire popcount24_3wel_core_177;

  assign popcount24_3wel_core_026 = ~(input_a[1] ^ input_a[12]);
  assign popcount24_3wel_core_027 = input_a[11] | input_a[10];
  assign popcount24_3wel_core_028 = ~(input_a[7] ^ input_a[14]);
  assign popcount24_3wel_core_029 = input_a[21] | input_a[9];
  assign popcount24_3wel_core_030 = input_a[20] ^ input_a[5];
  assign popcount24_3wel_core_031 = input_a[0] & input_a[16];
  assign popcount24_3wel_core_032 = ~(input_a[20] & input_a[4]);
  assign popcount24_3wel_core_034 = ~(input_a[4] ^ input_a[15]);
  assign popcount24_3wel_core_035 = ~input_a[16];
  assign popcount24_3wel_core_036 = input_a[3] & input_a[23];
  assign popcount24_3wel_core_037 = input_a[8] | input_a[6];
  assign popcount24_3wel_core_038 = input_a[4] ^ input_a[19];
  assign popcount24_3wel_core_040 = ~(input_a[11] ^ input_a[9]);
  assign popcount24_3wel_core_042 = ~input_a[17];
  assign popcount24_3wel_core_046 = ~input_a[16];
  assign popcount24_3wel_core_047 = ~(input_a[8] ^ input_a[23]);
  assign popcount24_3wel_core_051 = ~(input_a[1] | input_a[17]);
  assign popcount24_3wel_core_053 = ~(input_a[3] & input_a[18]);
  assign popcount24_3wel_core_054 = ~(input_a[14] | input_a[12]);
  assign popcount24_3wel_core_055 = input_a[7] ^ input_a[15];
  assign popcount24_3wel_core_056 = ~input_a[4];
  assign popcount24_3wel_core_058 = input_a[18] ^ input_a[16];
  assign popcount24_3wel_core_060 = ~(input_a[8] | input_a[22]);
  assign popcount24_3wel_core_064 = ~(input_a[18] | input_a[14]);
  assign popcount24_3wel_core_065 = ~(input_a[9] & input_a[4]);
  assign popcount24_3wel_core_066 = input_a[6] | input_a[10];
  assign popcount24_3wel_core_068 = ~(input_a[10] | input_a[17]);
  assign popcount24_3wel_core_069 = input_a[10] ^ input_a[21];
  assign popcount24_3wel_core_075 = input_a[0] ^ input_a[7];
  assign popcount24_3wel_core_076 = input_a[14] ^ input_a[8];
  assign popcount24_3wel_core_077 = input_a[13] & input_a[17];
  assign popcount24_3wel_core_079 = input_a[11] & input_a[4];
  assign popcount24_3wel_core_081 = input_a[1] ^ input_a[21];
  assign popcount24_3wel_core_082 = input_a[13] | input_a[17];
  assign popcount24_3wel_core_088 = ~input_a[2];
  assign popcount24_3wel_core_089 = input_a[10] ^ input_a[4];
  assign popcount24_3wel_core_090 = ~(input_a[8] & input_a[11]);
  assign popcount24_3wel_core_091 = ~(input_a[21] ^ input_a[2]);
  assign popcount24_3wel_core_092 = ~(input_a[10] ^ input_a[2]);
  assign popcount24_3wel_core_093 = ~input_a[18];
  assign popcount24_3wel_core_095_not = ~input_a[14];
  assign popcount24_3wel_core_096 = input_a[10] & input_a[21];
  assign popcount24_3wel_core_097 = ~(input_a[9] & input_a[12]);
  assign popcount24_3wel_core_098 = input_a[16] ^ input_a[8];
  assign popcount24_3wel_core_100 = ~(input_a[12] & input_a[0]);
  assign popcount24_3wel_core_101_not = ~input_a[15];
  assign popcount24_3wel_core_102 = input_a[20] & input_a[19];
  assign popcount24_3wel_core_103 = ~(input_a[20] | input_a[14]);
  assign popcount24_3wel_core_105 = ~input_a[16];
  assign popcount24_3wel_core_106 = ~(input_a[9] | input_a[4]);
  assign popcount24_3wel_core_107 = ~(input_a[3] | input_a[2]);
  assign popcount24_3wel_core_109 = ~(input_a[4] & input_a[8]);
  assign popcount24_3wel_core_112 = input_a[17] & input_a[9];
  assign popcount24_3wel_core_113_not = ~input_a[5];
  assign popcount24_3wel_core_115 = ~(input_a[22] ^ input_a[4]);
  assign popcount24_3wel_core_117 = ~(input_a[17] & input_a[2]);
  assign popcount24_3wel_core_119 = ~input_a[13];
  assign popcount24_3wel_core_125 = ~(input_a[8] | input_a[11]);
  assign popcount24_3wel_core_126 = ~(input_a[0] ^ input_a[8]);
  assign popcount24_3wel_core_128 = input_a[5] | input_a[15];
  assign popcount24_3wel_core_129 = input_a[1] & input_a[14];
  assign popcount24_3wel_core_131 = ~(input_a[22] | input_a[13]);
  assign popcount24_3wel_core_133 = ~(input_a[15] ^ input_a[3]);
  assign popcount24_3wel_core_136 = input_a[6] | input_a[14];
  assign popcount24_3wel_core_139_not = ~input_a[22];
  assign popcount24_3wel_core_140 = ~(input_a[19] & input_a[20]);
  assign popcount24_3wel_core_142 = ~(input_a[4] ^ input_a[9]);
  assign popcount24_3wel_core_143 = ~input_a[1];
  assign popcount24_3wel_core_144 = ~(input_a[4] & input_a[20]);
  assign popcount24_3wel_core_146 = ~(input_a[10] | input_a[10]);
  assign popcount24_3wel_core_147 = ~(input_a[21] | input_a[23]);
  assign popcount24_3wel_core_149 = ~(input_a[1] ^ input_a[8]);
  assign popcount24_3wel_core_150 = input_a[10] & input_a[3];
  assign popcount24_3wel_core_151 = ~(input_a[9] & input_a[21]);
  assign popcount24_3wel_core_153 = ~(input_a[23] & input_a[15]);
  assign popcount24_3wel_core_155 = ~(input_a[23] | input_a[5]);
  assign popcount24_3wel_core_156 = input_a[13] & input_a[0];
  assign popcount24_3wel_core_157_not = ~input_a[1];
  assign popcount24_3wel_core_160 = input_a[13] & input_a[1];
  assign popcount24_3wel_core_161 = ~(input_a[9] & input_a[11]);
  assign popcount24_3wel_core_164 = ~(input_a[4] & input_a[16]);
  assign popcount24_3wel_core_165_not = ~input_a[6];
  assign popcount24_3wel_core_166 = ~(input_a[20] ^ input_a[3]);
  assign popcount24_3wel_core_167_not = ~input_a[16];
  assign popcount24_3wel_core_171 = ~input_a[14];
  assign popcount24_3wel_core_172 = input_a[11] & input_a[8];
  assign popcount24_3wel_core_175 = input_a[6] & input_a[8];
  assign popcount24_3wel_core_177 = input_a[22] & input_a[9];

  assign popcount24_3wel_out[0] = 1'b1;
  assign popcount24_3wel_out[1] = 1'b1;
  assign popcount24_3wel_out[2] = input_a[20];
  assign popcount24_3wel_out[3] = 1'b1;
  assign popcount24_3wel_out[4] = 1'b0;
endmodule