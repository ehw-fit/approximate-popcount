// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.59507
// WCE=27.0
// EP=0.973691%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_95r9(input [32:0] input_a, output [5:0] popcount33_95r9_out);
  wire popcount33_95r9_core_036;
  wire popcount33_95r9_core_037;
  wire popcount33_95r9_core_039;
  wire popcount33_95r9_core_041;
  wire popcount33_95r9_core_044;
  wire popcount33_95r9_core_045;
  wire popcount33_95r9_core_048;
  wire popcount33_95r9_core_050;
  wire popcount33_95r9_core_052;
  wire popcount33_95r9_core_053;
  wire popcount33_95r9_core_055;
  wire popcount33_95r9_core_056;
  wire popcount33_95r9_core_057;
  wire popcount33_95r9_core_058;
  wire popcount33_95r9_core_060;
  wire popcount33_95r9_core_061;
  wire popcount33_95r9_core_062;
  wire popcount33_95r9_core_063;
  wire popcount33_95r9_core_065;
  wire popcount33_95r9_core_068;
  wire popcount33_95r9_core_069;
  wire popcount33_95r9_core_072;
  wire popcount33_95r9_core_074;
  wire popcount33_95r9_core_075;
  wire popcount33_95r9_core_076;
  wire popcount33_95r9_core_077;
  wire popcount33_95r9_core_080;
  wire popcount33_95r9_core_081;
  wire popcount33_95r9_core_083;
  wire popcount33_95r9_core_085;
  wire popcount33_95r9_core_086;
  wire popcount33_95r9_core_087;
  wire popcount33_95r9_core_088;
  wire popcount33_95r9_core_089;
  wire popcount33_95r9_core_090;
  wire popcount33_95r9_core_091;
  wire popcount33_95r9_core_092;
  wire popcount33_95r9_core_095;
  wire popcount33_95r9_core_097;
  wire popcount33_95r9_core_100;
  wire popcount33_95r9_core_101;
  wire popcount33_95r9_core_102;
  wire popcount33_95r9_core_103;
  wire popcount33_95r9_core_105;
  wire popcount33_95r9_core_108;
  wire popcount33_95r9_core_114;
  wire popcount33_95r9_core_115;
  wire popcount33_95r9_core_116;
  wire popcount33_95r9_core_117;
  wire popcount33_95r9_core_118;
  wire popcount33_95r9_core_119;
  wire popcount33_95r9_core_122;
  wire popcount33_95r9_core_124;
  wire popcount33_95r9_core_125;
  wire popcount33_95r9_core_126;
  wire popcount33_95r9_core_127;
  wire popcount33_95r9_core_128;
  wire popcount33_95r9_core_129;
  wire popcount33_95r9_core_130;
  wire popcount33_95r9_core_131;
  wire popcount33_95r9_core_135;
  wire popcount33_95r9_core_137;
  wire popcount33_95r9_core_141;
  wire popcount33_95r9_core_142;
  wire popcount33_95r9_core_143;
  wire popcount33_95r9_core_144;
  wire popcount33_95r9_core_145;
  wire popcount33_95r9_core_147;
  wire popcount33_95r9_core_148;
  wire popcount33_95r9_core_153;
  wire popcount33_95r9_core_154;
  wire popcount33_95r9_core_155;
  wire popcount33_95r9_core_156;
  wire popcount33_95r9_core_157;
  wire popcount33_95r9_core_158;
  wire popcount33_95r9_core_159;
  wire popcount33_95r9_core_160;
  wire popcount33_95r9_core_162;
  wire popcount33_95r9_core_163;
  wire popcount33_95r9_core_164;
  wire popcount33_95r9_core_165;
  wire popcount33_95r9_core_166;
  wire popcount33_95r9_core_170;
  wire popcount33_95r9_core_171;
  wire popcount33_95r9_core_173;
  wire popcount33_95r9_core_175;
  wire popcount33_95r9_core_176;
  wire popcount33_95r9_core_178;
  wire popcount33_95r9_core_180;
  wire popcount33_95r9_core_181;
  wire popcount33_95r9_core_183;
  wire popcount33_95r9_core_184;
  wire popcount33_95r9_core_185;
  wire popcount33_95r9_core_187;
  wire popcount33_95r9_core_188;
  wire popcount33_95r9_core_190;
  wire popcount33_95r9_core_192;
  wire popcount33_95r9_core_193;
  wire popcount33_95r9_core_195;
  wire popcount33_95r9_core_196;
  wire popcount33_95r9_core_197;
  wire popcount33_95r9_core_199;
  wire popcount33_95r9_core_200;
  wire popcount33_95r9_core_201;
  wire popcount33_95r9_core_202;
  wire popcount33_95r9_core_204;
  wire popcount33_95r9_core_205;
  wire popcount33_95r9_core_209;
  wire popcount33_95r9_core_210;
  wire popcount33_95r9_core_214;
  wire popcount33_95r9_core_215;
  wire popcount33_95r9_core_216;
  wire popcount33_95r9_core_218;
  wire popcount33_95r9_core_219;
  wire popcount33_95r9_core_222;
  wire popcount33_95r9_core_223;
  wire popcount33_95r9_core_225;
  wire popcount33_95r9_core_227;
  wire popcount33_95r9_core_228;
  wire popcount33_95r9_core_232;
  wire popcount33_95r9_core_233;
  wire popcount33_95r9_core_234;
  wire popcount33_95r9_core_236;
  wire popcount33_95r9_core_238;

  assign popcount33_95r9_core_036 = ~(input_a[25] ^ input_a[1]);
  assign popcount33_95r9_core_037 = input_a[17] | input_a[13];
  assign popcount33_95r9_core_039 = ~(input_a[12] ^ input_a[2]);
  assign popcount33_95r9_core_041 = input_a[28] ^ input_a[5];
  assign popcount33_95r9_core_044 = ~(input_a[14] & input_a[32]);
  assign popcount33_95r9_core_045 = ~(input_a[21] & input_a[25]);
  assign popcount33_95r9_core_048 = ~input_a[28];
  assign popcount33_95r9_core_050 = ~input_a[26];
  assign popcount33_95r9_core_052 = ~(input_a[24] ^ input_a[20]);
  assign popcount33_95r9_core_053 = ~input_a[12];
  assign popcount33_95r9_core_055 = ~(input_a[27] & input_a[23]);
  assign popcount33_95r9_core_056 = ~(input_a[27] & input_a[21]);
  assign popcount33_95r9_core_057 = ~(input_a[2] & input_a[1]);
  assign popcount33_95r9_core_058 = input_a[29] | input_a[30];
  assign popcount33_95r9_core_060 = input_a[12] ^ input_a[25];
  assign popcount33_95r9_core_061 = ~input_a[6];
  assign popcount33_95r9_core_062 = input_a[6] & input_a[14];
  assign popcount33_95r9_core_063 = input_a[9] ^ input_a[13];
  assign popcount33_95r9_core_065 = input_a[30] & input_a[22];
  assign popcount33_95r9_core_068 = input_a[27] ^ input_a[12];
  assign popcount33_95r9_core_069 = ~(input_a[10] & input_a[23]);
  assign popcount33_95r9_core_072 = ~(input_a[32] | input_a[7]);
  assign popcount33_95r9_core_074 = input_a[1] ^ input_a[17];
  assign popcount33_95r9_core_075 = input_a[32] | input_a[17];
  assign popcount33_95r9_core_076 = ~(input_a[2] | input_a[0]);
  assign popcount33_95r9_core_077 = input_a[29] ^ input_a[20];
  assign popcount33_95r9_core_080 = ~(input_a[1] & input_a[26]);
  assign popcount33_95r9_core_081 = ~input_a[24];
  assign popcount33_95r9_core_083 = input_a[11] | input_a[5];
  assign popcount33_95r9_core_085 = ~input_a[32];
  assign popcount33_95r9_core_086 = input_a[26] & input_a[10];
  assign popcount33_95r9_core_087 = ~(input_a[8] & input_a[10]);
  assign popcount33_95r9_core_088 = input_a[16] & input_a[4];
  assign popcount33_95r9_core_089 = ~(input_a[2] | input_a[29]);
  assign popcount33_95r9_core_090 = ~(input_a[17] ^ input_a[23]);
  assign popcount33_95r9_core_091 = input_a[2] ^ input_a[2];
  assign popcount33_95r9_core_092 = input_a[22] ^ input_a[6];
  assign popcount33_95r9_core_095 = ~(input_a[6] | input_a[28]);
  assign popcount33_95r9_core_097 = input_a[27] & input_a[8];
  assign popcount33_95r9_core_100 = input_a[23] ^ input_a[10];
  assign popcount33_95r9_core_101 = ~(input_a[28] ^ input_a[7]);
  assign popcount33_95r9_core_102 = ~(input_a[29] & input_a[13]);
  assign popcount33_95r9_core_103 = ~(input_a[3] ^ input_a[9]);
  assign popcount33_95r9_core_105 = ~(input_a[24] ^ input_a[20]);
  assign popcount33_95r9_core_108 = input_a[31] ^ input_a[20];
  assign popcount33_95r9_core_114 = ~(input_a[4] & input_a[17]);
  assign popcount33_95r9_core_115 = ~(input_a[4] | input_a[5]);
  assign popcount33_95r9_core_116 = input_a[13] & input_a[23];
  assign popcount33_95r9_core_117 = input_a[7] ^ input_a[10];
  assign popcount33_95r9_core_118 = ~(input_a[28] | input_a[31]);
  assign popcount33_95r9_core_119 = ~input_a[17];
  assign popcount33_95r9_core_122 = input_a[24] ^ input_a[17];
  assign popcount33_95r9_core_124 = ~(input_a[25] & input_a[2]);
  assign popcount33_95r9_core_125 = ~(input_a[5] & input_a[3]);
  assign popcount33_95r9_core_126 = input_a[26] | input_a[18];
  assign popcount33_95r9_core_127 = ~(input_a[29] | input_a[31]);
  assign popcount33_95r9_core_128 = ~(input_a[0] & input_a[21]);
  assign popcount33_95r9_core_129 = input_a[12] | input_a[15];
  assign popcount33_95r9_core_130 = ~(input_a[4] ^ input_a[17]);
  assign popcount33_95r9_core_131 = input_a[27] | input_a[2];
  assign popcount33_95r9_core_135 = input_a[4] & input_a[17];
  assign popcount33_95r9_core_137 = input_a[5] & input_a[24];
  assign popcount33_95r9_core_141 = ~input_a[20];
  assign popcount33_95r9_core_142 = ~input_a[32];
  assign popcount33_95r9_core_143 = input_a[5] ^ input_a[16];
  assign popcount33_95r9_core_144 = input_a[9] ^ input_a[18];
  assign popcount33_95r9_core_145 = input_a[13] | input_a[1];
  assign popcount33_95r9_core_147 = input_a[0] ^ input_a[31];
  assign popcount33_95r9_core_148 = input_a[18] ^ input_a[25];
  assign popcount33_95r9_core_153 = ~(input_a[26] & input_a[23]);
  assign popcount33_95r9_core_154 = input_a[31] & input_a[10];
  assign popcount33_95r9_core_155 = input_a[28] | input_a[3];
  assign popcount33_95r9_core_156 = input_a[6] | input_a[23];
  assign popcount33_95r9_core_157 = ~(input_a[24] | input_a[15]);
  assign popcount33_95r9_core_158 = ~(input_a[6] | input_a[21]);
  assign popcount33_95r9_core_159 = input_a[28] ^ input_a[30];
  assign popcount33_95r9_core_160 = ~(input_a[26] ^ input_a[7]);
  assign popcount33_95r9_core_162 = input_a[20] | input_a[6];
  assign popcount33_95r9_core_163 = ~(input_a[32] ^ input_a[3]);
  assign popcount33_95r9_core_164 = ~(input_a[0] ^ input_a[29]);
  assign popcount33_95r9_core_165 = ~input_a[23];
  assign popcount33_95r9_core_166 = input_a[18] & input_a[5];
  assign popcount33_95r9_core_170 = input_a[2] | input_a[1];
  assign popcount33_95r9_core_171 = ~(input_a[13] | input_a[13]);
  assign popcount33_95r9_core_173 = ~(input_a[23] ^ input_a[2]);
  assign popcount33_95r9_core_175 = ~input_a[2];
  assign popcount33_95r9_core_176 = ~(input_a[11] ^ input_a[12]);
  assign popcount33_95r9_core_178 = ~(input_a[25] & input_a[18]);
  assign popcount33_95r9_core_180 = ~(input_a[15] & input_a[4]);
  assign popcount33_95r9_core_181 = input_a[5] ^ input_a[10];
  assign popcount33_95r9_core_183 = ~(input_a[23] | input_a[4]);
  assign popcount33_95r9_core_184 = ~input_a[19];
  assign popcount33_95r9_core_185 = ~input_a[26];
  assign popcount33_95r9_core_187 = input_a[0] | input_a[23];
  assign popcount33_95r9_core_188 = input_a[13] ^ input_a[23];
  assign popcount33_95r9_core_190 = ~(input_a[30] ^ input_a[25]);
  assign popcount33_95r9_core_192 = ~input_a[1];
  assign popcount33_95r9_core_193 = ~(input_a[13] & input_a[26]);
  assign popcount33_95r9_core_195 = ~(input_a[2] | input_a[18]);
  assign popcount33_95r9_core_196 = ~input_a[24];
  assign popcount33_95r9_core_197 = ~(input_a[14] ^ input_a[10]);
  assign popcount33_95r9_core_199 = input_a[5] & input_a[30];
  assign popcount33_95r9_core_200 = input_a[30] & input_a[13];
  assign popcount33_95r9_core_201 = ~input_a[4];
  assign popcount33_95r9_core_202 = input_a[14] ^ input_a[20];
  assign popcount33_95r9_core_204 = ~(input_a[11] ^ input_a[2]);
  assign popcount33_95r9_core_205 = input_a[19] ^ input_a[2];
  assign popcount33_95r9_core_209 = input_a[15] | input_a[15];
  assign popcount33_95r9_core_210 = input_a[23] ^ input_a[2];
  assign popcount33_95r9_core_214 = ~(input_a[25] & input_a[2]);
  assign popcount33_95r9_core_215 = ~input_a[6];
  assign popcount33_95r9_core_216 = ~input_a[32];
  assign popcount33_95r9_core_218 = ~(input_a[3] & input_a[22]);
  assign popcount33_95r9_core_219 = input_a[32] ^ input_a[25];
  assign popcount33_95r9_core_222 = ~(input_a[19] | input_a[12]);
  assign popcount33_95r9_core_223 = input_a[0] ^ input_a[11];
  assign popcount33_95r9_core_225 = ~(input_a[15] ^ input_a[23]);
  assign popcount33_95r9_core_227 = input_a[15] | input_a[14];
  assign popcount33_95r9_core_228 = input_a[6] ^ input_a[10];
  assign popcount33_95r9_core_232 = ~(input_a[15] | input_a[0]);
  assign popcount33_95r9_core_233 = ~(input_a[13] & input_a[14]);
  assign popcount33_95r9_core_234 = input_a[11] & input_a[14];
  assign popcount33_95r9_core_236 = input_a[24] ^ input_a[32];
  assign popcount33_95r9_core_238 = ~(input_a[0] | input_a[23]);

  assign popcount33_95r9_out[0] = 1'b0;
  assign popcount33_95r9_out[1] = input_a[13];
  assign popcount33_95r9_out[2] = 1'b1;
  assign popcount33_95r9_out[3] = input_a[6];
  assign popcount33_95r9_out[4] = input_a[19];
  assign popcount33_95r9_out[5] = 1'b0;
endmodule