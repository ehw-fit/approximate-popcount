// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5285
// WCE=43.0
// EP=0.992257%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_q8j1(input [33:0] input_a, output [5:0] popcount34_q8j1_out);
  wire popcount34_q8j1_core_037;
  wire popcount34_q8j1_core_038;
  wire popcount34_q8j1_core_039;
  wire popcount34_q8j1_core_040;
  wire popcount34_q8j1_core_041;
  wire popcount34_q8j1_core_042;
  wire popcount34_q8j1_core_043;
  wire popcount34_q8j1_core_044;
  wire popcount34_q8j1_core_045;
  wire popcount34_q8j1_core_046;
  wire popcount34_q8j1_core_047;
  wire popcount34_q8j1_core_049;
  wire popcount34_q8j1_core_050;
  wire popcount34_q8j1_core_051;
  wire popcount34_q8j1_core_052;
  wire popcount34_q8j1_core_053;
  wire popcount34_q8j1_core_056;
  wire popcount34_q8j1_core_058;
  wire popcount34_q8j1_core_060;
  wire popcount34_q8j1_core_061;
  wire popcount34_q8j1_core_063;
  wire popcount34_q8j1_core_064;
  wire popcount34_q8j1_core_065;
  wire popcount34_q8j1_core_066;
  wire popcount34_q8j1_core_067;
  wire popcount34_q8j1_core_069;
  wire popcount34_q8j1_core_070;
  wire popcount34_q8j1_core_071;
  wire popcount34_q8j1_core_072;
  wire popcount34_q8j1_core_073;
  wire popcount34_q8j1_core_075;
  wire popcount34_q8j1_core_076;
  wire popcount34_q8j1_core_077;
  wire popcount34_q8j1_core_080;
  wire popcount34_q8j1_core_082;
  wire popcount34_q8j1_core_083;
  wire popcount34_q8j1_core_084;
  wire popcount34_q8j1_core_086;
  wire popcount34_q8j1_core_088;
  wire popcount34_q8j1_core_090;
  wire popcount34_q8j1_core_091;
  wire popcount34_q8j1_core_093;
  wire popcount34_q8j1_core_095;
  wire popcount34_q8j1_core_096;
  wire popcount34_q8j1_core_098;
  wire popcount34_q8j1_core_099;
  wire popcount34_q8j1_core_100;
  wire popcount34_q8j1_core_101;
  wire popcount34_q8j1_core_102;
  wire popcount34_q8j1_core_104;
  wire popcount34_q8j1_core_106;
  wire popcount34_q8j1_core_107;
  wire popcount34_q8j1_core_108;
  wire popcount34_q8j1_core_110;
  wire popcount34_q8j1_core_112;
  wire popcount34_q8j1_core_114;
  wire popcount34_q8j1_core_115;
  wire popcount34_q8j1_core_116;
  wire popcount34_q8j1_core_119;
  wire popcount34_q8j1_core_120;
  wire popcount34_q8j1_core_121;
  wire popcount34_q8j1_core_122;
  wire popcount34_q8j1_core_123;
  wire popcount34_q8j1_core_124;
  wire popcount34_q8j1_core_125;
  wire popcount34_q8j1_core_126;
  wire popcount34_q8j1_core_127;
  wire popcount34_q8j1_core_128;
  wire popcount34_q8j1_core_129;
  wire popcount34_q8j1_core_130;
  wire popcount34_q8j1_core_132;
  wire popcount34_q8j1_core_133;
  wire popcount34_q8j1_core_138;
  wire popcount34_q8j1_core_141;
  wire popcount34_q8j1_core_142;
  wire popcount34_q8j1_core_144;
  wire popcount34_q8j1_core_145;
  wire popcount34_q8j1_core_147;
  wire popcount34_q8j1_core_148;
  wire popcount34_q8j1_core_152;
  wire popcount34_q8j1_core_153;
  wire popcount34_q8j1_core_156;
  wire popcount34_q8j1_core_157_not;
  wire popcount34_q8j1_core_159;
  wire popcount34_q8j1_core_160;
  wire popcount34_q8j1_core_161;
  wire popcount34_q8j1_core_162;
  wire popcount34_q8j1_core_163;
  wire popcount34_q8j1_core_164_not;
  wire popcount34_q8j1_core_165_not;
  wire popcount34_q8j1_core_166;
  wire popcount34_q8j1_core_167;
  wire popcount34_q8j1_core_168;
  wire popcount34_q8j1_core_175;
  wire popcount34_q8j1_core_177;
  wire popcount34_q8j1_core_178;
  wire popcount34_q8j1_core_179;
  wire popcount34_q8j1_core_180;
  wire popcount34_q8j1_core_181;
  wire popcount34_q8j1_core_183;
  wire popcount34_q8j1_core_184;
  wire popcount34_q8j1_core_186;
  wire popcount34_q8j1_core_187;
  wire popcount34_q8j1_core_188;
  wire popcount34_q8j1_core_190;
  wire popcount34_q8j1_core_191;
  wire popcount34_q8j1_core_192;
  wire popcount34_q8j1_core_193;
  wire popcount34_q8j1_core_194;
  wire popcount34_q8j1_core_195;
  wire popcount34_q8j1_core_196;
  wire popcount34_q8j1_core_197;
  wire popcount34_q8j1_core_198;
  wire popcount34_q8j1_core_199;
  wire popcount34_q8j1_core_201;
  wire popcount34_q8j1_core_202;
  wire popcount34_q8j1_core_206;
  wire popcount34_q8j1_core_208;
  wire popcount34_q8j1_core_209;
  wire popcount34_q8j1_core_210;
  wire popcount34_q8j1_core_211;
  wire popcount34_q8j1_core_212;
  wire popcount34_q8j1_core_214;
  wire popcount34_q8j1_core_215;
  wire popcount34_q8j1_core_216;
  wire popcount34_q8j1_core_219;
  wire popcount34_q8j1_core_220;
  wire popcount34_q8j1_core_221;
  wire popcount34_q8j1_core_225;
  wire popcount34_q8j1_core_226;
  wire popcount34_q8j1_core_228;
  wire popcount34_q8j1_core_229;
  wire popcount34_q8j1_core_230;
  wire popcount34_q8j1_core_231;
  wire popcount34_q8j1_core_233;
  wire popcount34_q8j1_core_234;
  wire popcount34_q8j1_core_235;
  wire popcount34_q8j1_core_236;
  wire popcount34_q8j1_core_239;
  wire popcount34_q8j1_core_240_not;
  wire popcount34_q8j1_core_241_not;
  wire popcount34_q8j1_core_243;
  wire popcount34_q8j1_core_244;
  wire popcount34_q8j1_core_245;
  wire popcount34_q8j1_core_246;
  wire popcount34_q8j1_core_247;
  wire popcount34_q8j1_core_248;
  wire popcount34_q8j1_core_250;
  wire popcount34_q8j1_core_251;

  assign popcount34_q8j1_core_037 = ~(input_a[9] | input_a[5]);
  assign popcount34_q8j1_core_038 = input_a[26] ^ input_a[28];
  assign popcount34_q8j1_core_039 = ~(input_a[27] | input_a[16]);
  assign popcount34_q8j1_core_040 = ~(input_a[31] & input_a[21]);
  assign popcount34_q8j1_core_041 = ~(input_a[29] ^ input_a[27]);
  assign popcount34_q8j1_core_042 = ~(input_a[12] ^ input_a[3]);
  assign popcount34_q8j1_core_043 = ~(input_a[0] | input_a[30]);
  assign popcount34_q8j1_core_044 = input_a[21] ^ input_a[0];
  assign popcount34_q8j1_core_045 = ~(input_a[8] ^ input_a[25]);
  assign popcount34_q8j1_core_046 = ~(input_a[3] ^ input_a[33]);
  assign popcount34_q8j1_core_047 = input_a[6] ^ input_a[5];
  assign popcount34_q8j1_core_049 = input_a[25] | input_a[12];
  assign popcount34_q8j1_core_050 = ~(input_a[4] & input_a[17]);
  assign popcount34_q8j1_core_051 = input_a[20] | input_a[31];
  assign popcount34_q8j1_core_052 = ~(input_a[30] | input_a[15]);
  assign popcount34_q8j1_core_053 = ~(input_a[22] | input_a[29]);
  assign popcount34_q8j1_core_056 = ~(input_a[16] | input_a[16]);
  assign popcount34_q8j1_core_058 = input_a[3] ^ input_a[5];
  assign popcount34_q8j1_core_060 = input_a[31] & input_a[26];
  assign popcount34_q8j1_core_061 = ~(input_a[28] & input_a[24]);
  assign popcount34_q8j1_core_063 = ~(input_a[1] | input_a[8]);
  assign popcount34_q8j1_core_064 = ~(input_a[3] & input_a[28]);
  assign popcount34_q8j1_core_065 = input_a[33] | input_a[25];
  assign popcount34_q8j1_core_066 = input_a[11] ^ input_a[31];
  assign popcount34_q8j1_core_067 = input_a[22] | input_a[30];
  assign popcount34_q8j1_core_069 = ~(input_a[9] ^ input_a[30]);
  assign popcount34_q8j1_core_070 = ~input_a[32];
  assign popcount34_q8j1_core_071 = ~(input_a[17] & input_a[22]);
  assign popcount34_q8j1_core_072 = ~(input_a[16] & input_a[6]);
  assign popcount34_q8j1_core_073 = ~(input_a[15] ^ input_a[33]);
  assign popcount34_q8j1_core_075 = input_a[13] ^ input_a[26];
  assign popcount34_q8j1_core_076 = ~(input_a[12] | input_a[25]);
  assign popcount34_q8j1_core_077 = ~(input_a[28] | input_a[2]);
  assign popcount34_q8j1_core_080 = ~(input_a[7] & input_a[18]);
  assign popcount34_q8j1_core_082 = ~(input_a[11] | input_a[11]);
  assign popcount34_q8j1_core_083 = input_a[15] ^ input_a[12];
  assign popcount34_q8j1_core_084 = ~(input_a[12] & input_a[0]);
  assign popcount34_q8j1_core_086 = input_a[16] | input_a[28];
  assign popcount34_q8j1_core_088 = input_a[19] & input_a[3];
  assign popcount34_q8j1_core_090 = input_a[9] ^ input_a[2];
  assign popcount34_q8j1_core_091 = input_a[22] & input_a[24];
  assign popcount34_q8j1_core_093 = input_a[31] ^ input_a[25];
  assign popcount34_q8j1_core_095 = ~input_a[22];
  assign popcount34_q8j1_core_096 = input_a[31] & input_a[23];
  assign popcount34_q8j1_core_098 = ~input_a[33];
  assign popcount34_q8j1_core_099 = ~(input_a[24] ^ input_a[6]);
  assign popcount34_q8j1_core_100 = ~(input_a[1] & input_a[16]);
  assign popcount34_q8j1_core_101 = ~(input_a[5] & input_a[18]);
  assign popcount34_q8j1_core_102 = ~(input_a[17] | input_a[7]);
  assign popcount34_q8j1_core_104 = ~(input_a[19] & input_a[24]);
  assign popcount34_q8j1_core_106 = ~input_a[3];
  assign popcount34_q8j1_core_107 = input_a[28] | input_a[12];
  assign popcount34_q8j1_core_108 = ~(input_a[0] | input_a[0]);
  assign popcount34_q8j1_core_110 = ~(input_a[19] & input_a[23]);
  assign popcount34_q8j1_core_112 = ~(input_a[8] ^ input_a[6]);
  assign popcount34_q8j1_core_114 = ~(input_a[0] & input_a[19]);
  assign popcount34_q8j1_core_115 = ~(input_a[17] | input_a[23]);
  assign popcount34_q8j1_core_116 = ~(input_a[8] & input_a[12]);
  assign popcount34_q8j1_core_119 = ~(input_a[13] & input_a[14]);
  assign popcount34_q8j1_core_120 = ~(input_a[31] & input_a[6]);
  assign popcount34_q8j1_core_121 = input_a[25] ^ input_a[24];
  assign popcount34_q8j1_core_122 = input_a[30] | input_a[19];
  assign popcount34_q8j1_core_123 = ~(input_a[4] ^ input_a[14]);
  assign popcount34_q8j1_core_124 = input_a[9] ^ input_a[10];
  assign popcount34_q8j1_core_125 = input_a[26] ^ input_a[20];
  assign popcount34_q8j1_core_126 = input_a[11] & input_a[30];
  assign popcount34_q8j1_core_127 = input_a[23] | input_a[33];
  assign popcount34_q8j1_core_128 = ~(input_a[3] & input_a[10]);
  assign popcount34_q8j1_core_129 = ~input_a[28];
  assign popcount34_q8j1_core_130 = ~(input_a[3] ^ input_a[16]);
  assign popcount34_q8j1_core_132 = input_a[8] | input_a[23];
  assign popcount34_q8j1_core_133 = ~(input_a[6] & input_a[18]);
  assign popcount34_q8j1_core_138 = ~(input_a[32] ^ input_a[13]);
  assign popcount34_q8j1_core_141 = ~(input_a[28] & input_a[33]);
  assign popcount34_q8j1_core_142 = ~(input_a[3] | input_a[20]);
  assign popcount34_q8j1_core_144 = input_a[22] | input_a[11];
  assign popcount34_q8j1_core_145 = ~input_a[28];
  assign popcount34_q8j1_core_147 = input_a[21] ^ input_a[26];
  assign popcount34_q8j1_core_148 = input_a[17] & input_a[25];
  assign popcount34_q8j1_core_152 = input_a[6] ^ input_a[3];
  assign popcount34_q8j1_core_153 = ~input_a[5];
  assign popcount34_q8j1_core_156 = input_a[0] & input_a[17];
  assign popcount34_q8j1_core_157_not = ~input_a[27];
  assign popcount34_q8j1_core_159 = ~(input_a[25] | input_a[31]);
  assign popcount34_q8j1_core_160 = input_a[11] ^ input_a[22];
  assign popcount34_q8j1_core_161 = input_a[23] ^ input_a[2];
  assign popcount34_q8j1_core_162 = ~(input_a[33] & input_a[1]);
  assign popcount34_q8j1_core_163 = input_a[14] ^ input_a[23];
  assign popcount34_q8j1_core_164_not = ~input_a[11];
  assign popcount34_q8j1_core_165_not = ~input_a[24];
  assign popcount34_q8j1_core_166 = ~(input_a[5] ^ input_a[28]);
  assign popcount34_q8j1_core_167 = ~input_a[25];
  assign popcount34_q8j1_core_168 = input_a[13] | input_a[0];
  assign popcount34_q8j1_core_175 = ~(input_a[11] & input_a[28]);
  assign popcount34_q8j1_core_177 = ~(input_a[9] ^ input_a[19]);
  assign popcount34_q8j1_core_178 = input_a[5] | input_a[29];
  assign popcount34_q8j1_core_179 = input_a[33] | input_a[10];
  assign popcount34_q8j1_core_180 = ~(input_a[33] & input_a[25]);
  assign popcount34_q8j1_core_181 = ~(input_a[18] & input_a[18]);
  assign popcount34_q8j1_core_183 = input_a[7] ^ input_a[5];
  assign popcount34_q8j1_core_184 = ~(input_a[24] | input_a[19]);
  assign popcount34_q8j1_core_186 = input_a[27] ^ input_a[24];
  assign popcount34_q8j1_core_187 = ~input_a[33];
  assign popcount34_q8j1_core_188 = ~input_a[2];
  assign popcount34_q8j1_core_190 = ~(input_a[15] | input_a[19]);
  assign popcount34_q8j1_core_191 = ~(input_a[30] ^ input_a[24]);
  assign popcount34_q8j1_core_192 = ~input_a[28];
  assign popcount34_q8j1_core_193 = ~(input_a[32] | input_a[13]);
  assign popcount34_q8j1_core_194 = ~(input_a[16] & input_a[16]);
  assign popcount34_q8j1_core_195 = ~input_a[2];
  assign popcount34_q8j1_core_196 = input_a[26] | input_a[6];
  assign popcount34_q8j1_core_197 = ~(input_a[14] | input_a[10]);
  assign popcount34_q8j1_core_198 = ~input_a[29];
  assign popcount34_q8j1_core_199 = ~(input_a[21] & input_a[20]);
  assign popcount34_q8j1_core_201 = ~input_a[12];
  assign popcount34_q8j1_core_202 = input_a[19] ^ input_a[16];
  assign popcount34_q8j1_core_206 = input_a[15] ^ input_a[31];
  assign popcount34_q8j1_core_208 = ~(input_a[29] | input_a[21]);
  assign popcount34_q8j1_core_209 = input_a[20] | input_a[1];
  assign popcount34_q8j1_core_210 = input_a[13] & input_a[28];
  assign popcount34_q8j1_core_211 = input_a[19] | input_a[7];
  assign popcount34_q8j1_core_212 = input_a[9] ^ input_a[27];
  assign popcount34_q8j1_core_214 = ~input_a[23];
  assign popcount34_q8j1_core_215 = ~input_a[28];
  assign popcount34_q8j1_core_216 = input_a[13] | input_a[14];
  assign popcount34_q8j1_core_219 = ~(input_a[23] ^ input_a[25]);
  assign popcount34_q8j1_core_220 = ~(input_a[17] ^ input_a[14]);
  assign popcount34_q8j1_core_221 = ~input_a[25];
  assign popcount34_q8j1_core_225 = ~(input_a[16] | input_a[17]);
  assign popcount34_q8j1_core_226 = input_a[3] | input_a[19];
  assign popcount34_q8j1_core_228 = ~(input_a[12] | input_a[29]);
  assign popcount34_q8j1_core_229 = input_a[25] ^ input_a[3];
  assign popcount34_q8j1_core_230 = input_a[6] ^ input_a[4];
  assign popcount34_q8j1_core_231 = ~(input_a[8] & input_a[20]);
  assign popcount34_q8j1_core_233 = ~(input_a[12] ^ input_a[33]);
  assign popcount34_q8j1_core_234 = ~(input_a[16] & input_a[22]);
  assign popcount34_q8j1_core_235 = input_a[23] ^ input_a[25];
  assign popcount34_q8j1_core_236 = ~(input_a[23] & input_a[20]);
  assign popcount34_q8j1_core_239 = ~(input_a[17] ^ input_a[1]);
  assign popcount34_q8j1_core_240_not = ~input_a[20];
  assign popcount34_q8j1_core_241_not = ~input_a[2];
  assign popcount34_q8j1_core_243 = ~(input_a[28] | input_a[23]);
  assign popcount34_q8j1_core_244 = input_a[31] & input_a[21];
  assign popcount34_q8j1_core_245 = input_a[29] & input_a[30];
  assign popcount34_q8j1_core_246 = ~(input_a[13] & input_a[33]);
  assign popcount34_q8j1_core_247 = input_a[31] ^ input_a[21];
  assign popcount34_q8j1_core_248 = input_a[15] ^ input_a[4];
  assign popcount34_q8j1_core_250 = ~(input_a[28] & input_a[16]);
  assign popcount34_q8j1_core_251 = ~input_a[10];

  assign popcount34_q8j1_out[0] = input_a[1];
  assign popcount34_q8j1_out[1] = 1'b0;
  assign popcount34_q8j1_out[2] = input_a[11];
  assign popcount34_q8j1_out[3] = input_a[3];
  assign popcount34_q8j1_out[4] = 1'b0;
  assign popcount34_q8j1_out[5] = input_a[22];
endmodule