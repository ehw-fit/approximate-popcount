// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.24169
// WCE=15.0
// EP=0.860517%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_pk69(input [27:0] input_a, output [4:0] popcount28_pk69_out);
  wire popcount28_pk69_core_030;
  wire popcount28_pk69_core_031;
  wire popcount28_pk69_core_032;
  wire popcount28_pk69_core_033;
  wire popcount28_pk69_core_035;
  wire popcount28_pk69_core_037;
  wire popcount28_pk69_core_039;
  wire popcount28_pk69_core_040;
  wire popcount28_pk69_core_042;
  wire popcount28_pk69_core_044;
  wire popcount28_pk69_core_049;
  wire popcount28_pk69_core_051;
  wire popcount28_pk69_core_054;
  wire popcount28_pk69_core_055;
  wire popcount28_pk69_core_057;
  wire popcount28_pk69_core_058;
  wire popcount28_pk69_core_059;
  wire popcount28_pk69_core_063;
  wire popcount28_pk69_core_065;
  wire popcount28_pk69_core_068;
  wire popcount28_pk69_core_069;
  wire popcount28_pk69_core_071;
  wire popcount28_pk69_core_072;
  wire popcount28_pk69_core_073;
  wire popcount28_pk69_core_074;
  wire popcount28_pk69_core_077_not;
  wire popcount28_pk69_core_078;
  wire popcount28_pk69_core_079;
  wire popcount28_pk69_core_081;
  wire popcount28_pk69_core_083;
  wire popcount28_pk69_core_084;
  wire popcount28_pk69_core_086;
  wire popcount28_pk69_core_088;
  wire popcount28_pk69_core_089;
  wire popcount28_pk69_core_090;
  wire popcount28_pk69_core_092;
  wire popcount28_pk69_core_093;
  wire popcount28_pk69_core_094;
  wire popcount28_pk69_core_095;
  wire popcount28_pk69_core_097;
  wire popcount28_pk69_core_098;
  wire popcount28_pk69_core_099;
  wire popcount28_pk69_core_100;
  wire popcount28_pk69_core_102;
  wire popcount28_pk69_core_104;
  wire popcount28_pk69_core_105;
  wire popcount28_pk69_core_106;
  wire popcount28_pk69_core_107;
  wire popcount28_pk69_core_109;
  wire popcount28_pk69_core_111;
  wire popcount28_pk69_core_112;
  wire popcount28_pk69_core_113;
  wire popcount28_pk69_core_114;
  wire popcount28_pk69_core_116;
  wire popcount28_pk69_core_117;
  wire popcount28_pk69_core_118;
  wire popcount28_pk69_core_119;
  wire popcount28_pk69_core_126;
  wire popcount28_pk69_core_128;
  wire popcount28_pk69_core_129;
  wire popcount28_pk69_core_130;
  wire popcount28_pk69_core_131;
  wire popcount28_pk69_core_132;
  wire popcount28_pk69_core_134_not;
  wire popcount28_pk69_core_135;
  wire popcount28_pk69_core_136;
  wire popcount28_pk69_core_138;
  wire popcount28_pk69_core_139;
  wire popcount28_pk69_core_140;
  wire popcount28_pk69_core_142;
  wire popcount28_pk69_core_144;
  wire popcount28_pk69_core_145;
  wire popcount28_pk69_core_146;
  wire popcount28_pk69_core_147_not;
  wire popcount28_pk69_core_149;
  wire popcount28_pk69_core_152;
  wire popcount28_pk69_core_153;
  wire popcount28_pk69_core_154;
  wire popcount28_pk69_core_155;
  wire popcount28_pk69_core_157;
  wire popcount28_pk69_core_159;
  wire popcount28_pk69_core_160;
  wire popcount28_pk69_core_161;
  wire popcount28_pk69_core_162;
  wire popcount28_pk69_core_163;
  wire popcount28_pk69_core_164;
  wire popcount28_pk69_core_165;
  wire popcount28_pk69_core_169;
  wire popcount28_pk69_core_171;
  wire popcount28_pk69_core_172;
  wire popcount28_pk69_core_176;
  wire popcount28_pk69_core_179;
  wire popcount28_pk69_core_181;
  wire popcount28_pk69_core_182_not;
  wire popcount28_pk69_core_183;
  wire popcount28_pk69_core_185;
  wire popcount28_pk69_core_186;
  wire popcount28_pk69_core_188;
  wire popcount28_pk69_core_194;
  wire popcount28_pk69_core_196;
  wire popcount28_pk69_core_197;
  wire popcount28_pk69_core_198;
  wire popcount28_pk69_core_200;
  wire popcount28_pk69_core_201;

  assign popcount28_pk69_core_030 = input_a[20] | input_a[4];
  assign popcount28_pk69_core_031 = input_a[14] | input_a[21];
  assign popcount28_pk69_core_032 = input_a[13] | input_a[21];
  assign popcount28_pk69_core_033 = ~(input_a[0] & input_a[8]);
  assign popcount28_pk69_core_035 = ~(input_a[13] & input_a[23]);
  assign popcount28_pk69_core_037 = ~input_a[25];
  assign popcount28_pk69_core_039 = ~(input_a[5] | input_a[13]);
  assign popcount28_pk69_core_040 = input_a[25] & input_a[21];
  assign popcount28_pk69_core_042 = ~(input_a[4] | input_a[24]);
  assign popcount28_pk69_core_044 = ~(input_a[1] & input_a[27]);
  assign popcount28_pk69_core_049 = ~input_a[3];
  assign popcount28_pk69_core_051 = input_a[18] | input_a[27];
  assign popcount28_pk69_core_054 = ~(input_a[25] | input_a[6]);
  assign popcount28_pk69_core_055 = input_a[18] | input_a[24];
  assign popcount28_pk69_core_057 = ~(input_a[17] ^ input_a[1]);
  assign popcount28_pk69_core_058 = input_a[16] | input_a[27];
  assign popcount28_pk69_core_059 = ~(input_a[13] | input_a[9]);
  assign popcount28_pk69_core_063 = ~(input_a[21] & input_a[21]);
  assign popcount28_pk69_core_065 = input_a[15] ^ input_a[4];
  assign popcount28_pk69_core_068 = ~(input_a[25] ^ input_a[27]);
  assign popcount28_pk69_core_069 = input_a[7] & input_a[21];
  assign popcount28_pk69_core_071 = ~(input_a[25] ^ input_a[26]);
  assign popcount28_pk69_core_072 = ~(input_a[2] ^ input_a[5]);
  assign popcount28_pk69_core_073 = input_a[26] | input_a[23];
  assign popcount28_pk69_core_074 = ~(input_a[18] | input_a[9]);
  assign popcount28_pk69_core_077_not = ~input_a[18];
  assign popcount28_pk69_core_078 = ~(input_a[16] & input_a[14]);
  assign popcount28_pk69_core_079 = input_a[26] ^ input_a[23];
  assign popcount28_pk69_core_081 = ~(input_a[2] ^ input_a[12]);
  assign popcount28_pk69_core_083 = ~(input_a[2] | input_a[19]);
  assign popcount28_pk69_core_084 = ~input_a[11];
  assign popcount28_pk69_core_086 = ~(input_a[19] | input_a[15]);
  assign popcount28_pk69_core_088 = input_a[3] & input_a[13];
  assign popcount28_pk69_core_089 = input_a[2] & input_a[9];
  assign popcount28_pk69_core_090 = ~(input_a[6] & input_a[22]);
  assign popcount28_pk69_core_092 = input_a[25] ^ input_a[10];
  assign popcount28_pk69_core_093 = ~(input_a[12] ^ input_a[3]);
  assign popcount28_pk69_core_094 = ~(input_a[4] ^ input_a[18]);
  assign popcount28_pk69_core_095 = ~(input_a[14] | input_a[17]);
  assign popcount28_pk69_core_097 = ~(input_a[24] & input_a[14]);
  assign popcount28_pk69_core_098 = input_a[23] & input_a[27];
  assign popcount28_pk69_core_099 = input_a[7] & input_a[17];
  assign popcount28_pk69_core_100 = ~(input_a[23] & input_a[27]);
  assign popcount28_pk69_core_102 = ~(input_a[5] & input_a[19]);
  assign popcount28_pk69_core_104 = ~(input_a[19] ^ input_a[18]);
  assign popcount28_pk69_core_105 = ~(input_a[3] ^ input_a[1]);
  assign popcount28_pk69_core_106 = input_a[9] & input_a[27];
  assign popcount28_pk69_core_107 = input_a[6] ^ input_a[14];
  assign popcount28_pk69_core_109 = input_a[7] ^ input_a[2];
  assign popcount28_pk69_core_111 = ~(input_a[22] & input_a[27]);
  assign popcount28_pk69_core_112 = ~(input_a[8] & input_a[26]);
  assign popcount28_pk69_core_113 = input_a[12] & input_a[24];
  assign popcount28_pk69_core_114 = ~input_a[12];
  assign popcount28_pk69_core_116 = input_a[4] ^ input_a[20];
  assign popcount28_pk69_core_117 = ~(input_a[1] | input_a[20]);
  assign popcount28_pk69_core_118 = input_a[10] | input_a[5];
  assign popcount28_pk69_core_119 = ~(input_a[23] & input_a[11]);
  assign popcount28_pk69_core_126 = ~(input_a[10] | input_a[1]);
  assign popcount28_pk69_core_128 = input_a[7] ^ input_a[7];
  assign popcount28_pk69_core_129 = input_a[26] ^ input_a[8];
  assign popcount28_pk69_core_130 = input_a[3] ^ input_a[23];
  assign popcount28_pk69_core_131 = input_a[9] ^ input_a[26];
  assign popcount28_pk69_core_132 = input_a[8] ^ input_a[17];
  assign popcount28_pk69_core_134_not = ~input_a[15];
  assign popcount28_pk69_core_135 = input_a[27] | input_a[5];
  assign popcount28_pk69_core_136 = input_a[9] | input_a[21];
  assign popcount28_pk69_core_138 = ~input_a[8];
  assign popcount28_pk69_core_139 = ~(input_a[5] & input_a[11]);
  assign popcount28_pk69_core_140 = ~(input_a[13] | input_a[11]);
  assign popcount28_pk69_core_142 = input_a[20] | input_a[5];
  assign popcount28_pk69_core_144 = ~(input_a[6] ^ input_a[20]);
  assign popcount28_pk69_core_145 = ~input_a[10];
  assign popcount28_pk69_core_146 = input_a[25] ^ input_a[0];
  assign popcount28_pk69_core_147_not = ~input_a[5];
  assign popcount28_pk69_core_149 = ~(input_a[17] ^ input_a[4]);
  assign popcount28_pk69_core_152 = input_a[3] ^ input_a[17];
  assign popcount28_pk69_core_153 = input_a[18] & input_a[9];
  assign popcount28_pk69_core_154 = ~(input_a[20] & input_a[19]);
  assign popcount28_pk69_core_155 = ~(input_a[10] ^ input_a[6]);
  assign popcount28_pk69_core_157 = ~input_a[7];
  assign popcount28_pk69_core_159 = input_a[20] ^ input_a[8];
  assign popcount28_pk69_core_160 = ~input_a[3];
  assign popcount28_pk69_core_161 = input_a[15] & input_a[19];
  assign popcount28_pk69_core_162 = input_a[14] | input_a[16];
  assign popcount28_pk69_core_163 = ~(input_a[10] | input_a[16]);
  assign popcount28_pk69_core_164 = input_a[3] ^ input_a[16];
  assign popcount28_pk69_core_165 = ~(input_a[7] | input_a[14]);
  assign popcount28_pk69_core_169 = ~(input_a[14] | input_a[27]);
  assign popcount28_pk69_core_171 = input_a[5] ^ input_a[14];
  assign popcount28_pk69_core_172 = ~input_a[10];
  assign popcount28_pk69_core_176 = input_a[11] & input_a[14];
  assign popcount28_pk69_core_179 = ~(input_a[15] & input_a[22]);
  assign popcount28_pk69_core_181 = input_a[13] ^ input_a[26];
  assign popcount28_pk69_core_182_not = ~input_a[26];
  assign popcount28_pk69_core_183 = ~input_a[24];
  assign popcount28_pk69_core_185 = ~input_a[10];
  assign popcount28_pk69_core_186 = ~(input_a[19] & input_a[11]);
  assign popcount28_pk69_core_188 = input_a[13] | input_a[19];
  assign popcount28_pk69_core_194 = input_a[2] ^ input_a[0];
  assign popcount28_pk69_core_196 = input_a[3] | input_a[8];
  assign popcount28_pk69_core_197 = input_a[15] | input_a[12];
  assign popcount28_pk69_core_198 = input_a[16] | input_a[5];
  assign popcount28_pk69_core_200 = input_a[26] ^ input_a[18];
  assign popcount28_pk69_core_201 = input_a[8] ^ input_a[1];

  assign popcount28_pk69_out[0] = 1'b1;
  assign popcount28_pk69_out[1] = 1'b1;
  assign popcount28_pk69_out[2] = 1'b1;
  assign popcount28_pk69_out[3] = 1'b1;
  assign popcount28_pk69_out[4] = 1'b0;
endmodule