// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.93817
// WCE=11.0
// EP=0.839821%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_mjel(input [20:0] input_a, output [4:0] popcount21_mjel_out);
  wire popcount21_mjel_core_023;
  wire popcount21_mjel_core_026;
  wire popcount21_mjel_core_030;
  wire popcount21_mjel_core_032;
  wire popcount21_mjel_core_033;
  wire popcount21_mjel_core_034;
  wire popcount21_mjel_core_035;
  wire popcount21_mjel_core_036;
  wire popcount21_mjel_core_038;
  wire popcount21_mjel_core_042;
  wire popcount21_mjel_core_043;
  wire popcount21_mjel_core_044;
  wire popcount21_mjel_core_045;
  wire popcount21_mjel_core_046;
  wire popcount21_mjel_core_049;
  wire popcount21_mjel_core_053;
  wire popcount21_mjel_core_055;
  wire popcount21_mjel_core_056;
  wire popcount21_mjel_core_058;
  wire popcount21_mjel_core_059;
  wire popcount21_mjel_core_060;
  wire popcount21_mjel_core_061;
  wire popcount21_mjel_core_063;
  wire popcount21_mjel_core_066;
  wire popcount21_mjel_core_067;
  wire popcount21_mjel_core_068;
  wire popcount21_mjel_core_069;
  wire popcount21_mjel_core_070;
  wire popcount21_mjel_core_073;
  wire popcount21_mjel_core_074;
  wire popcount21_mjel_core_075;
  wire popcount21_mjel_core_077;
  wire popcount21_mjel_core_078_not;
  wire popcount21_mjel_core_079;
  wire popcount21_mjel_core_081;
  wire popcount21_mjel_core_082;
  wire popcount21_mjel_core_085;
  wire popcount21_mjel_core_086;
  wire popcount21_mjel_core_089;
  wire popcount21_mjel_core_091;
  wire popcount21_mjel_core_095;
  wire popcount21_mjel_core_098;
  wire popcount21_mjel_core_099;
  wire popcount21_mjel_core_100;
  wire popcount21_mjel_core_101;
  wire popcount21_mjel_core_103;
  wire popcount21_mjel_core_104;
  wire popcount21_mjel_core_105_not;
  wire popcount21_mjel_core_108;
  wire popcount21_mjel_core_112;
  wire popcount21_mjel_core_114;
  wire popcount21_mjel_core_116;
  wire popcount21_mjel_core_117;
  wire popcount21_mjel_core_120;
  wire popcount21_mjel_core_122;
  wire popcount21_mjel_core_124;
  wire popcount21_mjel_core_125;
  wire popcount21_mjel_core_133;
  wire popcount21_mjel_core_134;
  wire popcount21_mjel_core_135;
  wire popcount21_mjel_core_137_not;
  wire popcount21_mjel_core_138;
  wire popcount21_mjel_core_139;
  wire popcount21_mjel_core_140;
  wire popcount21_mjel_core_141;
  wire popcount21_mjel_core_142;
  wire popcount21_mjel_core_144;
  wire popcount21_mjel_core_147;
  wire popcount21_mjel_core_148;
  wire popcount21_mjel_core_150;
  wire popcount21_mjel_core_151;
  wire popcount21_mjel_core_153;

  assign popcount21_mjel_core_023 = ~(input_a[18] & input_a[13]);
  assign popcount21_mjel_core_026 = ~(input_a[11] | input_a[9]);
  assign popcount21_mjel_core_030 = input_a[13] | input_a[1];
  assign popcount21_mjel_core_032 = input_a[20] ^ input_a[20];
  assign popcount21_mjel_core_033 = input_a[14] ^ input_a[9];
  assign popcount21_mjel_core_034 = input_a[0] | input_a[3];
  assign popcount21_mjel_core_035 = ~(input_a[17] ^ input_a[4]);
  assign popcount21_mjel_core_036 = ~(input_a[6] ^ input_a[10]);
  assign popcount21_mjel_core_038 = ~(input_a[8] ^ input_a[0]);
  assign popcount21_mjel_core_042 = ~(input_a[6] ^ input_a[6]);
  assign popcount21_mjel_core_043 = ~input_a[0];
  assign popcount21_mjel_core_044 = ~(input_a[15] | input_a[5]);
  assign popcount21_mjel_core_045 = input_a[7] | input_a[9];
  assign popcount21_mjel_core_046 = ~(input_a[9] ^ input_a[6]);
  assign popcount21_mjel_core_049 = input_a[1] | input_a[10];
  assign popcount21_mjel_core_053 = ~(input_a[6] | input_a[7]);
  assign popcount21_mjel_core_055 = ~(input_a[13] | input_a[1]);
  assign popcount21_mjel_core_056 = ~(input_a[7] ^ input_a[1]);
  assign popcount21_mjel_core_058 = ~(input_a[14] ^ input_a[2]);
  assign popcount21_mjel_core_059 = ~input_a[1];
  assign popcount21_mjel_core_060 = input_a[13] | input_a[4];
  assign popcount21_mjel_core_061 = ~(input_a[3] & input_a[15]);
  assign popcount21_mjel_core_063 = ~input_a[10];
  assign popcount21_mjel_core_066 = input_a[16] | input_a[7];
  assign popcount21_mjel_core_067 = input_a[8] & input_a[16];
  assign popcount21_mjel_core_068 = input_a[9] ^ input_a[16];
  assign popcount21_mjel_core_069 = ~(input_a[4] & input_a[3]);
  assign popcount21_mjel_core_070 = input_a[10] & input_a[15];
  assign popcount21_mjel_core_073 = ~input_a[3];
  assign popcount21_mjel_core_074 = input_a[14] & input_a[9];
  assign popcount21_mjel_core_075 = input_a[20] & input_a[1];
  assign popcount21_mjel_core_077 = ~input_a[18];
  assign popcount21_mjel_core_078_not = ~input_a[16];
  assign popcount21_mjel_core_079 = ~(input_a[14] & input_a[18]);
  assign popcount21_mjel_core_081 = input_a[13] ^ input_a[14];
  assign popcount21_mjel_core_082 = ~(input_a[8] & input_a[7]);
  assign popcount21_mjel_core_085 = input_a[11] & input_a[4];
  assign popcount21_mjel_core_086 = input_a[11] & input_a[5];
  assign popcount21_mjel_core_089 = ~input_a[6];
  assign popcount21_mjel_core_091 = ~input_a[7];
  assign popcount21_mjel_core_095 = input_a[1] ^ input_a[20];
  assign popcount21_mjel_core_098 = input_a[9] | input_a[7];
  assign popcount21_mjel_core_099 = input_a[0] ^ input_a[18];
  assign popcount21_mjel_core_100 = ~input_a[16];
  assign popcount21_mjel_core_101 = input_a[20] | input_a[16];
  assign popcount21_mjel_core_103 = input_a[3] & input_a[12];
  assign popcount21_mjel_core_104 = ~input_a[15];
  assign popcount21_mjel_core_105_not = ~input_a[18];
  assign popcount21_mjel_core_108 = ~(input_a[0] & input_a[11]);
  assign popcount21_mjel_core_112 = ~(input_a[12] ^ input_a[3]);
  assign popcount21_mjel_core_114 = input_a[16] | input_a[14];
  assign popcount21_mjel_core_116 = ~(input_a[13] ^ input_a[17]);
  assign popcount21_mjel_core_117 = ~(input_a[9] | input_a[0]);
  assign popcount21_mjel_core_120 = ~input_a[11];
  assign popcount21_mjel_core_122 = ~(input_a[13] ^ input_a[14]);
  assign popcount21_mjel_core_124 = input_a[6] | input_a[20];
  assign popcount21_mjel_core_125 = input_a[9] | input_a[0];
  assign popcount21_mjel_core_133 = input_a[18] & input_a[9];
  assign popcount21_mjel_core_134 = input_a[5] | input_a[2];
  assign popcount21_mjel_core_135 = input_a[13] & input_a[16];
  assign popcount21_mjel_core_137_not = ~input_a[4];
  assign popcount21_mjel_core_138 = input_a[20] & input_a[2];
  assign popcount21_mjel_core_139 = input_a[17] ^ input_a[10];
  assign popcount21_mjel_core_140 = ~input_a[2];
  assign popcount21_mjel_core_141 = ~input_a[6];
  assign popcount21_mjel_core_142 = ~input_a[2];
  assign popcount21_mjel_core_144 = input_a[14] | input_a[3];
  assign popcount21_mjel_core_147 = input_a[20] | input_a[14];
  assign popcount21_mjel_core_148 = ~(input_a[2] & input_a[20]);
  assign popcount21_mjel_core_150 = input_a[2] ^ input_a[11];
  assign popcount21_mjel_core_151 = input_a[16] ^ input_a[16];
  assign popcount21_mjel_core_153 = input_a[1] ^ input_a[14];

  assign popcount21_mjel_out[0] = input_a[10];
  assign popcount21_mjel_out[1] = input_a[20];
  assign popcount21_mjel_out[2] = 1'b0;
  assign popcount21_mjel_out[3] = 1'b1;
  assign popcount21_mjel_out[4] = 1'b0;
endmodule