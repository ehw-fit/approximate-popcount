// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.50348
// WCE=20.0
// EP=0.921015%
// Printed PDK parameters:
//  Area=3684610.0
//  Delay=10759810.0
//  Power=121440.0

module popcount39_8ad7(input [38:0] input_a, output [5:0] popcount39_8ad7_out);
  wire popcount39_8ad7_core_041;
  wire popcount39_8ad7_core_042;
  wire popcount39_8ad7_core_043_not;
  wire popcount39_8ad7_core_045;
  wire popcount39_8ad7_core_046;
  wire popcount39_8ad7_core_047;
  wire popcount39_8ad7_core_050;
  wire popcount39_8ad7_core_052;
  wire popcount39_8ad7_core_056;
  wire popcount39_8ad7_core_058;
  wire popcount39_8ad7_core_059;
  wire popcount39_8ad7_core_062;
  wire popcount39_8ad7_core_064;
  wire popcount39_8ad7_core_065;
  wire popcount39_8ad7_core_066;
  wire popcount39_8ad7_core_067;
  wire popcount39_8ad7_core_069;
  wire popcount39_8ad7_core_070;
  wire popcount39_8ad7_core_071;
  wire popcount39_8ad7_core_072;
  wire popcount39_8ad7_core_073;
  wire popcount39_8ad7_core_074;
  wire popcount39_8ad7_core_075;
  wire popcount39_8ad7_core_079;
  wire popcount39_8ad7_core_080;
  wire popcount39_8ad7_core_081;
  wire popcount39_8ad7_core_083;
  wire popcount39_8ad7_core_086;
  wire popcount39_8ad7_core_089;
  wire popcount39_8ad7_core_091;
  wire popcount39_8ad7_core_092;
  wire popcount39_8ad7_core_093;
  wire popcount39_8ad7_core_094;
  wire popcount39_8ad7_core_095;
  wire popcount39_8ad7_core_096;
  wire popcount39_8ad7_core_097;
  wire popcount39_8ad7_core_098;
  wire popcount39_8ad7_core_099;
  wire popcount39_8ad7_core_100;
  wire popcount39_8ad7_core_103;
  wire popcount39_8ad7_core_106;
  wire popcount39_8ad7_core_107;
  wire popcount39_8ad7_core_108;
  wire popcount39_8ad7_core_109;
  wire popcount39_8ad7_core_111;
  wire popcount39_8ad7_core_112;
  wire popcount39_8ad7_core_114;
  wire popcount39_8ad7_core_115;
  wire popcount39_8ad7_core_116;
  wire popcount39_8ad7_core_117;
  wire popcount39_8ad7_core_118;
  wire popcount39_8ad7_core_119;
  wire popcount39_8ad7_core_120;
  wire popcount39_8ad7_core_121;
  wire popcount39_8ad7_core_123;
  wire popcount39_8ad7_core_125;
  wire popcount39_8ad7_core_126;
  wire popcount39_8ad7_core_127;
  wire popcount39_8ad7_core_128;
  wire popcount39_8ad7_core_129;
  wire popcount39_8ad7_core_132;
  wire popcount39_8ad7_core_133;
  wire popcount39_8ad7_core_134;
  wire popcount39_8ad7_core_135;
  wire popcount39_8ad7_core_136_not;
  wire popcount39_8ad7_core_137;
  wire popcount39_8ad7_core_138;
  wire popcount39_8ad7_core_140_not;
  wire popcount39_8ad7_core_141;
  wire popcount39_8ad7_core_142;
  wire popcount39_8ad7_core_143;
  wire popcount39_8ad7_core_144;
  wire popcount39_8ad7_core_145;
  wire popcount39_8ad7_core_146;
  wire popcount39_8ad7_core_149;
  wire popcount39_8ad7_core_154;
  wire popcount39_8ad7_core_155;
  wire popcount39_8ad7_core_156;
  wire popcount39_8ad7_core_157;
  wire popcount39_8ad7_core_159;
  wire popcount39_8ad7_core_160;
  wire popcount39_8ad7_core_161;
  wire popcount39_8ad7_core_162;
  wire popcount39_8ad7_core_165;
  wire popcount39_8ad7_core_166;
  wire popcount39_8ad7_core_167;
  wire popcount39_8ad7_core_168;
  wire popcount39_8ad7_core_169;
  wire popcount39_8ad7_core_170;
  wire popcount39_8ad7_core_172;
  wire popcount39_8ad7_core_173;
  wire popcount39_8ad7_core_177;
  wire popcount39_8ad7_core_178;
  wire popcount39_8ad7_core_180;
  wire popcount39_8ad7_core_181;
  wire popcount39_8ad7_core_182;
  wire popcount39_8ad7_core_183;
  wire popcount39_8ad7_core_185;
  wire popcount39_8ad7_core_189;
  wire popcount39_8ad7_core_190;
  wire popcount39_8ad7_core_192;
  wire popcount39_8ad7_core_193;
  wire popcount39_8ad7_core_194_not;
  wire popcount39_8ad7_core_195;
  wire popcount39_8ad7_core_196;
  wire popcount39_8ad7_core_198;
  wire popcount39_8ad7_core_200;
  wire popcount39_8ad7_core_203;
  wire popcount39_8ad7_core_210;
  wire popcount39_8ad7_core_212;
  wire popcount39_8ad7_core_213;
  wire popcount39_8ad7_core_215;
  wire popcount39_8ad7_core_216;
  wire popcount39_8ad7_core_217;
  wire popcount39_8ad7_core_221_not;
  wire popcount39_8ad7_core_223;
  wire popcount39_8ad7_core_224;
  wire popcount39_8ad7_core_227;
  wire popcount39_8ad7_core_228;
  wire popcount39_8ad7_core_230;
  wire popcount39_8ad7_core_232;
  wire popcount39_8ad7_core_236_not;
  wire popcount39_8ad7_core_238;
  wire popcount39_8ad7_core_239;
  wire popcount39_8ad7_core_246;
  wire popcount39_8ad7_core_247;
  wire popcount39_8ad7_core_248;
  wire popcount39_8ad7_core_249;
  wire popcount39_8ad7_core_250;
  wire popcount39_8ad7_core_251;
  wire popcount39_8ad7_core_252;
  wire popcount39_8ad7_core_253;
  wire popcount39_8ad7_core_258;
  wire popcount39_8ad7_core_260;
  wire popcount39_8ad7_core_261;
  wire popcount39_8ad7_core_262;
  wire popcount39_8ad7_core_265;
  wire popcount39_8ad7_core_266;
  wire popcount39_8ad7_core_267;
  wire popcount39_8ad7_core_268;
  wire popcount39_8ad7_core_269;
  wire popcount39_8ad7_core_271;
  wire popcount39_8ad7_core_272;
  wire popcount39_8ad7_core_273;
  wire popcount39_8ad7_core_274;
  wire popcount39_8ad7_core_279;
  wire popcount39_8ad7_core_280;
  wire popcount39_8ad7_core_282;
  wire popcount39_8ad7_core_283;
  wire popcount39_8ad7_core_284;
  wire popcount39_8ad7_core_287;
  wire popcount39_8ad7_core_288;
  wire popcount39_8ad7_core_290;
  wire popcount39_8ad7_core_292_not;
  wire popcount39_8ad7_core_294;
  wire popcount39_8ad7_core_296;
  wire popcount39_8ad7_core_300;
  wire popcount39_8ad7_core_301;
  wire popcount39_8ad7_core_303;
  wire popcount39_8ad7_core_304;
  wire popcount39_8ad7_core_305;
  wire popcount39_8ad7_core_306;

  assign popcount39_8ad7_core_041 = ~(input_a[22] | input_a[9]);
  assign popcount39_8ad7_core_042 = ~(input_a[16] & input_a[28]);
  assign popcount39_8ad7_core_043_not = ~input_a[36];
  assign popcount39_8ad7_core_045 = input_a[22] | input_a[2];
  assign popcount39_8ad7_core_046 = input_a[2] ^ input_a[35];
  assign popcount39_8ad7_core_047 = ~input_a[8];
  assign popcount39_8ad7_core_050 = ~(input_a[36] | input_a[18]);
  assign popcount39_8ad7_core_052 = ~(input_a[30] | input_a[3]);
  assign popcount39_8ad7_core_056 = input_a[20] & input_a[25];
  assign popcount39_8ad7_core_058 = ~input_a[34];
  assign popcount39_8ad7_core_059 = input_a[4] | input_a[33];
  assign popcount39_8ad7_core_062 = ~(input_a[4] & input_a[25]);
  assign popcount39_8ad7_core_064 = ~(input_a[8] ^ input_a[25]);
  assign popcount39_8ad7_core_065 = ~(input_a[32] & input_a[4]);
  assign popcount39_8ad7_core_066 = input_a[0] | input_a[9];
  assign popcount39_8ad7_core_067 = input_a[12] ^ input_a[14];
  assign popcount39_8ad7_core_069 = input_a[32] ^ input_a[17];
  assign popcount39_8ad7_core_070 = input_a[35] | input_a[5];
  assign popcount39_8ad7_core_071 = ~(input_a[34] ^ input_a[17]);
  assign popcount39_8ad7_core_072 = input_a[15] | input_a[38];
  assign popcount39_8ad7_core_073 = ~(input_a[29] & input_a[25]);
  assign popcount39_8ad7_core_074 = input_a[13] & input_a[2];
  assign popcount39_8ad7_core_075 = input_a[33] ^ input_a[9];
  assign popcount39_8ad7_core_079 = ~(input_a[13] & input_a[30]);
  assign popcount39_8ad7_core_080 = ~(input_a[1] ^ input_a[28]);
  assign popcount39_8ad7_core_081 = input_a[38] ^ input_a[29];
  assign popcount39_8ad7_core_083 = ~(input_a[36] | input_a[7]);
  assign popcount39_8ad7_core_086 = input_a[30] & input_a[18];
  assign popcount39_8ad7_core_089 = ~input_a[23];
  assign popcount39_8ad7_core_091 = ~(input_a[20] ^ input_a[0]);
  assign popcount39_8ad7_core_092 = input_a[3] | input_a[32];
  assign popcount39_8ad7_core_093 = input_a[26] & input_a[32];
  assign popcount39_8ad7_core_094 = input_a[15] & input_a[2];
  assign popcount39_8ad7_core_095 = ~(input_a[27] & input_a[14]);
  assign popcount39_8ad7_core_096 = input_a[27] ^ input_a[26];
  assign popcount39_8ad7_core_097 = ~(input_a[38] | input_a[0]);
  assign popcount39_8ad7_core_098 = ~(input_a[6] | input_a[38]);
  assign popcount39_8ad7_core_099 = input_a[19] | input_a[2];
  assign popcount39_8ad7_core_100 = input_a[7] | input_a[21];
  assign popcount39_8ad7_core_103 = input_a[33] & input_a[35];
  assign popcount39_8ad7_core_106 = ~(input_a[36] & input_a[28]);
  assign popcount39_8ad7_core_107 = input_a[20] | input_a[37];
  assign popcount39_8ad7_core_108 = input_a[22] ^ input_a[28];
  assign popcount39_8ad7_core_109 = ~input_a[21];
  assign popcount39_8ad7_core_111 = ~(input_a[18] ^ input_a[23]);
  assign popcount39_8ad7_core_112 = ~(input_a[5] & input_a[35]);
  assign popcount39_8ad7_core_114 = input_a[0] & input_a[19];
  assign popcount39_8ad7_core_115 = input_a[26] & input_a[23];
  assign popcount39_8ad7_core_116 = input_a[35] ^ input_a[14];
  assign popcount39_8ad7_core_117 = ~(input_a[25] & input_a[8]);
  assign popcount39_8ad7_core_118 = ~(input_a[2] & input_a[16]);
  assign popcount39_8ad7_core_119 = ~(input_a[5] & input_a[11]);
  assign popcount39_8ad7_core_120 = ~(input_a[6] ^ input_a[0]);
  assign popcount39_8ad7_core_121 = ~(input_a[36] ^ input_a[23]);
  assign popcount39_8ad7_core_123 = ~input_a[33];
  assign popcount39_8ad7_core_125 = input_a[28] ^ input_a[27];
  assign popcount39_8ad7_core_126 = ~(input_a[15] & input_a[20]);
  assign popcount39_8ad7_core_127 = ~(input_a[1] | input_a[34]);
  assign popcount39_8ad7_core_128 = input_a[34] ^ input_a[26];
  assign popcount39_8ad7_core_129 = ~input_a[37];
  assign popcount39_8ad7_core_132 = ~(input_a[38] & input_a[10]);
  assign popcount39_8ad7_core_133 = input_a[33] & input_a[25];
  assign popcount39_8ad7_core_134 = input_a[36] | input_a[34];
  assign popcount39_8ad7_core_135 = ~(input_a[31] ^ input_a[11]);
  assign popcount39_8ad7_core_136_not = ~input_a[33];
  assign popcount39_8ad7_core_137 = input_a[8] | input_a[5];
  assign popcount39_8ad7_core_138 = ~(input_a[38] | input_a[18]);
  assign popcount39_8ad7_core_140_not = ~input_a[32];
  assign popcount39_8ad7_core_141 = input_a[20] ^ input_a[35];
  assign popcount39_8ad7_core_142 = ~(input_a[33] & input_a[33]);
  assign popcount39_8ad7_core_143 = input_a[29] ^ input_a[30];
  assign popcount39_8ad7_core_144 = ~(input_a[23] ^ input_a[21]);
  assign popcount39_8ad7_core_145 = input_a[24] & input_a[36];
  assign popcount39_8ad7_core_146 = input_a[24] ^ input_a[0];
  assign popcount39_8ad7_core_149 = input_a[34] | input_a[33];
  assign popcount39_8ad7_core_154 = input_a[35] ^ input_a[32];
  assign popcount39_8ad7_core_155 = ~(input_a[18] ^ input_a[18]);
  assign popcount39_8ad7_core_156 = ~(input_a[18] & input_a[36]);
  assign popcount39_8ad7_core_157 = input_a[10] | input_a[3];
  assign popcount39_8ad7_core_159 = ~(input_a[16] | input_a[32]);
  assign popcount39_8ad7_core_160 = ~(input_a[24] & input_a[16]);
  assign popcount39_8ad7_core_161 = ~input_a[35];
  assign popcount39_8ad7_core_162 = ~(input_a[11] | input_a[2]);
  assign popcount39_8ad7_core_165 = ~(input_a[27] & input_a[37]);
  assign popcount39_8ad7_core_166 = input_a[34] & input_a[35];
  assign popcount39_8ad7_core_167 = input_a[2] & input_a[34];
  assign popcount39_8ad7_core_168 = ~(input_a[17] & input_a[14]);
  assign popcount39_8ad7_core_169 = input_a[35] & input_a[29];
  assign popcount39_8ad7_core_170 = popcount39_8ad7_core_167 | popcount39_8ad7_core_169;
  assign popcount39_8ad7_core_172 = ~(input_a[6] | input_a[23]);
  assign popcount39_8ad7_core_173 = ~(input_a[3] ^ input_a[35]);
  assign popcount39_8ad7_core_177 = input_a[28] & input_a[19];
  assign popcount39_8ad7_core_178 = ~input_a[14];
  assign popcount39_8ad7_core_180 = ~(input_a[32] & input_a[21]);
  assign popcount39_8ad7_core_181 = ~(input_a[7] & input_a[1]);
  assign popcount39_8ad7_core_182 = ~(input_a[13] ^ input_a[20]);
  assign popcount39_8ad7_core_183 = ~(input_a[6] ^ input_a[17]);
  assign popcount39_8ad7_core_185 = ~(input_a[13] ^ input_a[1]);
  assign popcount39_8ad7_core_189 = ~(input_a[8] & input_a[4]);
  assign popcount39_8ad7_core_190 = input_a[3] | input_a[34];
  assign popcount39_8ad7_core_192 = ~(input_a[3] | input_a[4]);
  assign popcount39_8ad7_core_193 = input_a[31] ^ input_a[22];
  assign popcount39_8ad7_core_194_not = ~input_a[25];
  assign popcount39_8ad7_core_195 = input_a[1] | input_a[20];
  assign popcount39_8ad7_core_196 = ~(input_a[38] ^ input_a[9]);
  assign popcount39_8ad7_core_198 = popcount39_8ad7_core_170 & input_a[23];
  assign popcount39_8ad7_core_200 = ~input_a[3];
  assign popcount39_8ad7_core_203 = ~(input_a[22] ^ input_a[22]);
  assign popcount39_8ad7_core_210 = input_a[2] & input_a[11];
  assign popcount39_8ad7_core_212 = input_a[15] & input_a[4];
  assign popcount39_8ad7_core_213 = ~(input_a[21] ^ input_a[2]);
  assign popcount39_8ad7_core_215 = input_a[18] | input_a[35];
  assign popcount39_8ad7_core_216 = input_a[22] & input_a[29];
  assign popcount39_8ad7_core_217 = ~input_a[12];
  assign popcount39_8ad7_core_221_not = ~input_a[14];
  assign popcount39_8ad7_core_223 = ~(input_a[28] & input_a[36]);
  assign popcount39_8ad7_core_224 = ~input_a[27];
  assign popcount39_8ad7_core_227 = ~(input_a[30] ^ input_a[7]);
  assign popcount39_8ad7_core_228 = input_a[8] | input_a[4];
  assign popcount39_8ad7_core_230 = input_a[33] | input_a[34];
  assign popcount39_8ad7_core_232 = input_a[3] ^ input_a[26];
  assign popcount39_8ad7_core_236_not = ~input_a[16];
  assign popcount39_8ad7_core_238 = ~(input_a[25] | input_a[36]);
  assign popcount39_8ad7_core_239 = input_a[27] | input_a[33];
  assign popcount39_8ad7_core_246 = input_a[36] | input_a[4];
  assign popcount39_8ad7_core_247 = ~(input_a[19] | input_a[15]);
  assign popcount39_8ad7_core_248 = input_a[24] | input_a[37];
  assign popcount39_8ad7_core_249 = ~input_a[32];
  assign popcount39_8ad7_core_250 = ~(input_a[38] | input_a[8]);
  assign popcount39_8ad7_core_251 = ~input_a[15];
  assign popcount39_8ad7_core_252 = ~(input_a[32] | input_a[33]);
  assign popcount39_8ad7_core_253 = input_a[31] ^ input_a[11];
  assign popcount39_8ad7_core_258 = ~(input_a[9] & input_a[16]);
  assign popcount39_8ad7_core_260 = ~(input_a[5] & input_a[12]);
  assign popcount39_8ad7_core_261 = input_a[36] & input_a[3];
  assign popcount39_8ad7_core_262 = ~(input_a[16] ^ input_a[13]);
  assign popcount39_8ad7_core_265 = input_a[16] & input_a[32];
  assign popcount39_8ad7_core_266 = popcount39_8ad7_core_170 & input_a[20];
  assign popcount39_8ad7_core_267 = ~(input_a[4] & input_a[30]);
  assign popcount39_8ad7_core_268 = input_a[11] & popcount39_8ad7_core_261;
  assign popcount39_8ad7_core_269 = popcount39_8ad7_core_266 | popcount39_8ad7_core_268;
  assign popcount39_8ad7_core_271 = ~(input_a[8] & input_a[0]);
  assign popcount39_8ad7_core_272 = popcount39_8ad7_core_198 | popcount39_8ad7_core_269;
  assign popcount39_8ad7_core_273 = input_a[14] ^ input_a[9];
  assign popcount39_8ad7_core_274 = input_a[13] & input_a[14];
  assign popcount39_8ad7_core_279 = ~(input_a[35] & input_a[32]);
  assign popcount39_8ad7_core_280 = ~(input_a[15] & input_a[4]);
  assign popcount39_8ad7_core_282 = ~(input_a[28] | input_a[37]);
  assign popcount39_8ad7_core_283 = ~(input_a[3] & input_a[35]);
  assign popcount39_8ad7_core_284 = input_a[34] ^ input_a[21];
  assign popcount39_8ad7_core_287 = input_a[35] & input_a[23];
  assign popcount39_8ad7_core_288 = ~(input_a[20] | input_a[37]);
  assign popcount39_8ad7_core_290 = ~(input_a[19] | input_a[37]);
  assign popcount39_8ad7_core_292_not = ~popcount39_8ad7_core_272;
  assign popcount39_8ad7_core_294 = popcount39_8ad7_core_292_not ^ input_a[32];
  assign popcount39_8ad7_core_296 = popcount39_8ad7_core_272 | input_a[32];
  assign popcount39_8ad7_core_300 = input_a[23] & input_a[1];
  assign popcount39_8ad7_core_301 = ~(input_a[24] & input_a[21]);
  assign popcount39_8ad7_core_303 = input_a[25] & input_a[37];
  assign popcount39_8ad7_core_304 = input_a[35] & input_a[22];
  assign popcount39_8ad7_core_305 = input_a[28] ^ input_a[1];
  assign popcount39_8ad7_core_306 = ~(input_a[18] ^ input_a[32]);

  assign popcount39_8ad7_out[0] = input_a[27];
  assign popcount39_8ad7_out[1] = popcount39_8ad7_core_249;
  assign popcount39_8ad7_out[2] = popcount39_8ad7_core_249;
  assign popcount39_8ad7_out[3] = popcount39_8ad7_core_294;
  assign popcount39_8ad7_out[4] = popcount39_8ad7_core_296;
  assign popcount39_8ad7_out[5] = 1'b0;
endmodule