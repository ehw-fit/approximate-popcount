// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.14092
// WCE=27.0
// EP=0.930441%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount47_um3q(input [46:0] input_a, output [5:0] popcount47_um3q_out);
  wire popcount47_um3q_core_049;
  wire popcount47_um3q_core_050;
  wire popcount47_um3q_core_051;
  wire popcount47_um3q_core_054;
  wire popcount47_um3q_core_056;
  wire popcount47_um3q_core_057;
  wire popcount47_um3q_core_058;
  wire popcount47_um3q_core_059;
  wire popcount47_um3q_core_060;
  wire popcount47_um3q_core_064;
  wire popcount47_um3q_core_065;
  wire popcount47_um3q_core_067;
  wire popcount47_um3q_core_068;
  wire popcount47_um3q_core_069;
  wire popcount47_um3q_core_070;
  wire popcount47_um3q_core_071;
  wire popcount47_um3q_core_072;
  wire popcount47_um3q_core_073;
  wire popcount47_um3q_core_074;
  wire popcount47_um3q_core_075;
  wire popcount47_um3q_core_076;
  wire popcount47_um3q_core_077;
  wire popcount47_um3q_core_079;
  wire popcount47_um3q_core_080;
  wire popcount47_um3q_core_081;
  wire popcount47_um3q_core_082;
  wire popcount47_um3q_core_083;
  wire popcount47_um3q_core_084;
  wire popcount47_um3q_core_088_not;
  wire popcount47_um3q_core_092;
  wire popcount47_um3q_core_095_not;
  wire popcount47_um3q_core_097;
  wire popcount47_um3q_core_098;
  wire popcount47_um3q_core_100;
  wire popcount47_um3q_core_101;
  wire popcount47_um3q_core_102;
  wire popcount47_um3q_core_106;
  wire popcount47_um3q_core_107;
  wire popcount47_um3q_core_111;
  wire popcount47_um3q_core_113;
  wire popcount47_um3q_core_115;
  wire popcount47_um3q_core_118;
  wire popcount47_um3q_core_119;
  wire popcount47_um3q_core_120_not;
  wire popcount47_um3q_core_121;
  wire popcount47_um3q_core_122;
  wire popcount47_um3q_core_125;
  wire popcount47_um3q_core_127;
  wire popcount47_um3q_core_128;
  wire popcount47_um3q_core_129;
  wire popcount47_um3q_core_130;
  wire popcount47_um3q_core_131;
  wire popcount47_um3q_core_134;
  wire popcount47_um3q_core_136;
  wire popcount47_um3q_core_137;
  wire popcount47_um3q_core_138;
  wire popcount47_um3q_core_139;
  wire popcount47_um3q_core_140;
  wire popcount47_um3q_core_141;
  wire popcount47_um3q_core_143;
  wire popcount47_um3q_core_144;
  wire popcount47_um3q_core_145;
  wire popcount47_um3q_core_147;
  wire popcount47_um3q_core_148;
  wire popcount47_um3q_core_149;
  wire popcount47_um3q_core_152;
  wire popcount47_um3q_core_153;
  wire popcount47_um3q_core_154;
  wire popcount47_um3q_core_155;
  wire popcount47_um3q_core_156;
  wire popcount47_um3q_core_157;
  wire popcount47_um3q_core_158;
  wire popcount47_um3q_core_160;
  wire popcount47_um3q_core_161;
  wire popcount47_um3q_core_162;
  wire popcount47_um3q_core_163;
  wire popcount47_um3q_core_164;
  wire popcount47_um3q_core_165;
  wire popcount47_um3q_core_168;
  wire popcount47_um3q_core_169;
  wire popcount47_um3q_core_170;
  wire popcount47_um3q_core_171;
  wire popcount47_um3q_core_172;
  wire popcount47_um3q_core_173;
  wire popcount47_um3q_core_174;
  wire popcount47_um3q_core_175;
  wire popcount47_um3q_core_177;
  wire popcount47_um3q_core_181;
  wire popcount47_um3q_core_184;
  wire popcount47_um3q_core_185;
  wire popcount47_um3q_core_187;
  wire popcount47_um3q_core_189;
  wire popcount47_um3q_core_190;
  wire popcount47_um3q_core_191;
  wire popcount47_um3q_core_192;
  wire popcount47_um3q_core_193;
  wire popcount47_um3q_core_197;
  wire popcount47_um3q_core_198;
  wire popcount47_um3q_core_199;
  wire popcount47_um3q_core_201;
  wire popcount47_um3q_core_202;
  wire popcount47_um3q_core_204;
  wire popcount47_um3q_core_205;
  wire popcount47_um3q_core_208;
  wire popcount47_um3q_core_210;
  wire popcount47_um3q_core_215;
  wire popcount47_um3q_core_216;
  wire popcount47_um3q_core_217;
  wire popcount47_um3q_core_219;
  wire popcount47_um3q_core_220;
  wire popcount47_um3q_core_221_not;
  wire popcount47_um3q_core_223;
  wire popcount47_um3q_core_225;
  wire popcount47_um3q_core_230;
  wire popcount47_um3q_core_232;
  wire popcount47_um3q_core_234;
  wire popcount47_um3q_core_235;
  wire popcount47_um3q_core_236;
  wire popcount47_um3q_core_239;
  wire popcount47_um3q_core_242;
  wire popcount47_um3q_core_244;
  wire popcount47_um3q_core_245;
  wire popcount47_um3q_core_249;
  wire popcount47_um3q_core_250;
  wire popcount47_um3q_core_251;
  wire popcount47_um3q_core_252;
  wire popcount47_um3q_core_253;
  wire popcount47_um3q_core_254;
  wire popcount47_um3q_core_260;
  wire popcount47_um3q_core_261;
  wire popcount47_um3q_core_265;
  wire popcount47_um3q_core_266;
  wire popcount47_um3q_core_268;
  wire popcount47_um3q_core_269;
  wire popcount47_um3q_core_270;
  wire popcount47_um3q_core_271;
  wire popcount47_um3q_core_272;
  wire popcount47_um3q_core_273;
  wire popcount47_um3q_core_274;
  wire popcount47_um3q_core_276_not;
  wire popcount47_um3q_core_279;
  wire popcount47_um3q_core_280;
  wire popcount47_um3q_core_283;
  wire popcount47_um3q_core_284_not;
  wire popcount47_um3q_core_289;
  wire popcount47_um3q_core_293;
  wire popcount47_um3q_core_296;
  wire popcount47_um3q_core_297;
  wire popcount47_um3q_core_298;
  wire popcount47_um3q_core_300;
  wire popcount47_um3q_core_301;
  wire popcount47_um3q_core_302;
  wire popcount47_um3q_core_303;
  wire popcount47_um3q_core_305;
  wire popcount47_um3q_core_306;
  wire popcount47_um3q_core_307;
  wire popcount47_um3q_core_308;
  wire popcount47_um3q_core_315;
  wire popcount47_um3q_core_318;
  wire popcount47_um3q_core_319;
  wire popcount47_um3q_core_320;
  wire popcount47_um3q_core_322;
  wire popcount47_um3q_core_323;
  wire popcount47_um3q_core_324;
  wire popcount47_um3q_core_326;
  wire popcount47_um3q_core_327;
  wire popcount47_um3q_core_329;
  wire popcount47_um3q_core_330;
  wire popcount47_um3q_core_333;
  wire popcount47_um3q_core_334;
  wire popcount47_um3q_core_335;
  wire popcount47_um3q_core_336;
  wire popcount47_um3q_core_337;
  wire popcount47_um3q_core_339;
  wire popcount47_um3q_core_341;
  wire popcount47_um3q_core_342;
  wire popcount47_um3q_core_343;
  wire popcount47_um3q_core_344;
  wire popcount47_um3q_core_347;
  wire popcount47_um3q_core_348;
  wire popcount47_um3q_core_349;
  wire popcount47_um3q_core_350;
  wire popcount47_um3q_core_351;
  wire popcount47_um3q_core_352;
  wire popcount47_um3q_core_354;
  wire popcount47_um3q_core_355;
  wire popcount47_um3q_core_356;
  wire popcount47_um3q_core_357;
  wire popcount47_um3q_core_358;
  wire popcount47_um3q_core_359;
  wire popcount47_um3q_core_360;
  wire popcount47_um3q_core_361;
  wire popcount47_um3q_core_362;
  wire popcount47_um3q_core_363;
  wire popcount47_um3q_core_364;
  wire popcount47_um3q_core_365;
  wire popcount47_um3q_core_366;
  wire popcount47_um3q_core_367;
  wire popcount47_um3q_core_369;
  wire popcount47_um3q_core_370;

  assign popcount47_um3q_core_049 = ~(input_a[36] | input_a[3]);
  assign popcount47_um3q_core_050 = input_a[7] | input_a[27];
  assign popcount47_um3q_core_051 = ~input_a[23];
  assign popcount47_um3q_core_054 = ~input_a[2];
  assign popcount47_um3q_core_056 = input_a[15] & input_a[15];
  assign popcount47_um3q_core_057 = ~input_a[34];
  assign popcount47_um3q_core_058 = input_a[25] & input_a[38];
  assign popcount47_um3q_core_059 = ~input_a[7];
  assign popcount47_um3q_core_060 = input_a[23] & input_a[16];
  assign popcount47_um3q_core_064 = ~input_a[7];
  assign popcount47_um3q_core_065 = input_a[5] | input_a[33];
  assign popcount47_um3q_core_067 = input_a[23] ^ input_a[41];
  assign popcount47_um3q_core_068 = input_a[46] ^ input_a[31];
  assign popcount47_um3q_core_069 = ~input_a[34];
  assign popcount47_um3q_core_070 = ~(input_a[44] & input_a[41]);
  assign popcount47_um3q_core_071 = ~(input_a[45] & input_a[0]);
  assign popcount47_um3q_core_072 = ~(input_a[27] | input_a[37]);
  assign popcount47_um3q_core_073 = input_a[11] & input_a[14];
  assign popcount47_um3q_core_074 = ~(input_a[23] | input_a[39]);
  assign popcount47_um3q_core_075 = ~(input_a[39] | input_a[37]);
  assign popcount47_um3q_core_076 = input_a[37] & input_a[16];
  assign popcount47_um3q_core_077 = ~(input_a[19] ^ input_a[26]);
  assign popcount47_um3q_core_079 = input_a[18] | input_a[40];
  assign popcount47_um3q_core_080 = ~input_a[36];
  assign popcount47_um3q_core_081 = ~(input_a[33] | input_a[31]);
  assign popcount47_um3q_core_082 = input_a[18] & input_a[12];
  assign popcount47_um3q_core_083 = ~(input_a[32] ^ input_a[29]);
  assign popcount47_um3q_core_084 = input_a[16] & input_a[9];
  assign popcount47_um3q_core_088_not = ~input_a[34];
  assign popcount47_um3q_core_092 = input_a[5] | input_a[29];
  assign popcount47_um3q_core_095_not = ~input_a[0];
  assign popcount47_um3q_core_097 = ~(input_a[44] ^ input_a[32]);
  assign popcount47_um3q_core_098 = ~(input_a[28] | input_a[8]);
  assign popcount47_um3q_core_100 = input_a[18] ^ input_a[12];
  assign popcount47_um3q_core_101 = input_a[8] | input_a[28];
  assign popcount47_um3q_core_102 = input_a[15] ^ input_a[37];
  assign popcount47_um3q_core_106 = ~(input_a[3] | input_a[11]);
  assign popcount47_um3q_core_107 = input_a[42] ^ input_a[31];
  assign popcount47_um3q_core_111 = ~(input_a[8] & input_a[3]);
  assign popcount47_um3q_core_113 = input_a[4] | input_a[5];
  assign popcount47_um3q_core_115 = input_a[44] | input_a[39];
  assign popcount47_um3q_core_118 = input_a[30] ^ input_a[12];
  assign popcount47_um3q_core_119 = ~input_a[1];
  assign popcount47_um3q_core_120_not = ~input_a[30];
  assign popcount47_um3q_core_121 = input_a[15] | input_a[25];
  assign popcount47_um3q_core_122 = input_a[36] & input_a[8];
  assign popcount47_um3q_core_125 = ~(input_a[17] ^ input_a[45]);
  assign popcount47_um3q_core_127 = ~input_a[44];
  assign popcount47_um3q_core_128 = input_a[10] ^ input_a[19];
  assign popcount47_um3q_core_129 = ~input_a[29];
  assign popcount47_um3q_core_130 = input_a[18] & input_a[9];
  assign popcount47_um3q_core_131 = input_a[0] ^ input_a[15];
  assign popcount47_um3q_core_134 = ~(input_a[37] & input_a[1]);
  assign popcount47_um3q_core_136 = input_a[18] ^ input_a[42];
  assign popcount47_um3q_core_137 = ~(input_a[2] & input_a[37]);
  assign popcount47_um3q_core_138 = input_a[3] | input_a[34];
  assign popcount47_um3q_core_139 = ~(input_a[15] & input_a[35]);
  assign popcount47_um3q_core_140 = input_a[5] ^ input_a[41];
  assign popcount47_um3q_core_141 = input_a[42] & input_a[21];
  assign popcount47_um3q_core_143 = input_a[14] | input_a[39];
  assign popcount47_um3q_core_144 = input_a[46] & input_a[5];
  assign popcount47_um3q_core_145 = input_a[41] ^ input_a[17];
  assign popcount47_um3q_core_147 = input_a[44] | input_a[25];
  assign popcount47_um3q_core_148 = ~input_a[7];
  assign popcount47_um3q_core_149 = ~input_a[5];
  assign popcount47_um3q_core_152 = ~input_a[21];
  assign popcount47_um3q_core_153 = ~(input_a[36] ^ input_a[17]);
  assign popcount47_um3q_core_154 = ~(input_a[14] | input_a[5]);
  assign popcount47_um3q_core_155 = input_a[43] ^ input_a[5];
  assign popcount47_um3q_core_156 = input_a[31] | input_a[35];
  assign popcount47_um3q_core_157 = ~(input_a[2] ^ input_a[38]);
  assign popcount47_um3q_core_158 = ~input_a[0];
  assign popcount47_um3q_core_160 = input_a[24] | input_a[20];
  assign popcount47_um3q_core_161 = ~(input_a[17] ^ input_a[25]);
  assign popcount47_um3q_core_162 = input_a[1] & input_a[24];
  assign popcount47_um3q_core_163 = ~input_a[38];
  assign popcount47_um3q_core_164 = ~input_a[5];
  assign popcount47_um3q_core_165 = ~input_a[1];
  assign popcount47_um3q_core_168 = input_a[14] & input_a[4];
  assign popcount47_um3q_core_169 = input_a[35] ^ input_a[5];
  assign popcount47_um3q_core_170 = ~(input_a[3] | input_a[37]);
  assign popcount47_um3q_core_171 = input_a[24] ^ input_a[11];
  assign popcount47_um3q_core_172 = ~(input_a[43] ^ input_a[14]);
  assign popcount47_um3q_core_173 = input_a[40] & input_a[3];
  assign popcount47_um3q_core_174 = ~(input_a[24] ^ input_a[22]);
  assign popcount47_um3q_core_175 = input_a[0] | input_a[5];
  assign popcount47_um3q_core_177 = ~(input_a[30] ^ input_a[11]);
  assign popcount47_um3q_core_181 = ~(input_a[24] & input_a[44]);
  assign popcount47_um3q_core_184 = input_a[23] ^ input_a[33];
  assign popcount47_um3q_core_185 = ~(input_a[1] & input_a[35]);
  assign popcount47_um3q_core_187 = ~(input_a[23] ^ input_a[5]);
  assign popcount47_um3q_core_189 = input_a[39] ^ input_a[30];
  assign popcount47_um3q_core_190 = input_a[33] | input_a[12];
  assign popcount47_um3q_core_191 = input_a[29] & input_a[38];
  assign popcount47_um3q_core_192 = ~input_a[17];
  assign popcount47_um3q_core_193 = ~(input_a[35] & input_a[41]);
  assign popcount47_um3q_core_197 = input_a[11] & input_a[13];
  assign popcount47_um3q_core_198 = ~(input_a[17] | input_a[10]);
  assign popcount47_um3q_core_199 = input_a[15] ^ input_a[34];
  assign popcount47_um3q_core_201 = ~(input_a[2] ^ input_a[39]);
  assign popcount47_um3q_core_202 = input_a[46] & input_a[41];
  assign popcount47_um3q_core_204 = ~input_a[21];
  assign popcount47_um3q_core_205 = ~(input_a[46] | input_a[7]);
  assign popcount47_um3q_core_208 = ~(input_a[14] | input_a[40]);
  assign popcount47_um3q_core_210 = ~(input_a[35] & input_a[8]);
  assign popcount47_um3q_core_215 = ~(input_a[18] | input_a[17]);
  assign popcount47_um3q_core_216 = ~input_a[6];
  assign popcount47_um3q_core_217 = input_a[10] & input_a[43];
  assign popcount47_um3q_core_219 = ~input_a[44];
  assign popcount47_um3q_core_220 = ~(input_a[10] ^ input_a[1]);
  assign popcount47_um3q_core_221_not = ~input_a[21];
  assign popcount47_um3q_core_223 = input_a[21] | input_a[19];
  assign popcount47_um3q_core_225 = ~input_a[32];
  assign popcount47_um3q_core_230 = ~(input_a[43] & input_a[14]);
  assign popcount47_um3q_core_232 = ~(input_a[23] | input_a[35]);
  assign popcount47_um3q_core_234 = ~input_a[15];
  assign popcount47_um3q_core_235 = ~(input_a[33] | input_a[21]);
  assign popcount47_um3q_core_236 = input_a[34] ^ input_a[37];
  assign popcount47_um3q_core_239 = input_a[45] ^ input_a[26];
  assign popcount47_um3q_core_242 = ~(input_a[41] & input_a[1]);
  assign popcount47_um3q_core_244 = ~(input_a[29] & input_a[10]);
  assign popcount47_um3q_core_245 = ~(input_a[15] ^ input_a[33]);
  assign popcount47_um3q_core_249 = ~(input_a[13] & input_a[15]);
  assign popcount47_um3q_core_250 = ~(input_a[39] ^ input_a[42]);
  assign popcount47_um3q_core_251 = input_a[20] ^ input_a[13];
  assign popcount47_um3q_core_252 = input_a[30] ^ input_a[45];
  assign popcount47_um3q_core_253 = input_a[1] | input_a[29];
  assign popcount47_um3q_core_254 = ~(input_a[0] | input_a[11]);
  assign popcount47_um3q_core_260 = input_a[10] ^ input_a[15];
  assign popcount47_um3q_core_261 = ~input_a[20];
  assign popcount47_um3q_core_265 = input_a[35] ^ input_a[6];
  assign popcount47_um3q_core_266 = input_a[33] ^ input_a[30];
  assign popcount47_um3q_core_268 = input_a[13] | input_a[15];
  assign popcount47_um3q_core_269 = ~(input_a[8] ^ input_a[39]);
  assign popcount47_um3q_core_270 = input_a[14] & input_a[17];
  assign popcount47_um3q_core_271 = input_a[12] & input_a[11];
  assign popcount47_um3q_core_272 = input_a[38] | input_a[5];
  assign popcount47_um3q_core_273 = ~(input_a[36] | input_a[45]);
  assign popcount47_um3q_core_274 = ~(input_a[33] & input_a[35]);
  assign popcount47_um3q_core_276_not = ~input_a[41];
  assign popcount47_um3q_core_279 = ~(input_a[7] ^ input_a[44]);
  assign popcount47_um3q_core_280 = ~(input_a[12] & input_a[19]);
  assign popcount47_um3q_core_283 = input_a[2] ^ input_a[2];
  assign popcount47_um3q_core_284_not = ~input_a[16];
  assign popcount47_um3q_core_289 = ~(input_a[40] ^ input_a[26]);
  assign popcount47_um3q_core_293 = input_a[12] | input_a[6];
  assign popcount47_um3q_core_296 = input_a[14] ^ input_a[9];
  assign popcount47_um3q_core_297 = input_a[26] | input_a[6];
  assign popcount47_um3q_core_298 = ~(input_a[31] ^ input_a[31]);
  assign popcount47_um3q_core_300 = input_a[35] & input_a[44];
  assign popcount47_um3q_core_301 = ~(input_a[37] & input_a[35]);
  assign popcount47_um3q_core_302 = input_a[31] ^ input_a[15];
  assign popcount47_um3q_core_303 = ~(input_a[15] & input_a[41]);
  assign popcount47_um3q_core_305 = input_a[0] ^ input_a[27];
  assign popcount47_um3q_core_306 = ~input_a[28];
  assign popcount47_um3q_core_307 = ~(input_a[38] & input_a[14]);
  assign popcount47_um3q_core_308 = input_a[23] | input_a[10];
  assign popcount47_um3q_core_315 = ~(input_a[41] | input_a[42]);
  assign popcount47_um3q_core_318 = input_a[14] & input_a[44];
  assign popcount47_um3q_core_319 = ~(input_a[12] ^ input_a[35]);
  assign popcount47_um3q_core_320 = input_a[32] & input_a[18];
  assign popcount47_um3q_core_322 = input_a[20] | input_a[8];
  assign popcount47_um3q_core_323 = ~input_a[25];
  assign popcount47_um3q_core_324 = ~input_a[44];
  assign popcount47_um3q_core_326 = ~input_a[31];
  assign popcount47_um3q_core_327 = input_a[4] & input_a[43];
  assign popcount47_um3q_core_329 = ~(input_a[30] ^ input_a[44]);
  assign popcount47_um3q_core_330 = input_a[38] & input_a[21];
  assign popcount47_um3q_core_333 = input_a[38] & input_a[6];
  assign popcount47_um3q_core_334 = input_a[4] & input_a[33];
  assign popcount47_um3q_core_335 = input_a[30] ^ input_a[27];
  assign popcount47_um3q_core_336 = ~(input_a[16] | input_a[0]);
  assign popcount47_um3q_core_337 = ~input_a[22];
  assign popcount47_um3q_core_339 = ~(input_a[10] & input_a[42]);
  assign popcount47_um3q_core_341 = ~input_a[16];
  assign popcount47_um3q_core_342 = ~input_a[21];
  assign popcount47_um3q_core_343 = input_a[35] & input_a[25];
  assign popcount47_um3q_core_344 = ~(input_a[31] | input_a[27]);
  assign popcount47_um3q_core_347 = input_a[41] & input_a[6];
  assign popcount47_um3q_core_348 = input_a[41] | input_a[30];
  assign popcount47_um3q_core_349 = input_a[44] & input_a[43];
  assign popcount47_um3q_core_350 = ~input_a[28];
  assign popcount47_um3q_core_351 = ~(input_a[37] | input_a[17]);
  assign popcount47_um3q_core_352 = input_a[5] | input_a[44];
  assign popcount47_um3q_core_354 = ~(input_a[30] | input_a[40]);
  assign popcount47_um3q_core_355 = input_a[9] & input_a[8];
  assign popcount47_um3q_core_356 = ~(input_a[21] ^ input_a[45]);
  assign popcount47_um3q_core_357 = input_a[19] & input_a[26];
  assign popcount47_um3q_core_358 = input_a[19] | input_a[9];
  assign popcount47_um3q_core_359 = input_a[4] & input_a[44];
  assign popcount47_um3q_core_360 = ~(input_a[40] | input_a[46]);
  assign popcount47_um3q_core_361 = ~(input_a[17] & input_a[11]);
  assign popcount47_um3q_core_362 = ~(input_a[25] | input_a[28]);
  assign popcount47_um3q_core_363 = ~input_a[16];
  assign popcount47_um3q_core_364 = ~(input_a[46] | input_a[9]);
  assign popcount47_um3q_core_365 = input_a[22] & input_a[42];
  assign popcount47_um3q_core_366 = input_a[2] ^ input_a[17];
  assign popcount47_um3q_core_367 = ~(input_a[23] | input_a[15]);
  assign popcount47_um3q_core_369 = input_a[29] & input_a[37];
  assign popcount47_um3q_core_370 = input_a[23] & input_a[43];

  assign popcount47_um3q_out[0] = input_a[10];
  assign popcount47_um3q_out[1] = input_a[36];
  assign popcount47_um3q_out[2] = input_a[4];
  assign popcount47_um3q_out[3] = input_a[34];
  assign popcount47_um3q_out[4] = 1'b1;
  assign popcount47_um3q_out[5] = 1'b0;
endmodule