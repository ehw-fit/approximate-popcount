// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.76197
// WCE=10.0
// EP=0.823803%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount20_3nqq(input [19:0] input_a, output [4:0] popcount20_3nqq_out);
  wire popcount20_3nqq_core_023;
  wire popcount20_3nqq_core_024;
  wire popcount20_3nqq_core_025;
  wire popcount20_3nqq_core_026;
  wire popcount20_3nqq_core_030_not;
  wire popcount20_3nqq_core_031;
  wire popcount20_3nqq_core_032;
  wire popcount20_3nqq_core_033;
  wire popcount20_3nqq_core_034;
  wire popcount20_3nqq_core_035;
  wire popcount20_3nqq_core_037;
  wire popcount20_3nqq_core_039;
  wire popcount20_3nqq_core_040;
  wire popcount20_3nqq_core_042;
  wire popcount20_3nqq_core_044;
  wire popcount20_3nqq_core_046;
  wire popcount20_3nqq_core_048;
  wire popcount20_3nqq_core_050;
  wire popcount20_3nqq_core_052;
  wire popcount20_3nqq_core_053;
  wire popcount20_3nqq_core_055;
  wire popcount20_3nqq_core_057;
  wire popcount20_3nqq_core_058;
  wire popcount20_3nqq_core_059;
  wire popcount20_3nqq_core_060;
  wire popcount20_3nqq_core_061;
  wire popcount20_3nqq_core_062;
  wire popcount20_3nqq_core_063;
  wire popcount20_3nqq_core_064;
  wire popcount20_3nqq_core_066;
  wire popcount20_3nqq_core_067;
  wire popcount20_3nqq_core_068;
  wire popcount20_3nqq_core_069;
  wire popcount20_3nqq_core_071;
  wire popcount20_3nqq_core_072;
  wire popcount20_3nqq_core_073;
  wire popcount20_3nqq_core_075;
  wire popcount20_3nqq_core_076;
  wire popcount20_3nqq_core_078;
  wire popcount20_3nqq_core_079;
  wire popcount20_3nqq_core_081;
  wire popcount20_3nqq_core_082;
  wire popcount20_3nqq_core_083;
  wire popcount20_3nqq_core_085;
  wire popcount20_3nqq_core_087_not;
  wire popcount20_3nqq_core_088;
  wire popcount20_3nqq_core_089;
  wire popcount20_3nqq_core_090;
  wire popcount20_3nqq_core_092;
  wire popcount20_3nqq_core_093;
  wire popcount20_3nqq_core_094;
  wire popcount20_3nqq_core_097;
  wire popcount20_3nqq_core_098;
  wire popcount20_3nqq_core_103;
  wire popcount20_3nqq_core_104;
  wire popcount20_3nqq_core_105;
  wire popcount20_3nqq_core_108;
  wire popcount20_3nqq_core_109;
  wire popcount20_3nqq_core_110;
  wire popcount20_3nqq_core_112;
  wire popcount20_3nqq_core_113;
  wire popcount20_3nqq_core_114;
  wire popcount20_3nqq_core_115;
  wire popcount20_3nqq_core_117;
  wire popcount20_3nqq_core_118_not;
  wire popcount20_3nqq_core_121;
  wire popcount20_3nqq_core_122;
  wire popcount20_3nqq_core_125;
  wire popcount20_3nqq_core_128_not;
  wire popcount20_3nqq_core_131;
  wire popcount20_3nqq_core_132;
  wire popcount20_3nqq_core_133;
  wire popcount20_3nqq_core_134;
  wire popcount20_3nqq_core_135;
  wire popcount20_3nqq_core_137;
  wire popcount20_3nqq_core_138_not;
  wire popcount20_3nqq_core_139;
  wire popcount20_3nqq_core_140;
  wire popcount20_3nqq_core_141;
  wire popcount20_3nqq_core_143;
  wire popcount20_3nqq_core_145;

  assign popcount20_3nqq_core_023 = input_a[11] ^ input_a[18];
  assign popcount20_3nqq_core_024 = ~(input_a[12] | input_a[13]);
  assign popcount20_3nqq_core_025 = input_a[1] & input_a[17];
  assign popcount20_3nqq_core_026 = ~input_a[2];
  assign popcount20_3nqq_core_030_not = ~input_a[14];
  assign popcount20_3nqq_core_031 = ~input_a[1];
  assign popcount20_3nqq_core_032 = ~(input_a[10] ^ input_a[6]);
  assign popcount20_3nqq_core_033 = input_a[11] | input_a[14];
  assign popcount20_3nqq_core_034 = ~(input_a[12] | input_a[8]);
  assign popcount20_3nqq_core_035 = ~(input_a[3] & input_a[7]);
  assign popcount20_3nqq_core_037 = input_a[7] | input_a[4];
  assign popcount20_3nqq_core_039 = input_a[5] & input_a[5];
  assign popcount20_3nqq_core_040 = ~input_a[1];
  assign popcount20_3nqq_core_042 = ~input_a[18];
  assign popcount20_3nqq_core_044 = ~(input_a[11] ^ input_a[11]);
  assign popcount20_3nqq_core_046 = input_a[4] & input_a[0];
  assign popcount20_3nqq_core_048 = ~(input_a[11] | input_a[2]);
  assign popcount20_3nqq_core_050 = ~(input_a[2] ^ input_a[0]);
  assign popcount20_3nqq_core_052 = ~(input_a[8] & input_a[8]);
  assign popcount20_3nqq_core_053 = ~(input_a[12] ^ input_a[10]);
  assign popcount20_3nqq_core_055 = input_a[4] & input_a[17];
  assign popcount20_3nqq_core_057 = input_a[15] & input_a[14];
  assign popcount20_3nqq_core_058 = input_a[12] | input_a[12];
  assign popcount20_3nqq_core_059 = input_a[18] & input_a[1];
  assign popcount20_3nqq_core_060 = ~(input_a[11] & input_a[14]);
  assign popcount20_3nqq_core_061 = input_a[2] & input_a[11];
  assign popcount20_3nqq_core_062 = input_a[9] | input_a[2];
  assign popcount20_3nqq_core_063 = input_a[1] & input_a[7];
  assign popcount20_3nqq_core_064 = ~input_a[16];
  assign popcount20_3nqq_core_066 = ~(input_a[18] & input_a[2]);
  assign popcount20_3nqq_core_067 = input_a[11] | input_a[4];
  assign popcount20_3nqq_core_068 = ~(input_a[19] ^ input_a[5]);
  assign popcount20_3nqq_core_069 = input_a[7] | input_a[18];
  assign popcount20_3nqq_core_071 = ~input_a[7];
  assign popcount20_3nqq_core_072 = input_a[0] ^ input_a[2];
  assign popcount20_3nqq_core_073 = input_a[2] ^ input_a[18];
  assign popcount20_3nqq_core_075 = ~(input_a[4] | input_a[4]);
  assign popcount20_3nqq_core_076 = input_a[8] ^ input_a[1];
  assign popcount20_3nqq_core_078 = ~input_a[4];
  assign popcount20_3nqq_core_079 = ~input_a[1];
  assign popcount20_3nqq_core_081 = ~(input_a[3] ^ input_a[12]);
  assign popcount20_3nqq_core_082 = input_a[14] ^ input_a[3];
  assign popcount20_3nqq_core_083 = input_a[5] & input_a[2];
  assign popcount20_3nqq_core_085 = ~input_a[12];
  assign popcount20_3nqq_core_087_not = ~input_a[14];
  assign popcount20_3nqq_core_088 = ~(input_a[1] | input_a[3]);
  assign popcount20_3nqq_core_089 = ~(input_a[5] ^ input_a[9]);
  assign popcount20_3nqq_core_090 = input_a[5] ^ input_a[14];
  assign popcount20_3nqq_core_092 = ~input_a[5];
  assign popcount20_3nqq_core_093 = input_a[18] ^ input_a[7];
  assign popcount20_3nqq_core_094 = input_a[18] & input_a[2];
  assign popcount20_3nqq_core_097 = ~input_a[9];
  assign popcount20_3nqq_core_098 = input_a[18] | input_a[4];
  assign popcount20_3nqq_core_103 = ~input_a[1];
  assign popcount20_3nqq_core_104 = input_a[17] | input_a[4];
  assign popcount20_3nqq_core_105 = input_a[6] ^ input_a[17];
  assign popcount20_3nqq_core_108 = ~(input_a[13] | input_a[3]);
  assign popcount20_3nqq_core_109 = ~(input_a[7] | input_a[3]);
  assign popcount20_3nqq_core_110 = input_a[18] ^ input_a[4];
  assign popcount20_3nqq_core_112 = input_a[10] | input_a[17];
  assign popcount20_3nqq_core_113 = ~(input_a[16] | input_a[10]);
  assign popcount20_3nqq_core_114 = ~(input_a[14] ^ input_a[18]);
  assign popcount20_3nqq_core_115 = input_a[1] ^ input_a[1];
  assign popcount20_3nqq_core_117 = input_a[2] | input_a[12];
  assign popcount20_3nqq_core_118_not = ~input_a[13];
  assign popcount20_3nqq_core_121 = ~(input_a[14] & input_a[3]);
  assign popcount20_3nqq_core_122 = input_a[0] | input_a[0];
  assign popcount20_3nqq_core_125 = ~input_a[14];
  assign popcount20_3nqq_core_128_not = ~input_a[10];
  assign popcount20_3nqq_core_131 = ~(input_a[0] & input_a[12]);
  assign popcount20_3nqq_core_132 = ~(input_a[8] & input_a[3]);
  assign popcount20_3nqq_core_133 = ~(input_a[15] | input_a[2]);
  assign popcount20_3nqq_core_134 = ~(input_a[9] ^ input_a[1]);
  assign popcount20_3nqq_core_135 = input_a[9] & input_a[8];
  assign popcount20_3nqq_core_137 = input_a[5] & input_a[14];
  assign popcount20_3nqq_core_138_not = ~input_a[19];
  assign popcount20_3nqq_core_139 = ~(input_a[2] | input_a[15]);
  assign popcount20_3nqq_core_140 = ~(input_a[8] ^ input_a[13]);
  assign popcount20_3nqq_core_141 = ~input_a[18];
  assign popcount20_3nqq_core_143 = ~(input_a[9] & input_a[3]);
  assign popcount20_3nqq_core_145 = ~(input_a[3] & input_a[16]);

  assign popcount20_3nqq_out[0] = input_a[0];
  assign popcount20_3nqq_out[1] = input_a[19];
  assign popcount20_3nqq_out[2] = 1'b0;
  assign popcount20_3nqq_out[3] = 1'b1;
  assign popcount20_3nqq_out[4] = 1'b0;
endmodule