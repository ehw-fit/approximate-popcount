// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.72677
// WCE=17.0
// EP=0.888465%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount30_3jmp(input [29:0] input_a, output [4:0] popcount30_3jmp_out);
  wire popcount30_3jmp_core_035;
  wire popcount30_3jmp_core_036;
  wire popcount30_3jmp_core_037;
  wire popcount30_3jmp_core_044;
  wire popcount30_3jmp_core_045;
  wire popcount30_3jmp_core_046;
  wire popcount30_3jmp_core_047_not;
  wire popcount30_3jmp_core_048;
  wire popcount30_3jmp_core_049;
  wire popcount30_3jmp_core_055;
  wire popcount30_3jmp_core_058;
  wire popcount30_3jmp_core_062;
  wire popcount30_3jmp_core_063;
  wire popcount30_3jmp_core_064;
  wire popcount30_3jmp_core_066;
  wire popcount30_3jmp_core_067;
  wire popcount30_3jmp_core_068;
  wire popcount30_3jmp_core_069;
  wire popcount30_3jmp_core_070;
  wire popcount30_3jmp_core_071;
  wire popcount30_3jmp_core_072;
  wire popcount30_3jmp_core_073;
  wire popcount30_3jmp_core_075;
  wire popcount30_3jmp_core_077;
  wire popcount30_3jmp_core_078;
  wire popcount30_3jmp_core_079;
  wire popcount30_3jmp_core_080;
  wire popcount30_3jmp_core_081;
  wire popcount30_3jmp_core_082;
  wire popcount30_3jmp_core_083;
  wire popcount30_3jmp_core_088;
  wire popcount30_3jmp_core_089;
  wire popcount30_3jmp_core_091;
  wire popcount30_3jmp_core_092;
  wire popcount30_3jmp_core_093;
  wire popcount30_3jmp_core_094;
  wire popcount30_3jmp_core_095;
  wire popcount30_3jmp_core_096;
  wire popcount30_3jmp_core_097;
  wire popcount30_3jmp_core_098;
  wire popcount30_3jmp_core_099;
  wire popcount30_3jmp_core_100;
  wire popcount30_3jmp_core_102;
  wire popcount30_3jmp_core_103;
  wire popcount30_3jmp_core_104;
  wire popcount30_3jmp_core_107;
  wire popcount30_3jmp_core_108;
  wire popcount30_3jmp_core_110;
  wire popcount30_3jmp_core_111;
  wire popcount30_3jmp_core_112;
  wire popcount30_3jmp_core_113;
  wire popcount30_3jmp_core_116;
  wire popcount30_3jmp_core_120;
  wire popcount30_3jmp_core_121;
  wire popcount30_3jmp_core_122;
  wire popcount30_3jmp_core_123;
  wire popcount30_3jmp_core_125;
  wire popcount30_3jmp_core_126;
  wire popcount30_3jmp_core_133;
  wire popcount30_3jmp_core_134;
  wire popcount30_3jmp_core_135;
  wire popcount30_3jmp_core_136;
  wire popcount30_3jmp_core_137;
  wire popcount30_3jmp_core_141;
  wire popcount30_3jmp_core_142;
  wire popcount30_3jmp_core_143;
  wire popcount30_3jmp_core_144;
  wire popcount30_3jmp_core_145;
  wire popcount30_3jmp_core_148;
  wire popcount30_3jmp_core_149;
  wire popcount30_3jmp_core_151;
  wire popcount30_3jmp_core_153;
  wire popcount30_3jmp_core_154;
  wire popcount30_3jmp_core_155;
  wire popcount30_3jmp_core_156;
  wire popcount30_3jmp_core_157;
  wire popcount30_3jmp_core_158;
  wire popcount30_3jmp_core_160;
  wire popcount30_3jmp_core_161;
  wire popcount30_3jmp_core_162;
  wire popcount30_3jmp_core_163;
  wire popcount30_3jmp_core_164;
  wire popcount30_3jmp_core_165;
  wire popcount30_3jmp_core_167;
  wire popcount30_3jmp_core_170;
  wire popcount30_3jmp_core_172;
  wire popcount30_3jmp_core_173;
  wire popcount30_3jmp_core_174;
  wire popcount30_3jmp_core_175;
  wire popcount30_3jmp_core_177;
  wire popcount30_3jmp_core_178;
  wire popcount30_3jmp_core_180_not;
  wire popcount30_3jmp_core_181;
  wire popcount30_3jmp_core_183;
  wire popcount30_3jmp_core_184;
  wire popcount30_3jmp_core_185;
  wire popcount30_3jmp_core_189;
  wire popcount30_3jmp_core_190;
  wire popcount30_3jmp_core_191;
  wire popcount30_3jmp_core_194;
  wire popcount30_3jmp_core_195;
  wire popcount30_3jmp_core_196;
  wire popcount30_3jmp_core_197;
  wire popcount30_3jmp_core_198;
  wire popcount30_3jmp_core_199;
  wire popcount30_3jmp_core_201;
  wire popcount30_3jmp_core_203;
  wire popcount30_3jmp_core_204;
  wire popcount30_3jmp_core_205;
  wire popcount30_3jmp_core_207;
  wire popcount30_3jmp_core_209;
  wire popcount30_3jmp_core_210;
  wire popcount30_3jmp_core_211;
  wire popcount30_3jmp_core_212;

  assign popcount30_3jmp_core_035 = ~(input_a[11] & input_a[17]);
  assign popcount30_3jmp_core_036 = ~input_a[21];
  assign popcount30_3jmp_core_037 = ~(input_a[12] | input_a[10]);
  assign popcount30_3jmp_core_044 = ~(input_a[10] & input_a[5]);
  assign popcount30_3jmp_core_045 = ~(input_a[19] ^ input_a[14]);
  assign popcount30_3jmp_core_046 = ~input_a[0];
  assign popcount30_3jmp_core_047_not = ~input_a[1];
  assign popcount30_3jmp_core_048 = input_a[15] & input_a[6];
  assign popcount30_3jmp_core_049 = ~(input_a[21] ^ input_a[10]);
  assign popcount30_3jmp_core_055 = ~(input_a[29] | input_a[10]);
  assign popcount30_3jmp_core_058 = ~(input_a[24] ^ input_a[22]);
  assign popcount30_3jmp_core_062 = ~input_a[26];
  assign popcount30_3jmp_core_063 = input_a[6] ^ input_a[12];
  assign popcount30_3jmp_core_064 = ~(input_a[20] & input_a[14]);
  assign popcount30_3jmp_core_066 = input_a[27] & input_a[28];
  assign popcount30_3jmp_core_067 = ~(input_a[23] ^ input_a[3]);
  assign popcount30_3jmp_core_068 = input_a[21] | input_a[6];
  assign popcount30_3jmp_core_069 = ~(input_a[28] & input_a[21]);
  assign popcount30_3jmp_core_070 = ~input_a[15];
  assign popcount30_3jmp_core_071 = input_a[21] | input_a[0];
  assign popcount30_3jmp_core_072 = input_a[16] ^ input_a[25];
  assign popcount30_3jmp_core_073 = ~(input_a[26] ^ input_a[19]);
  assign popcount30_3jmp_core_075 = ~input_a[14];
  assign popcount30_3jmp_core_077 = input_a[1] | input_a[10];
  assign popcount30_3jmp_core_078 = ~(input_a[8] | input_a[24]);
  assign popcount30_3jmp_core_079 = ~(input_a[24] | input_a[7]);
  assign popcount30_3jmp_core_080 = ~(input_a[1] ^ input_a[13]);
  assign popcount30_3jmp_core_081 = ~(input_a[5] & input_a[23]);
  assign popcount30_3jmp_core_082 = input_a[0] & input_a[20];
  assign popcount30_3jmp_core_083 = input_a[27] ^ input_a[21];
  assign popcount30_3jmp_core_088 = input_a[17] | input_a[4];
  assign popcount30_3jmp_core_089 = input_a[16] & input_a[13];
  assign popcount30_3jmp_core_091 = ~input_a[11];
  assign popcount30_3jmp_core_092 = ~(input_a[26] ^ input_a[18]);
  assign popcount30_3jmp_core_093 = input_a[17] ^ input_a[18];
  assign popcount30_3jmp_core_094 = input_a[18] ^ input_a[20];
  assign popcount30_3jmp_core_095 = ~(input_a[12] ^ input_a[3]);
  assign popcount30_3jmp_core_096 = input_a[26] & input_a[29];
  assign popcount30_3jmp_core_097 = ~(input_a[21] ^ input_a[21]);
  assign popcount30_3jmp_core_098 = input_a[8] & input_a[12];
  assign popcount30_3jmp_core_099 = input_a[15] | input_a[12];
  assign popcount30_3jmp_core_100 = input_a[26] ^ input_a[29];
  assign popcount30_3jmp_core_102 = ~(input_a[9] & input_a[27]);
  assign popcount30_3jmp_core_103 = ~(input_a[20] | input_a[3]);
  assign popcount30_3jmp_core_104 = input_a[22] | input_a[3];
  assign popcount30_3jmp_core_107 = ~(input_a[16] | input_a[26]);
  assign popcount30_3jmp_core_108 = input_a[8] | input_a[22];
  assign popcount30_3jmp_core_110 = ~(input_a[12] ^ input_a[10]);
  assign popcount30_3jmp_core_111 = input_a[3] & input_a[14];
  assign popcount30_3jmp_core_112 = input_a[1] ^ input_a[16];
  assign popcount30_3jmp_core_113 = input_a[20] ^ input_a[20];
  assign popcount30_3jmp_core_116 = ~(input_a[10] | input_a[28]);
  assign popcount30_3jmp_core_120 = ~(input_a[5] ^ input_a[25]);
  assign popcount30_3jmp_core_121 = input_a[15] & input_a[28];
  assign popcount30_3jmp_core_122 = ~(input_a[15] ^ input_a[17]);
  assign popcount30_3jmp_core_123 = ~(input_a[9] ^ input_a[24]);
  assign popcount30_3jmp_core_125 = ~(input_a[13] ^ input_a[4]);
  assign popcount30_3jmp_core_126 = ~input_a[14];
  assign popcount30_3jmp_core_133 = input_a[16] ^ input_a[19];
  assign popcount30_3jmp_core_134 = input_a[13] ^ input_a[23];
  assign popcount30_3jmp_core_135 = input_a[11] ^ input_a[11];
  assign popcount30_3jmp_core_136 = ~(input_a[22] | input_a[23]);
  assign popcount30_3jmp_core_137 = input_a[25] ^ input_a[19];
  assign popcount30_3jmp_core_141 = input_a[25] ^ input_a[14];
  assign popcount30_3jmp_core_142 = ~(input_a[0] ^ input_a[26]);
  assign popcount30_3jmp_core_143 = ~(input_a[17] & input_a[12]);
  assign popcount30_3jmp_core_144 = input_a[29] ^ input_a[0];
  assign popcount30_3jmp_core_145 = input_a[20] ^ input_a[7];
  assign popcount30_3jmp_core_148 = ~(input_a[27] & input_a[29]);
  assign popcount30_3jmp_core_149 = ~(input_a[7] | input_a[5]);
  assign popcount30_3jmp_core_151 = ~(input_a[23] & input_a[1]);
  assign popcount30_3jmp_core_153 = input_a[5] & input_a[6];
  assign popcount30_3jmp_core_154 = ~input_a[6];
  assign popcount30_3jmp_core_155 = ~(input_a[0] & input_a[23]);
  assign popcount30_3jmp_core_156 = ~(input_a[11] & input_a[13]);
  assign popcount30_3jmp_core_157 = ~(input_a[13] | input_a[6]);
  assign popcount30_3jmp_core_158 = ~input_a[12];
  assign popcount30_3jmp_core_160 = ~(input_a[5] ^ input_a[3]);
  assign popcount30_3jmp_core_161 = ~input_a[15];
  assign popcount30_3jmp_core_162 = input_a[11] & input_a[29];
  assign popcount30_3jmp_core_163 = ~(input_a[13] ^ input_a[21]);
  assign popcount30_3jmp_core_164 = ~input_a[28];
  assign popcount30_3jmp_core_165 = ~(input_a[15] ^ input_a[19]);
  assign popcount30_3jmp_core_167 = ~(input_a[18] & input_a[18]);
  assign popcount30_3jmp_core_170 = ~(input_a[12] ^ input_a[6]);
  assign popcount30_3jmp_core_172 = input_a[14] | input_a[25];
  assign popcount30_3jmp_core_173 = input_a[5] & input_a[11];
  assign popcount30_3jmp_core_174 = ~(input_a[28] | input_a[1]);
  assign popcount30_3jmp_core_175 = ~(input_a[27] | input_a[20]);
  assign popcount30_3jmp_core_177 = input_a[9] ^ input_a[13];
  assign popcount30_3jmp_core_178 = input_a[3] | input_a[9];
  assign popcount30_3jmp_core_180_not = ~input_a[2];
  assign popcount30_3jmp_core_181 = input_a[19] ^ input_a[20];
  assign popcount30_3jmp_core_183 = ~(input_a[5] & input_a[2]);
  assign popcount30_3jmp_core_184 = input_a[21] | input_a[20];
  assign popcount30_3jmp_core_185 = ~(input_a[7] ^ input_a[9]);
  assign popcount30_3jmp_core_189 = ~(input_a[19] | input_a[14]);
  assign popcount30_3jmp_core_190 = ~(input_a[6] & input_a[29]);
  assign popcount30_3jmp_core_191 = input_a[11] ^ input_a[29];
  assign popcount30_3jmp_core_194 = ~input_a[27];
  assign popcount30_3jmp_core_195 = ~(input_a[12] & input_a[23]);
  assign popcount30_3jmp_core_196 = ~input_a[27];
  assign popcount30_3jmp_core_197 = input_a[7] ^ input_a[15];
  assign popcount30_3jmp_core_198 = input_a[3] & input_a[6];
  assign popcount30_3jmp_core_199 = input_a[15] ^ input_a[23];
  assign popcount30_3jmp_core_201 = input_a[14] ^ input_a[25];
  assign popcount30_3jmp_core_203 = input_a[19] ^ input_a[23];
  assign popcount30_3jmp_core_204 = input_a[25] & input_a[18];
  assign popcount30_3jmp_core_205 = input_a[0] ^ input_a[6];
  assign popcount30_3jmp_core_207 = ~input_a[29];
  assign popcount30_3jmp_core_209 = ~(input_a[17] & input_a[8]);
  assign popcount30_3jmp_core_210 = input_a[23] ^ input_a[8];
  assign popcount30_3jmp_core_211 = ~(input_a[19] ^ input_a[26]);
  assign popcount30_3jmp_core_212 = input_a[15] & input_a[9];

  assign popcount30_3jmp_out[0] = 1'b1;
  assign popcount30_3jmp_out[1] = 1'b0;
  assign popcount30_3jmp_out[2] = 1'b0;
  assign popcount30_3jmp_out[3] = 1'b0;
  assign popcount30_3jmp_out[4] = 1'b1;
endmodule