// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.5701
// WCE=21.0
// EP=0.877614%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount43_0kbs(input [42:0] input_a, output [5:0] popcount43_0kbs_out);
  wire popcount43_0kbs_core_045;
  wire popcount43_0kbs_core_049;
  wire popcount43_0kbs_core_050;
  wire popcount43_0kbs_core_052;
  wire popcount43_0kbs_core_053;
  wire popcount43_0kbs_core_054;
  wire popcount43_0kbs_core_058;
  wire popcount43_0kbs_core_059;
  wire popcount43_0kbs_core_061;
  wire popcount43_0kbs_core_063;
  wire popcount43_0kbs_core_064;
  wire popcount43_0kbs_core_069;
  wire popcount43_0kbs_core_070;
  wire popcount43_0kbs_core_074;
  wire popcount43_0kbs_core_075;
  wire popcount43_0kbs_core_076;
  wire popcount43_0kbs_core_077;
  wire popcount43_0kbs_core_078;
  wire popcount43_0kbs_core_079;
  wire popcount43_0kbs_core_080;
  wire popcount43_0kbs_core_081;
  wire popcount43_0kbs_core_082;
  wire popcount43_0kbs_core_083;
  wire popcount43_0kbs_core_086;
  wire popcount43_0kbs_core_087;
  wire popcount43_0kbs_core_088;
  wire popcount43_0kbs_core_089;
  wire popcount43_0kbs_core_090;
  wire popcount43_0kbs_core_091;
  wire popcount43_0kbs_core_092;
  wire popcount43_0kbs_core_093;
  wire popcount43_0kbs_core_095;
  wire popcount43_0kbs_core_096;
  wire popcount43_0kbs_core_097;
  wire popcount43_0kbs_core_100;
  wire popcount43_0kbs_core_103;
  wire popcount43_0kbs_core_106;
  wire popcount43_0kbs_core_107;
  wire popcount43_0kbs_core_108;
  wire popcount43_0kbs_core_110;
  wire popcount43_0kbs_core_111;
  wire popcount43_0kbs_core_112;
  wire popcount43_0kbs_core_114;
  wire popcount43_0kbs_core_116;
  wire popcount43_0kbs_core_117;
  wire popcount43_0kbs_core_118;
  wire popcount43_0kbs_core_119;
  wire popcount43_0kbs_core_120;
  wire popcount43_0kbs_core_125;
  wire popcount43_0kbs_core_126;
  wire popcount43_0kbs_core_127;
  wire popcount43_0kbs_core_129;
  wire popcount43_0kbs_core_130;
  wire popcount43_0kbs_core_132;
  wire popcount43_0kbs_core_135;
  wire popcount43_0kbs_core_136;
  wire popcount43_0kbs_core_137;
  wire popcount43_0kbs_core_138;
  wire popcount43_0kbs_core_139;
  wire popcount43_0kbs_core_140;
  wire popcount43_0kbs_core_141;
  wire popcount43_0kbs_core_142;
  wire popcount43_0kbs_core_143;
  wire popcount43_0kbs_core_144;
  wire popcount43_0kbs_core_146;
  wire popcount43_0kbs_core_147;
  wire popcount43_0kbs_core_148;
  wire popcount43_0kbs_core_149;
  wire popcount43_0kbs_core_150_not;
  wire popcount43_0kbs_core_151;
  wire popcount43_0kbs_core_156;
  wire popcount43_0kbs_core_157;
  wire popcount43_0kbs_core_158;
  wire popcount43_0kbs_core_159_not;
  wire popcount43_0kbs_core_160;
  wire popcount43_0kbs_core_161;
  wire popcount43_0kbs_core_162;
  wire popcount43_0kbs_core_163;
  wire popcount43_0kbs_core_164;
  wire popcount43_0kbs_core_167;
  wire popcount43_0kbs_core_169;
  wire popcount43_0kbs_core_170;
  wire popcount43_0kbs_core_173;
  wire popcount43_0kbs_core_174;
  wire popcount43_0kbs_core_175;
  wire popcount43_0kbs_core_176;
  wire popcount43_0kbs_core_177;
  wire popcount43_0kbs_core_178;
  wire popcount43_0kbs_core_179;
  wire popcount43_0kbs_core_181;
  wire popcount43_0kbs_core_182;
  wire popcount43_0kbs_core_186;
  wire popcount43_0kbs_core_187;
  wire popcount43_0kbs_core_190;
  wire popcount43_0kbs_core_191;
  wire popcount43_0kbs_core_192;
  wire popcount43_0kbs_core_195;
  wire popcount43_0kbs_core_196;
  wire popcount43_0kbs_core_197;
  wire popcount43_0kbs_core_198;
  wire popcount43_0kbs_core_199;
  wire popcount43_0kbs_core_200;
  wire popcount43_0kbs_core_202;
  wire popcount43_0kbs_core_203;
  wire popcount43_0kbs_core_204;
  wire popcount43_0kbs_core_205;
  wire popcount43_0kbs_core_207;
  wire popcount43_0kbs_core_212;
  wire popcount43_0kbs_core_215;
  wire popcount43_0kbs_core_216;
  wire popcount43_0kbs_core_218;
  wire popcount43_0kbs_core_222;
  wire popcount43_0kbs_core_227;
  wire popcount43_0kbs_core_229;
  wire popcount43_0kbs_core_231_not;
  wire popcount43_0kbs_core_232;
  wire popcount43_0kbs_core_234;
  wire popcount43_0kbs_core_235;
  wire popcount43_0kbs_core_236;
  wire popcount43_0kbs_core_237;
  wire popcount43_0kbs_core_238;
  wire popcount43_0kbs_core_239;
  wire popcount43_0kbs_core_240;
  wire popcount43_0kbs_core_242;
  wire popcount43_0kbs_core_243;
  wire popcount43_0kbs_core_244;
  wire popcount43_0kbs_core_245;
  wire popcount43_0kbs_core_247;
  wire popcount43_0kbs_core_251;
  wire popcount43_0kbs_core_253;
  wire popcount43_0kbs_core_254;
  wire popcount43_0kbs_core_256;
  wire popcount43_0kbs_core_258;
  wire popcount43_0kbs_core_259_not;
  wire popcount43_0kbs_core_260;
  wire popcount43_0kbs_core_262;
  wire popcount43_0kbs_core_263;
  wire popcount43_0kbs_core_266;
  wire popcount43_0kbs_core_267;
  wire popcount43_0kbs_core_268;
  wire popcount43_0kbs_core_269;
  wire popcount43_0kbs_core_270;
  wire popcount43_0kbs_core_272;
  wire popcount43_0kbs_core_275;
  wire popcount43_0kbs_core_277;
  wire popcount43_0kbs_core_281;
  wire popcount43_0kbs_core_282;
  wire popcount43_0kbs_core_283;
  wire popcount43_0kbs_core_286;
  wire popcount43_0kbs_core_287;
  wire popcount43_0kbs_core_288;
  wire popcount43_0kbs_core_290;
  wire popcount43_0kbs_core_292;
  wire popcount43_0kbs_core_294;
  wire popcount43_0kbs_core_295;
  wire popcount43_0kbs_core_297;
  wire popcount43_0kbs_core_299;
  wire popcount43_0kbs_core_300;
  wire popcount43_0kbs_core_301_not;
  wire popcount43_0kbs_core_302;
  wire popcount43_0kbs_core_303;
  wire popcount43_0kbs_core_305;
  wire popcount43_0kbs_core_306;
  wire popcount43_0kbs_core_307;
  wire popcount43_0kbs_core_308;
  wire popcount43_0kbs_core_310;
  wire popcount43_0kbs_core_312;
  wire popcount43_0kbs_core_313;
  wire popcount43_0kbs_core_314;
  wire popcount43_0kbs_core_315;
  wire popcount43_0kbs_core_322;
  wire popcount43_0kbs_core_324;
  wire popcount43_0kbs_core_325;
  wire popcount43_0kbs_core_326;
  wire popcount43_0kbs_core_327;
  wire popcount43_0kbs_core_330;
  wire popcount43_0kbs_core_332;
  wire popcount43_0kbs_core_334;
  wire popcount43_0kbs_core_335;
  wire popcount43_0kbs_core_337;
  wire popcount43_0kbs_core_338;
  wire popcount43_0kbs_core_339;

  assign popcount43_0kbs_core_045 = input_a[13] ^ input_a[29];
  assign popcount43_0kbs_core_049 = input_a[20] ^ input_a[19];
  assign popcount43_0kbs_core_050 = input_a[21] | input_a[8];
  assign popcount43_0kbs_core_052 = ~(input_a[18] | input_a[40]);
  assign popcount43_0kbs_core_053 = ~(input_a[13] & input_a[12]);
  assign popcount43_0kbs_core_054 = input_a[22] & input_a[39];
  assign popcount43_0kbs_core_058 = ~(input_a[8] & input_a[36]);
  assign popcount43_0kbs_core_059 = ~input_a[30];
  assign popcount43_0kbs_core_061 = ~(input_a[12] | input_a[9]);
  assign popcount43_0kbs_core_063 = input_a[11] & input_a[22];
  assign popcount43_0kbs_core_064 = ~input_a[4];
  assign popcount43_0kbs_core_069 = ~(input_a[11] ^ input_a[15]);
  assign popcount43_0kbs_core_070 = ~(input_a[38] ^ input_a[41]);
  assign popcount43_0kbs_core_074 = ~input_a[17];
  assign popcount43_0kbs_core_075 = ~(input_a[37] & input_a[1]);
  assign popcount43_0kbs_core_076 = ~(input_a[16] & input_a[39]);
  assign popcount43_0kbs_core_077 = input_a[38] ^ input_a[11];
  assign popcount43_0kbs_core_078 = input_a[14] ^ input_a[6];
  assign popcount43_0kbs_core_079 = input_a[23] & input_a[39];
  assign popcount43_0kbs_core_080 = ~input_a[26];
  assign popcount43_0kbs_core_081 = ~(input_a[12] & input_a[13]);
  assign popcount43_0kbs_core_082 = input_a[1] & input_a[26];
  assign popcount43_0kbs_core_083 = ~input_a[15];
  assign popcount43_0kbs_core_086 = ~(input_a[7] & input_a[19]);
  assign popcount43_0kbs_core_087 = ~(input_a[15] & input_a[10]);
  assign popcount43_0kbs_core_088 = ~input_a[39];
  assign popcount43_0kbs_core_089 = ~(input_a[19] & input_a[26]);
  assign popcount43_0kbs_core_090 = input_a[6] ^ input_a[40];
  assign popcount43_0kbs_core_091 = ~(input_a[32] ^ input_a[25]);
  assign popcount43_0kbs_core_092 = input_a[20] | input_a[26];
  assign popcount43_0kbs_core_093 = ~(input_a[24] ^ input_a[16]);
  assign popcount43_0kbs_core_095 = ~input_a[7];
  assign popcount43_0kbs_core_096 = ~(input_a[4] & input_a[38]);
  assign popcount43_0kbs_core_097 = input_a[20] | input_a[19];
  assign popcount43_0kbs_core_100 = ~(input_a[3] & input_a[21]);
  assign popcount43_0kbs_core_103 = ~(input_a[26] & input_a[8]);
  assign popcount43_0kbs_core_106 = ~(input_a[40] ^ input_a[32]);
  assign popcount43_0kbs_core_107 = ~(input_a[5] | input_a[9]);
  assign popcount43_0kbs_core_108 = ~input_a[2];
  assign popcount43_0kbs_core_110 = input_a[27] | input_a[1];
  assign popcount43_0kbs_core_111 = input_a[16] ^ input_a[36];
  assign popcount43_0kbs_core_112 = input_a[7] & input_a[23];
  assign popcount43_0kbs_core_114 = ~(input_a[3] & input_a[30]);
  assign popcount43_0kbs_core_116 = input_a[29] & input_a[29];
  assign popcount43_0kbs_core_117 = input_a[5] & input_a[28];
  assign popcount43_0kbs_core_118 = ~input_a[14];
  assign popcount43_0kbs_core_119 = ~input_a[11];
  assign popcount43_0kbs_core_120 = ~(input_a[7] ^ input_a[24]);
  assign popcount43_0kbs_core_125 = input_a[12] ^ input_a[22];
  assign popcount43_0kbs_core_126 = ~input_a[35];
  assign popcount43_0kbs_core_127 = input_a[32] & input_a[9];
  assign popcount43_0kbs_core_129 = ~(input_a[11] ^ input_a[17]);
  assign popcount43_0kbs_core_130 = input_a[28] & input_a[26];
  assign popcount43_0kbs_core_132 = input_a[30] ^ input_a[33];
  assign popcount43_0kbs_core_135 = ~(input_a[10] | input_a[37]);
  assign popcount43_0kbs_core_136 = ~(input_a[29] & input_a[6]);
  assign popcount43_0kbs_core_137 = input_a[24] | input_a[10];
  assign popcount43_0kbs_core_138 = input_a[33] & input_a[38];
  assign popcount43_0kbs_core_139 = input_a[21] ^ input_a[17];
  assign popcount43_0kbs_core_140 = input_a[19] | input_a[13];
  assign popcount43_0kbs_core_141 = ~(input_a[22] ^ input_a[14]);
  assign popcount43_0kbs_core_142 = ~(input_a[34] ^ input_a[36]);
  assign popcount43_0kbs_core_143 = ~(input_a[28] & input_a[19]);
  assign popcount43_0kbs_core_144 = ~(input_a[33] | input_a[41]);
  assign popcount43_0kbs_core_146 = ~(input_a[11] | input_a[36]);
  assign popcount43_0kbs_core_147 = ~(input_a[14] ^ input_a[22]);
  assign popcount43_0kbs_core_148 = ~(input_a[5] ^ input_a[41]);
  assign popcount43_0kbs_core_149 = ~(input_a[32] & input_a[32]);
  assign popcount43_0kbs_core_150_not = ~input_a[21];
  assign popcount43_0kbs_core_151 = ~(input_a[31] ^ input_a[24]);
  assign popcount43_0kbs_core_156 = ~(input_a[40] & input_a[14]);
  assign popcount43_0kbs_core_157 = input_a[9] ^ input_a[40];
  assign popcount43_0kbs_core_158 = input_a[36] ^ input_a[41];
  assign popcount43_0kbs_core_159_not = ~input_a[29];
  assign popcount43_0kbs_core_160 = ~(input_a[6] | input_a[34]);
  assign popcount43_0kbs_core_161 = ~(input_a[13] | input_a[12]);
  assign popcount43_0kbs_core_162 = input_a[20] & input_a[10];
  assign popcount43_0kbs_core_163 = input_a[25] | input_a[33];
  assign popcount43_0kbs_core_164 = ~(input_a[39] | input_a[30]);
  assign popcount43_0kbs_core_167 = ~(input_a[5] | input_a[31]);
  assign popcount43_0kbs_core_169 = ~(input_a[31] & input_a[32]);
  assign popcount43_0kbs_core_170 = input_a[14] & input_a[33];
  assign popcount43_0kbs_core_173 = ~input_a[9];
  assign popcount43_0kbs_core_174 = input_a[30] & input_a[0];
  assign popcount43_0kbs_core_175 = input_a[20] | input_a[37];
  assign popcount43_0kbs_core_176 = ~(input_a[16] & input_a[34]);
  assign popcount43_0kbs_core_177 = input_a[12] | input_a[28];
  assign popcount43_0kbs_core_178 = input_a[10] & input_a[42];
  assign popcount43_0kbs_core_179 = input_a[1] ^ input_a[19];
  assign popcount43_0kbs_core_181 = ~input_a[0];
  assign popcount43_0kbs_core_182 = input_a[25] & input_a[35];
  assign popcount43_0kbs_core_186 = input_a[10] ^ input_a[39];
  assign popcount43_0kbs_core_187 = input_a[2] & input_a[24];
  assign popcount43_0kbs_core_190 = ~(input_a[27] | input_a[36]);
  assign popcount43_0kbs_core_191 = ~(input_a[22] | input_a[24]);
  assign popcount43_0kbs_core_192 = ~(input_a[35] ^ input_a[18]);
  assign popcount43_0kbs_core_195 = ~(input_a[0] & input_a[35]);
  assign popcount43_0kbs_core_196 = ~(input_a[38] ^ input_a[15]);
  assign popcount43_0kbs_core_197 = ~(input_a[42] | input_a[20]);
  assign popcount43_0kbs_core_198 = input_a[6] & input_a[1];
  assign popcount43_0kbs_core_199 = ~(input_a[20] ^ input_a[13]);
  assign popcount43_0kbs_core_200 = input_a[35] | input_a[7];
  assign popcount43_0kbs_core_202 = input_a[20] & input_a[34];
  assign popcount43_0kbs_core_203 = ~(input_a[41] | input_a[28]);
  assign popcount43_0kbs_core_204 = input_a[39] ^ input_a[25];
  assign popcount43_0kbs_core_205 = input_a[41] & input_a[42];
  assign popcount43_0kbs_core_207 = input_a[22] & input_a[36];
  assign popcount43_0kbs_core_212 = ~input_a[16];
  assign popcount43_0kbs_core_215 = input_a[27] | input_a[39];
  assign popcount43_0kbs_core_216 = ~(input_a[15] ^ input_a[35]);
  assign popcount43_0kbs_core_218 = ~input_a[3];
  assign popcount43_0kbs_core_222 = ~(input_a[11] ^ input_a[33]);
  assign popcount43_0kbs_core_227 = input_a[18] & input_a[7];
  assign popcount43_0kbs_core_229 = input_a[4] | input_a[39];
  assign popcount43_0kbs_core_231_not = ~input_a[42];
  assign popcount43_0kbs_core_232 = input_a[5] ^ input_a[1];
  assign popcount43_0kbs_core_234 = input_a[40] | input_a[32];
  assign popcount43_0kbs_core_235 = input_a[4] & input_a[38];
  assign popcount43_0kbs_core_236 = input_a[27] | input_a[35];
  assign popcount43_0kbs_core_237 = ~(input_a[8] ^ input_a[33]);
  assign popcount43_0kbs_core_238 = input_a[23] & input_a[25];
  assign popcount43_0kbs_core_239 = ~input_a[20];
  assign popcount43_0kbs_core_240 = input_a[10] ^ input_a[14];
  assign popcount43_0kbs_core_242 = input_a[14] & input_a[41];
  assign popcount43_0kbs_core_243 = input_a[35] | input_a[8];
  assign popcount43_0kbs_core_244 = ~(input_a[30] | input_a[7]);
  assign popcount43_0kbs_core_245 = ~(input_a[35] | input_a[23]);
  assign popcount43_0kbs_core_247 = ~(input_a[42] | input_a[15]);
  assign popcount43_0kbs_core_251 = input_a[25] & input_a[25];
  assign popcount43_0kbs_core_253 = input_a[22] & input_a[12];
  assign popcount43_0kbs_core_254 = ~input_a[34];
  assign popcount43_0kbs_core_256 = ~(input_a[25] & input_a[41]);
  assign popcount43_0kbs_core_258 = ~(input_a[10] | input_a[38]);
  assign popcount43_0kbs_core_259_not = ~input_a[6];
  assign popcount43_0kbs_core_260 = input_a[39] ^ input_a[41];
  assign popcount43_0kbs_core_262 = ~(input_a[41] ^ input_a[15]);
  assign popcount43_0kbs_core_263 = ~(input_a[4] | input_a[5]);
  assign popcount43_0kbs_core_266 = input_a[24] ^ input_a[35];
  assign popcount43_0kbs_core_267 = ~(input_a[20] ^ input_a[1]);
  assign popcount43_0kbs_core_268 = input_a[2] ^ input_a[41];
  assign popcount43_0kbs_core_269 = ~input_a[0];
  assign popcount43_0kbs_core_270 = ~input_a[41];
  assign popcount43_0kbs_core_272 = ~input_a[12];
  assign popcount43_0kbs_core_275 = ~(input_a[39] ^ input_a[7]);
  assign popcount43_0kbs_core_277 = input_a[15] & input_a[25];
  assign popcount43_0kbs_core_281 = input_a[27] | input_a[38];
  assign popcount43_0kbs_core_282 = ~(input_a[18] & input_a[33]);
  assign popcount43_0kbs_core_283 = input_a[33] & input_a[4];
  assign popcount43_0kbs_core_286 = input_a[22] | input_a[20];
  assign popcount43_0kbs_core_287 = ~input_a[34];
  assign popcount43_0kbs_core_288 = ~(input_a[39] & input_a[21]);
  assign popcount43_0kbs_core_290 = ~input_a[13];
  assign popcount43_0kbs_core_292 = input_a[12] & input_a[12];
  assign popcount43_0kbs_core_294 = input_a[17] ^ input_a[25];
  assign popcount43_0kbs_core_295 = ~(input_a[38] ^ input_a[13]);
  assign popcount43_0kbs_core_297 = ~input_a[6];
  assign popcount43_0kbs_core_299 = input_a[39] ^ input_a[27];
  assign popcount43_0kbs_core_300 = ~(input_a[16] ^ input_a[7]);
  assign popcount43_0kbs_core_301_not = ~input_a[7];
  assign popcount43_0kbs_core_302 = ~(input_a[22] ^ input_a[27]);
  assign popcount43_0kbs_core_303 = input_a[9] | input_a[8];
  assign popcount43_0kbs_core_305 = input_a[39] ^ input_a[31];
  assign popcount43_0kbs_core_306 = ~(input_a[11] & input_a[25]);
  assign popcount43_0kbs_core_307 = input_a[21] ^ input_a[28];
  assign popcount43_0kbs_core_308 = ~(input_a[16] ^ input_a[2]);
  assign popcount43_0kbs_core_310 = ~(input_a[22] & input_a[23]);
  assign popcount43_0kbs_core_312 = ~(input_a[23] & input_a[28]);
  assign popcount43_0kbs_core_313 = ~(input_a[10] | input_a[7]);
  assign popcount43_0kbs_core_314 = input_a[8] & input_a[5];
  assign popcount43_0kbs_core_315 = ~(input_a[23] | input_a[40]);
  assign popcount43_0kbs_core_322 = input_a[33] ^ input_a[32];
  assign popcount43_0kbs_core_324 = input_a[0] | input_a[32];
  assign popcount43_0kbs_core_325 = ~(input_a[15] | input_a[11]);
  assign popcount43_0kbs_core_326 = ~(input_a[35] ^ input_a[18]);
  assign popcount43_0kbs_core_327 = ~(input_a[34] ^ input_a[3]);
  assign popcount43_0kbs_core_330 = input_a[14] ^ input_a[40];
  assign popcount43_0kbs_core_332 = input_a[36] | input_a[37];
  assign popcount43_0kbs_core_334 = ~input_a[6];
  assign popcount43_0kbs_core_335 = ~input_a[31];
  assign popcount43_0kbs_core_337 = ~input_a[6];
  assign popcount43_0kbs_core_338 = ~(input_a[23] ^ input_a[5]);
  assign popcount43_0kbs_core_339 = ~(input_a[21] | input_a[21]);

  assign popcount43_0kbs_out[0] = input_a[34];
  assign popcount43_0kbs_out[1] = input_a[37];
  assign popcount43_0kbs_out[2] = 1'b1;
  assign popcount43_0kbs_out[3] = 1'b0;
  assign popcount43_0kbs_out[4] = 1'b1;
  assign popcount43_0kbs_out[5] = 1'b0;
endmodule