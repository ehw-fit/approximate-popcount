// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.31592
// WCE=5.0
// EP=0.770996%
// Printed PDK parameters:
//  Area=23899409.0
//  Delay=55256672.0
//  Power=1175500.0

module popcount21_m1cq(input [20:0] input_a, output [4:0] popcount21_m1cq_out);
  wire popcount21_m1cq_core_023;
  wire popcount21_m1cq_core_024;
  wire popcount21_m1cq_core_026;
  wire popcount21_m1cq_core_028;
  wire popcount21_m1cq_core_032;
  wire popcount21_m1cq_core_033;
  wire popcount21_m1cq_core_034;
  wire popcount21_m1cq_core_041;
  wire popcount21_m1cq_core_044;
  wire popcount21_m1cq_core_047;
  wire popcount21_m1cq_core_048;
  wire popcount21_m1cq_core_049;
  wire popcount21_m1cq_core_052;
  wire popcount21_m1cq_core_053;
  wire popcount21_m1cq_core_055;
  wire popcount21_m1cq_core_056;
  wire popcount21_m1cq_core_059;
  wire popcount21_m1cq_core_060;
  wire popcount21_m1cq_core_063;
  wire popcount21_m1cq_core_064;
  wire popcount21_m1cq_core_065;
  wire popcount21_m1cq_core_070;
  wire popcount21_m1cq_core_073;
  wire popcount21_m1cq_core_075;
  wire popcount21_m1cq_core_076;
  wire popcount21_m1cq_core_077;
  wire popcount21_m1cq_core_079;
  wire popcount21_m1cq_core_080;
  wire popcount21_m1cq_core_082;
  wire popcount21_m1cq_core_083;
  wire popcount21_m1cq_core_084;
  wire popcount21_m1cq_core_085;
  wire popcount21_m1cq_core_086;
  wire popcount21_m1cq_core_087;
  wire popcount21_m1cq_core_088;
  wire popcount21_m1cq_core_090;
  wire popcount21_m1cq_core_091;
  wire popcount21_m1cq_core_092;
  wire popcount21_m1cq_core_093;
  wire popcount21_m1cq_core_094;
  wire popcount21_m1cq_core_095;
  wire popcount21_m1cq_core_096;
  wire popcount21_m1cq_core_097;
  wire popcount21_m1cq_core_098;
  wire popcount21_m1cq_core_100;
  wire popcount21_m1cq_core_101;
  wire popcount21_m1cq_core_103;
  wire popcount21_m1cq_core_105;
  wire popcount21_m1cq_core_106;
  wire popcount21_m1cq_core_107;
  wire popcount21_m1cq_core_108;
  wire popcount21_m1cq_core_109;
  wire popcount21_m1cq_core_116;
  wire popcount21_m1cq_core_117;
  wire popcount21_m1cq_core_118;
  wire popcount21_m1cq_core_119;
  wire popcount21_m1cq_core_120;
  wire popcount21_m1cq_core_121;
  wire popcount21_m1cq_core_122;
  wire popcount21_m1cq_core_123;
  wire popcount21_m1cq_core_124;
  wire popcount21_m1cq_core_125;
  wire popcount21_m1cq_core_126;
  wire popcount21_m1cq_core_130;
  wire popcount21_m1cq_core_131;
  wire popcount21_m1cq_core_132;
  wire popcount21_m1cq_core_133;
  wire popcount21_m1cq_core_134;
  wire popcount21_m1cq_core_135;
  wire popcount21_m1cq_core_138;
  wire popcount21_m1cq_core_139;
  wire popcount21_m1cq_core_140;
  wire popcount21_m1cq_core_141;
  wire popcount21_m1cq_core_142;
  wire popcount21_m1cq_core_144;
  wire popcount21_m1cq_core_145;
  wire popcount21_m1cq_core_146;
  wire popcount21_m1cq_core_147;
  wire popcount21_m1cq_core_148;
  wire popcount21_m1cq_core_149;
  wire popcount21_m1cq_core_153;

  assign popcount21_m1cq_core_023 = input_a[17] & input_a[6];
  assign popcount21_m1cq_core_024 = ~(input_a[17] & input_a[1]);
  assign popcount21_m1cq_core_026 = input_a[3] & input_a[4];
  assign popcount21_m1cq_core_028 = input_a[8] & input_a[10];
  assign popcount21_m1cq_core_032 = ~input_a[9];
  assign popcount21_m1cq_core_033 = ~input_a[8];
  assign popcount21_m1cq_core_034 = input_a[1] & popcount21_m1cq_core_026;
  assign popcount21_m1cq_core_041 = input_a[14] & input_a[11];
  assign popcount21_m1cq_core_044 = input_a[0] & input_a[8];
  assign popcount21_m1cq_core_047 = input_a[5] | input_a[6];
  assign popcount21_m1cq_core_048 = input_a[8] ^ input_a[17];
  assign popcount21_m1cq_core_049 = ~(input_a[17] & input_a[9]);
  assign popcount21_m1cq_core_052 = input_a[11] | input_a[11];
  assign popcount21_m1cq_core_053 = input_a[13] ^ input_a[4];
  assign popcount21_m1cq_core_055 = ~input_a[5];
  assign popcount21_m1cq_core_056 = input_a[13] ^ input_a[14];
  assign popcount21_m1cq_core_059 = ~input_a[5];
  assign popcount21_m1cq_core_060 = ~(input_a[16] ^ input_a[19]);
  assign popcount21_m1cq_core_063 = input_a[0] & input_a[7];
  assign popcount21_m1cq_core_064 = ~(popcount21_m1cq_core_034 & input_a[6]);
  assign popcount21_m1cq_core_065 = popcount21_m1cq_core_034 & input_a[6];
  assign popcount21_m1cq_core_070 = ~input_a[18];
  assign popcount21_m1cq_core_073 = ~(input_a[1] | input_a[5]);
  assign popcount21_m1cq_core_075 = input_a[10] & input_a[2];
  assign popcount21_m1cq_core_076 = input_a[13] | input_a[14];
  assign popcount21_m1cq_core_077 = input_a[13] & input_a[14];
  assign popcount21_m1cq_core_079 = input_a[12] & popcount21_m1cq_core_076;
  assign popcount21_m1cq_core_080 = popcount21_m1cq_core_077 | popcount21_m1cq_core_079;
  assign popcount21_m1cq_core_082 = ~(input_a[16] ^ input_a[20]);
  assign popcount21_m1cq_core_083 = input_a[11] & input_a[7];
  assign popcount21_m1cq_core_084 = popcount21_m1cq_core_075 ^ popcount21_m1cq_core_080;
  assign popcount21_m1cq_core_085 = popcount21_m1cq_core_075 & popcount21_m1cq_core_080;
  assign popcount21_m1cq_core_086 = popcount21_m1cq_core_084 ^ popcount21_m1cq_core_083;
  assign popcount21_m1cq_core_087 = popcount21_m1cq_core_084 & popcount21_m1cq_core_083;
  assign popcount21_m1cq_core_088 = popcount21_m1cq_core_085 | popcount21_m1cq_core_087;
  assign popcount21_m1cq_core_090 = ~(input_a[16] & input_a[17]);
  assign popcount21_m1cq_core_091 = input_a[16] ^ input_a[17];
  assign popcount21_m1cq_core_092 = input_a[16] & input_a[17];
  assign popcount21_m1cq_core_093 = input_a[15] ^ popcount21_m1cq_core_091;
  assign popcount21_m1cq_core_094 = input_a[15] & popcount21_m1cq_core_091;
  assign popcount21_m1cq_core_095 = popcount21_m1cq_core_092 | popcount21_m1cq_core_094;
  assign popcount21_m1cq_core_096 = ~(input_a[8] & input_a[10]);
  assign popcount21_m1cq_core_097 = ~(input_a[8] | input_a[0]);
  assign popcount21_m1cq_core_098 = input_a[19] & input_a[20];
  assign popcount21_m1cq_core_100 = input_a[8] & input_a[18];
  assign popcount21_m1cq_core_101 = popcount21_m1cq_core_098 | popcount21_m1cq_core_100;
  assign popcount21_m1cq_core_103 = ~(input_a[6] ^ input_a[20]);
  assign popcount21_m1cq_core_105 = popcount21_m1cq_core_095 ^ popcount21_m1cq_core_101;
  assign popcount21_m1cq_core_106 = popcount21_m1cq_core_095 & popcount21_m1cq_core_101;
  assign popcount21_m1cq_core_107 = popcount21_m1cq_core_105 ^ popcount21_m1cq_core_093;
  assign popcount21_m1cq_core_108 = popcount21_m1cq_core_105 & popcount21_m1cq_core_093;
  assign popcount21_m1cq_core_109 = popcount21_m1cq_core_106 | popcount21_m1cq_core_108;
  assign popcount21_m1cq_core_116 = input_a[0] & input_a[9];
  assign popcount21_m1cq_core_117 = popcount21_m1cq_core_086 ^ popcount21_m1cq_core_107;
  assign popcount21_m1cq_core_118 = popcount21_m1cq_core_086 & popcount21_m1cq_core_107;
  assign popcount21_m1cq_core_119 = popcount21_m1cq_core_117 ^ popcount21_m1cq_core_116;
  assign popcount21_m1cq_core_120 = popcount21_m1cq_core_117 & popcount21_m1cq_core_116;
  assign popcount21_m1cq_core_121 = popcount21_m1cq_core_118 | popcount21_m1cq_core_120;
  assign popcount21_m1cq_core_122 = popcount21_m1cq_core_088 ^ popcount21_m1cq_core_109;
  assign popcount21_m1cq_core_123 = popcount21_m1cq_core_088 & popcount21_m1cq_core_109;
  assign popcount21_m1cq_core_124 = popcount21_m1cq_core_122 ^ popcount21_m1cq_core_121;
  assign popcount21_m1cq_core_125 = popcount21_m1cq_core_122 & popcount21_m1cq_core_121;
  assign popcount21_m1cq_core_126 = popcount21_m1cq_core_123 | popcount21_m1cq_core_125;
  assign popcount21_m1cq_core_130 = ~(input_a[14] & input_a[15]);
  assign popcount21_m1cq_core_131 = ~(input_a[18] ^ input_a[10]);
  assign popcount21_m1cq_core_132 = ~(input_a[20] | input_a[6]);
  assign popcount21_m1cq_core_133 = ~(input_a[11] ^ input_a[17]);
  assign popcount21_m1cq_core_134 = input_a[19] | input_a[20];
  assign popcount21_m1cq_core_135 = input_a[15] ^ input_a[0];
  assign popcount21_m1cq_core_138 = input_a[15] & input_a[2];
  assign popcount21_m1cq_core_139 = popcount21_m1cq_core_064 ^ popcount21_m1cq_core_124;
  assign popcount21_m1cq_core_140 = popcount21_m1cq_core_064 & popcount21_m1cq_core_124;
  assign popcount21_m1cq_core_141 = input_a[0] | input_a[14];
  assign popcount21_m1cq_core_142 = input_a[18] | input_a[12];
  assign popcount21_m1cq_core_144 = popcount21_m1cq_core_065 ^ popcount21_m1cq_core_126;
  assign popcount21_m1cq_core_145 = popcount21_m1cq_core_065 & popcount21_m1cq_core_126;
  assign popcount21_m1cq_core_146 = popcount21_m1cq_core_144 ^ popcount21_m1cq_core_140;
  assign popcount21_m1cq_core_147 = popcount21_m1cq_core_144 & popcount21_m1cq_core_140;
  assign popcount21_m1cq_core_148 = popcount21_m1cq_core_145 | popcount21_m1cq_core_147;
  assign popcount21_m1cq_core_149 = ~(input_a[9] & input_a[9]);
  assign popcount21_m1cq_core_153 = ~(input_a[9] | input_a[10]);

  assign popcount21_m1cq_out[0] = input_a[5];
  assign popcount21_m1cq_out[1] = popcount21_m1cq_core_119;
  assign popcount21_m1cq_out[2] = popcount21_m1cq_core_139;
  assign popcount21_m1cq_out[3] = popcount21_m1cq_core_146;
  assign popcount21_m1cq_out[4] = popcount21_m1cq_core_148;
endmodule