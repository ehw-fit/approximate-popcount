// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.18645
// WCE=12.0
// EP=0.859843%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount22_y1dy(input [21:0] input_a, output [4:0] popcount22_y1dy_out);
  wire popcount22_y1dy_core_025;
  wire popcount22_y1dy_core_027;
  wire popcount22_y1dy_core_029;
  wire popcount22_y1dy_core_031;
  wire popcount22_y1dy_core_032;
  wire popcount22_y1dy_core_033;
  wire popcount22_y1dy_core_034;
  wire popcount22_y1dy_core_035;
  wire popcount22_y1dy_core_037;
  wire popcount22_y1dy_core_038;
  wire popcount22_y1dy_core_040;
  wire popcount22_y1dy_core_041;
  wire popcount22_y1dy_core_042;
  wire popcount22_y1dy_core_043;
  wire popcount22_y1dy_core_045;
  wire popcount22_y1dy_core_048;
  wire popcount22_y1dy_core_049;
  wire popcount22_y1dy_core_051;
  wire popcount22_y1dy_core_052;
  wire popcount22_y1dy_core_053;
  wire popcount22_y1dy_core_055;
  wire popcount22_y1dy_core_057;
  wire popcount22_y1dy_core_059;
  wire popcount22_y1dy_core_061;
  wire popcount22_y1dy_core_062;
  wire popcount22_y1dy_core_063;
  wire popcount22_y1dy_core_064;
  wire popcount22_y1dy_core_065;
  wire popcount22_y1dy_core_067;
  wire popcount22_y1dy_core_070;
  wire popcount22_y1dy_core_072;
  wire popcount22_y1dy_core_075;
  wire popcount22_y1dy_core_076;
  wire popcount22_y1dy_core_077;
  wire popcount22_y1dy_core_081;
  wire popcount22_y1dy_core_083;
  wire popcount22_y1dy_core_084;
  wire popcount22_y1dy_core_087;
  wire popcount22_y1dy_core_088;
  wire popcount22_y1dy_core_089;
  wire popcount22_y1dy_core_091;
  wire popcount22_y1dy_core_092;
  wire popcount22_y1dy_core_093;
  wire popcount22_y1dy_core_096;
  wire popcount22_y1dy_core_098_not;
  wire popcount22_y1dy_core_101;
  wire popcount22_y1dy_core_103_not;
  wire popcount22_y1dy_core_104;
  wire popcount22_y1dy_core_105;
  wire popcount22_y1dy_core_106;
  wire popcount22_y1dy_core_109;
  wire popcount22_y1dy_core_112;
  wire popcount22_y1dy_core_115;
  wire popcount22_y1dy_core_116;
  wire popcount22_y1dy_core_118;
  wire popcount22_y1dy_core_119;
  wire popcount22_y1dy_core_120;
  wire popcount22_y1dy_core_123;
  wire popcount22_y1dy_core_125_not;
  wire popcount22_y1dy_core_126;
  wire popcount22_y1dy_core_129;
  wire popcount22_y1dy_core_130;
  wire popcount22_y1dy_core_132;
  wire popcount22_y1dy_core_133;
  wire popcount22_y1dy_core_139;
  wire popcount22_y1dy_core_141;
  wire popcount22_y1dy_core_142;
  wire popcount22_y1dy_core_143_not;
  wire popcount22_y1dy_core_144;
  wire popcount22_y1dy_core_145;
  wire popcount22_y1dy_core_151;
  wire popcount22_y1dy_core_152;
  wire popcount22_y1dy_core_153;
  wire popcount22_y1dy_core_154;
  wire popcount22_y1dy_core_155;
  wire popcount22_y1dy_core_157;
  wire popcount22_y1dy_core_158_not;
  wire popcount22_y1dy_core_161;

  assign popcount22_y1dy_core_025 = ~input_a[5];
  assign popcount22_y1dy_core_027 = ~(input_a[20] | input_a[10]);
  assign popcount22_y1dy_core_029 = input_a[9] ^ input_a[19];
  assign popcount22_y1dy_core_031 = input_a[2] ^ input_a[11];
  assign popcount22_y1dy_core_032 = input_a[11] | input_a[4];
  assign popcount22_y1dy_core_033 = ~input_a[21];
  assign popcount22_y1dy_core_034 = ~(input_a[4] ^ input_a[5]);
  assign popcount22_y1dy_core_035 = input_a[4] & input_a[21];
  assign popcount22_y1dy_core_037 = ~(input_a[4] & input_a[17]);
  assign popcount22_y1dy_core_038 = input_a[1] | input_a[5];
  assign popcount22_y1dy_core_040 = ~input_a[4];
  assign popcount22_y1dy_core_041 = input_a[10] | input_a[18];
  assign popcount22_y1dy_core_042 = ~(input_a[13] & input_a[20]);
  assign popcount22_y1dy_core_043 = ~(input_a[6] ^ input_a[0]);
  assign popcount22_y1dy_core_045 = ~(input_a[15] ^ input_a[1]);
  assign popcount22_y1dy_core_048 = ~(input_a[6] & input_a[9]);
  assign popcount22_y1dy_core_049 = ~input_a[8];
  assign popcount22_y1dy_core_051 = ~input_a[14];
  assign popcount22_y1dy_core_052 = input_a[20] ^ input_a[1];
  assign popcount22_y1dy_core_053 = ~(input_a[11] | input_a[15]);
  assign popcount22_y1dy_core_055 = ~input_a[5];
  assign popcount22_y1dy_core_057 = input_a[8] | input_a[6];
  assign popcount22_y1dy_core_059 = input_a[16] ^ input_a[10];
  assign popcount22_y1dy_core_061 = ~(input_a[14] ^ input_a[14]);
  assign popcount22_y1dy_core_062 = input_a[5] | input_a[2];
  assign popcount22_y1dy_core_063 = input_a[20] & input_a[11];
  assign popcount22_y1dy_core_064 = input_a[4] & input_a[15];
  assign popcount22_y1dy_core_065 = input_a[2] & input_a[1];
  assign popcount22_y1dy_core_067 = input_a[17] & input_a[13];
  assign popcount22_y1dy_core_070 = ~(input_a[11] | input_a[21]);
  assign popcount22_y1dy_core_072 = ~input_a[3];
  assign popcount22_y1dy_core_075 = input_a[0] & input_a[7];
  assign popcount22_y1dy_core_076 = input_a[10] & input_a[9];
  assign popcount22_y1dy_core_077 = input_a[4] | input_a[6];
  assign popcount22_y1dy_core_081 = input_a[13] ^ input_a[14];
  assign popcount22_y1dy_core_083 = input_a[8] & input_a[15];
  assign popcount22_y1dy_core_084 = ~(input_a[3] | input_a[7]);
  assign popcount22_y1dy_core_087 = input_a[5] & input_a[1];
  assign popcount22_y1dy_core_088 = ~(input_a[10] & input_a[14]);
  assign popcount22_y1dy_core_089 = input_a[14] | input_a[15];
  assign popcount22_y1dy_core_091 = ~input_a[8];
  assign popcount22_y1dy_core_092 = input_a[3] & input_a[10];
  assign popcount22_y1dy_core_093 = input_a[10] ^ input_a[11];
  assign popcount22_y1dy_core_096 = ~(input_a[10] | input_a[1]);
  assign popcount22_y1dy_core_098_not = ~input_a[18];
  assign popcount22_y1dy_core_101 = input_a[15] ^ input_a[13];
  assign popcount22_y1dy_core_103_not = ~input_a[4];
  assign popcount22_y1dy_core_104 = input_a[6] ^ input_a[11];
  assign popcount22_y1dy_core_105 = ~(input_a[2] | input_a[10]);
  assign popcount22_y1dy_core_106 = ~(input_a[4] & input_a[15]);
  assign popcount22_y1dy_core_109 = ~input_a[11];
  assign popcount22_y1dy_core_112 = ~(input_a[15] & input_a[11]);
  assign popcount22_y1dy_core_115 = ~(input_a[19] & input_a[18]);
  assign popcount22_y1dy_core_116 = ~input_a[12];
  assign popcount22_y1dy_core_118 = input_a[12] ^ input_a[2];
  assign popcount22_y1dy_core_119 = input_a[1] ^ input_a[1];
  assign popcount22_y1dy_core_120 = input_a[9] | input_a[9];
  assign popcount22_y1dy_core_123 = ~(input_a[11] ^ input_a[8]);
  assign popcount22_y1dy_core_125_not = ~input_a[7];
  assign popcount22_y1dy_core_126 = input_a[0] | input_a[5];
  assign popcount22_y1dy_core_129 = ~(input_a[9] ^ input_a[9]);
  assign popcount22_y1dy_core_130 = input_a[3] | input_a[16];
  assign popcount22_y1dy_core_132 = input_a[12] | input_a[11];
  assign popcount22_y1dy_core_133 = ~(input_a[15] & input_a[13]);
  assign popcount22_y1dy_core_139 = input_a[18] ^ input_a[8];
  assign popcount22_y1dy_core_141 = ~(input_a[16] | input_a[15]);
  assign popcount22_y1dy_core_142 = ~(input_a[13] & input_a[3]);
  assign popcount22_y1dy_core_143_not = ~input_a[15];
  assign popcount22_y1dy_core_144 = input_a[4] ^ input_a[18];
  assign popcount22_y1dy_core_145 = ~(input_a[17] & input_a[7]);
  assign popcount22_y1dy_core_151 = ~(input_a[17] & input_a[3]);
  assign popcount22_y1dy_core_152 = ~input_a[13];
  assign popcount22_y1dy_core_153 = ~input_a[6];
  assign popcount22_y1dy_core_154 = ~input_a[2];
  assign popcount22_y1dy_core_155 = ~(input_a[4] | input_a[13]);
  assign popcount22_y1dy_core_157 = ~(input_a[12] | input_a[13]);
  assign popcount22_y1dy_core_158_not = ~input_a[21];
  assign popcount22_y1dy_core_161 = input_a[18] & input_a[3];

  assign popcount22_y1dy_out[0] = input_a[10];
  assign popcount22_y1dy_out[1] = input_a[15];
  assign popcount22_y1dy_out[2] = input_a[0];
  assign popcount22_y1dy_out[3] = 1'b1;
  assign popcount22_y1dy_out[4] = 1'b0;
endmodule