
module cmp_pos(input [59:0] input_a, output [5:0] cgp_out);
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_111;
  wire cgp_core_113;
  wire cgp_core_114;
  wire cgp_core_115;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_118;
  wire cgp_core_119;
  wire cgp_core_120;
  wire cgp_core_121;
  wire cgp_core_122;
  wire cgp_core_123;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_129;
  wire cgp_core_130;
  wire cgp_core_131;
  wire cgp_core_132;
  wire cgp_core_133;
  wire cgp_core_134;
  wire cgp_core_135;
  wire cgp_core_136;
  wire cgp_core_138;
  wire cgp_core_139;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_146;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_150;
  wire cgp_core_151;
  wire cgp_core_152;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_161;
  wire cgp_core_162;
  wire cgp_core_163;
  wire cgp_core_164;
  wire cgp_core_165;
  wire cgp_core_168;
  wire cgp_core_169;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_188;
  wire cgp_core_189;
  wire cgp_core_190;
  wire cgp_core_191;
  wire cgp_core_193;
  wire cgp_core_194;
  wire cgp_core_195;
  wire cgp_core_196;
  wire cgp_core_197;
  wire cgp_core_198;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_205;
  wire cgp_core_206;
  wire cgp_core_207;
  wire cgp_core_208;
  wire cgp_core_209;
  wire cgp_core_210;
  wire cgp_core_211;
  wire cgp_core_212;
  wire cgp_core_213;
  wire cgp_core_214;
  wire cgp_core_215;
  wire cgp_core_216;
  wire cgp_core_219;
  wire cgp_core_220;
  wire cgp_core_221;
  wire cgp_core_222;
  wire cgp_core_223;
  wire cgp_core_224;
  wire cgp_core_225;
  wire cgp_core_226;
  wire cgp_core_227;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_230;
  wire cgp_core_231;
  wire cgp_core_232;
  wire cgp_core_233;
  wire cgp_core_234;
  wire cgp_core_235;
  wire cgp_core_236;
  wire cgp_core_237;
  wire cgp_core_238;
  wire cgp_core_240;
  wire cgp_core_242;
  wire cgp_core_243;
  wire cgp_core_244;
  wire cgp_core_245;
  wire cgp_core_246;
  wire cgp_core_247;
  wire cgp_core_248;
  wire cgp_core_250;
  wire cgp_core_251;
  wire cgp_core_252;
  wire cgp_core_253;
  wire cgp_core_254;
  wire cgp_core_255;
  wire cgp_core_256;
  wire cgp_core_257;
  wire cgp_core_258;
  wire cgp_core_261;
  wire cgp_core_262;
  wire cgp_core_263;
  wire cgp_core_264;
  wire cgp_core_265;
  wire cgp_core_266;
  wire cgp_core_267;
  wire cgp_core_269;
  wire cgp_core_270;
  wire cgp_core_271;
  wire cgp_core_273;
  wire cgp_core_274;
  wire cgp_core_275;
  wire cgp_core_276;
  wire cgp_core_277;
  wire cgp_core_278;
  wire cgp_core_279;
  wire cgp_core_280;
  wire cgp_core_281;
  wire cgp_core_282;
  wire cgp_core_284;
  wire cgp_core_285;
  wire cgp_core_286;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_290;
  wire cgp_core_291;
  wire cgp_core_292;
  wire cgp_core_293;
  wire cgp_core_295;
  wire cgp_core_296;
  wire cgp_core_297;
  wire cgp_core_298;
  wire cgp_core_299;
  wire cgp_core_300;
  wire cgp_core_301;
  wire cgp_core_302;
  wire cgp_core_303;
  wire cgp_core_304;
  wire cgp_core_307;
  wire cgp_core_308;
  wire cgp_core_309;
  wire cgp_core_310;
  wire cgp_core_311;
  wire cgp_core_312;
  wire cgp_core_313;
  wire cgp_core_314;
  wire cgp_core_315;
  wire cgp_core_316;
  wire cgp_core_317;
  wire cgp_core_318;
  wire cgp_core_320;
  wire cgp_core_321;
  wire cgp_core_323;
  wire cgp_core_324;
  wire cgp_core_325;
  wire cgp_core_326;
  wire cgp_core_327;
  wire cgp_core_328;
  wire cgp_core_330;
  wire cgp_core_331;
  wire cgp_core_332;
  wire cgp_core_333;
  wire cgp_core_334;
  wire cgp_core_335;
  wire cgp_core_336;
  wire cgp_core_337;
  wire cgp_core_338;
  wire cgp_core_341;
  wire cgp_core_342;
  wire cgp_core_343;
  wire cgp_core_344;
  wire cgp_core_345;
  wire cgp_core_346;
  wire cgp_core_347;
  wire cgp_core_349;
  wire cgp_core_350;
  wire cgp_core_353;
  wire cgp_core_354;
  wire cgp_core_355;
  wire cgp_core_356;
  wire cgp_core_357;
  wire cgp_core_358;
  wire cgp_core_359;
  wire cgp_core_360;
  wire cgp_core_361;
  wire cgp_core_362;
  wire cgp_core_364;
  wire cgp_core_365;
  wire cgp_core_366;
  wire cgp_core_367;
  wire cgp_core_368;
  wire cgp_core_369;
  wire cgp_core_370;
  wire cgp_core_371;
  wire cgp_core_372;
  wire cgp_core_373;
  wire cgp_core_375;
  wire cgp_core_376;
  wire cgp_core_377;
  wire cgp_core_378;
  wire cgp_core_379;
  wire cgp_core_380;
  wire cgp_core_381;
  wire cgp_core_382;
  wire cgp_core_383;
  wire cgp_core_384;
  wire cgp_core_385;
  wire cgp_core_387;
  wire cgp_core_388;
  wire cgp_core_389;
  wire cgp_core_390;
  wire cgp_core_391;
  wire cgp_core_392;
  wire cgp_core_393;
  wire cgp_core_394;
  wire cgp_core_395;
  wire cgp_core_396;
  wire cgp_core_397;
  wire cgp_core_398;
  wire cgp_core_400;
  wire cgp_core_401;
  wire cgp_core_403;
  wire cgp_core_404;
  wire cgp_core_405;
  wire cgp_core_406;
  wire cgp_core_407;
  wire cgp_core_408;
  wire cgp_core_409;
  wire cgp_core_410;
  wire cgp_core_411;
  wire cgp_core_412;
  wire cgp_core_413;
  wire cgp_core_414;
  wire cgp_core_415;
  wire cgp_core_416;
  wire cgp_core_417;
  wire cgp_core_418;
  wire cgp_core_419;
  wire cgp_core_420;
  wire cgp_core_422;
  wire cgp_core_424;
  wire cgp_core_426;
  wire cgp_core_427;
  wire cgp_core_428;
  wire cgp_core_429;
  wire cgp_core_430;
  wire cgp_core_431;
  wire cgp_core_432;
  wire cgp_core_433;
  wire cgp_core_434;
  wire cgp_core_435;
  wire cgp_core_436;
  wire cgp_core_437;
  wire cgp_core_438;
  wire cgp_core_439;
  wire cgp_core_440;
  wire cgp_core_441;
  wire cgp_core_442;
  wire cgp_core_443;
  wire cgp_core_444;
  wire cgp_core_445;
  wire cgp_core_446;
  wire cgp_core_447;
  wire cgp_core_448;
  wire cgp_core_449;
  wire cgp_core_450;
  wire cgp_core_452;

  assign cgp_core_062 = input_a[1] ^ input_a[2];
  assign cgp_core_063 = input_a[1] & input_a[2];
  assign cgp_core_064 = input_a[0] ^ cgp_core_062;
  assign cgp_core_065 = input_a[0] & cgp_core_062;
  assign cgp_core_066 = cgp_core_063 | cgp_core_065;
  assign cgp_core_068 = input_a[3] ^ input_a[4];
  assign cgp_core_069 = input_a[3] & input_a[4];
  assign cgp_core_070 = input_a[5] ^ input_a[6];
  assign cgp_core_071 = input_a[5] & input_a[6];
  assign cgp_core_072 = cgp_core_068 ^ cgp_core_070;
  assign cgp_core_073 = cgp_core_068 & cgp_core_070;
  assign cgp_core_074 = cgp_core_069 ^ cgp_core_071;
  assign cgp_core_075 = cgp_core_069 & cgp_core_071;
  assign cgp_core_076 = cgp_core_074 | cgp_core_073;
  assign cgp_core_077 = input_a[53] ^ input_a[39];
  assign cgp_core_079 = cgp_core_064 ^ cgp_core_072;
  assign cgp_core_080 = cgp_core_064 & cgp_core_072;
  assign cgp_core_081 = cgp_core_066 ^ cgp_core_076;
  assign cgp_core_082 = cgp_core_066 & cgp_core_076;
  assign cgp_core_083 = cgp_core_081 ^ cgp_core_080;
  assign cgp_core_084 = cgp_core_081 & cgp_core_080;
  assign cgp_core_085 = cgp_core_082 | cgp_core_084;
  assign cgp_core_087 = input_a[30] ^ input_a[46];
  assign cgp_core_088 = cgp_core_075 | cgp_core_085;
  assign cgp_core_089 = ~(input_a[14] ^ input_a[31]);
  assign cgp_core_091 = input_a[7] ^ input_a[8];
  assign cgp_core_092 = input_a[7] & input_a[8];
  assign cgp_core_093 = input_a[9] ^ input_a[10];
  assign cgp_core_094 = input_a[9] & input_a[10];
  assign cgp_core_095 = cgp_core_091 ^ cgp_core_093;
  assign cgp_core_096 = cgp_core_091 & cgp_core_093;
  assign cgp_core_097 = cgp_core_092 ^ cgp_core_094;
  assign cgp_core_098 = cgp_core_092 & cgp_core_094;
  assign cgp_core_099 = cgp_core_097 | cgp_core_096;
  assign cgp_core_100 = ~(input_a[52] & input_a[0]);
  assign cgp_core_102 = input_a[11] ^ input_a[12];
  assign cgp_core_103 = input_a[11] & input_a[12];
  assign cgp_core_104 = input_a[13] ^ input_a[14];
  assign cgp_core_105 = input_a[13] & input_a[14];
  assign cgp_core_106 = cgp_core_102 ^ cgp_core_104;
  assign cgp_core_107 = cgp_core_102 & cgp_core_104;
  assign cgp_core_108 = cgp_core_103 ^ cgp_core_105;
  assign cgp_core_109 = cgp_core_103 & cgp_core_105;
  assign cgp_core_110 = cgp_core_108 | cgp_core_107;
  assign cgp_core_111 = ~(input_a[25] | input_a[54]);
  assign cgp_core_113 = cgp_core_095 ^ cgp_core_106;
  assign cgp_core_114 = cgp_core_095 & cgp_core_106;
  assign cgp_core_115 = cgp_core_099 ^ cgp_core_110;
  assign cgp_core_116 = cgp_core_099 & cgp_core_110;
  assign cgp_core_117 = cgp_core_115 ^ cgp_core_114;
  assign cgp_core_118 = cgp_core_115 & cgp_core_114;
  assign cgp_core_119 = cgp_core_116 | cgp_core_118;
  assign cgp_core_120 = cgp_core_098 ^ cgp_core_109;
  assign cgp_core_121 = cgp_core_098 & cgp_core_109;
  assign cgp_core_122 = cgp_core_120 | cgp_core_119;
  assign cgp_core_123 = input_a[4] ^ input_a[32];
  assign cgp_core_125 = cgp_core_079 ^ cgp_core_113;
  assign cgp_core_126 = cgp_core_079 & cgp_core_113;
  assign cgp_core_127 = cgp_core_083 ^ cgp_core_117;
  assign cgp_core_128 = cgp_core_083 & cgp_core_117;
  assign cgp_core_129 = cgp_core_127 ^ cgp_core_126;
  assign cgp_core_130 = cgp_core_127 & cgp_core_126;
  assign cgp_core_131 = cgp_core_128 | cgp_core_130;
  assign cgp_core_132 = cgp_core_088 ^ cgp_core_122;
  assign cgp_core_133 = cgp_core_088 & cgp_core_122;
  assign cgp_core_134 = cgp_core_132 ^ cgp_core_131;
  assign cgp_core_135 = cgp_core_132 & cgp_core_131;
  assign cgp_core_136 = cgp_core_133 | cgp_core_135;
  assign cgp_core_138 = ~input_a[45];
  assign cgp_core_139 = cgp_core_121 | cgp_core_136;
  assign cgp_core_141 = ~(input_a[24] ^ input_a[38]);
  assign cgp_core_142 = input_a[16] ^ input_a[17];
  assign cgp_core_143 = input_a[16] & input_a[17];
  assign cgp_core_144 = input_a[15] ^ cgp_core_142;
  assign cgp_core_145 = input_a[15] & cgp_core_142;
  assign cgp_core_146 = cgp_core_143 | cgp_core_145;
  assign cgp_core_148 = input_a[18] ^ input_a[19];
  assign cgp_core_149 = input_a[18] & input_a[19];
  assign cgp_core_150 = input_a[20] ^ input_a[21];
  assign cgp_core_151 = input_a[20] & input_a[21];
  assign cgp_core_152 = cgp_core_148 ^ cgp_core_150;
  assign cgp_core_153 = cgp_core_148 & cgp_core_150;
  assign cgp_core_154 = cgp_core_149 ^ cgp_core_151;
  assign cgp_core_155 = cgp_core_149 & cgp_core_151;
  assign cgp_core_156 = cgp_core_154 | cgp_core_153;
  assign cgp_core_157 = ~(input_a[48] & input_a[51]);
  assign cgp_core_159 = cgp_core_144 ^ cgp_core_152;
  assign cgp_core_160 = cgp_core_144 & cgp_core_152;
  assign cgp_core_161 = cgp_core_146 ^ cgp_core_156;
  assign cgp_core_162 = cgp_core_146 & cgp_core_156;
  assign cgp_core_163 = cgp_core_161 ^ cgp_core_160;
  assign cgp_core_164 = cgp_core_161 & cgp_core_160;
  assign cgp_core_165 = cgp_core_162 | cgp_core_164;
  assign cgp_core_168 = cgp_core_155 | cgp_core_165;
  assign cgp_core_169 = input_a[30] | input_a[32];
  assign cgp_core_171 = input_a[22] ^ input_a[23];
  assign cgp_core_172 = input_a[22] & input_a[23];
  assign cgp_core_173 = input_a[24] ^ input_a[25];
  assign cgp_core_174 = input_a[24] & input_a[25];
  assign cgp_core_175 = cgp_core_171 ^ cgp_core_173;
  assign cgp_core_176 = cgp_core_171 & cgp_core_173;
  assign cgp_core_177 = cgp_core_172 ^ cgp_core_174;
  assign cgp_core_178 = cgp_core_172 & cgp_core_174;
  assign cgp_core_179 = cgp_core_177 | cgp_core_176;
  assign cgp_core_182 = input_a[26] ^ input_a[27];
  assign cgp_core_183 = input_a[26] & input_a[27];
  assign cgp_core_184 = input_a[28] ^ input_a[29];
  assign cgp_core_185 = input_a[28] & input_a[29];
  assign cgp_core_186 = cgp_core_182 ^ cgp_core_184;
  assign cgp_core_187 = cgp_core_182 & cgp_core_184;
  assign cgp_core_188 = cgp_core_183 ^ cgp_core_185;
  assign cgp_core_189 = cgp_core_183 & cgp_core_185;
  assign cgp_core_190 = cgp_core_188 | cgp_core_187;
  assign cgp_core_191 = ~input_a[9];
  assign cgp_core_193 = cgp_core_175 ^ cgp_core_186;
  assign cgp_core_194 = cgp_core_175 & cgp_core_186;
  assign cgp_core_195 = cgp_core_179 ^ cgp_core_190;
  assign cgp_core_196 = cgp_core_179 & cgp_core_190;
  assign cgp_core_197 = cgp_core_195 ^ cgp_core_194;
  assign cgp_core_198 = cgp_core_195 & cgp_core_194;
  assign cgp_core_199 = cgp_core_196 | cgp_core_198;
  assign cgp_core_200 = cgp_core_178 ^ cgp_core_189;
  assign cgp_core_201 = cgp_core_178 & cgp_core_189;
  assign cgp_core_202 = cgp_core_200 | cgp_core_199;
  assign cgp_core_205 = cgp_core_159 ^ cgp_core_193;
  assign cgp_core_206 = cgp_core_159 & cgp_core_193;
  assign cgp_core_207 = cgp_core_163 ^ cgp_core_197;
  assign cgp_core_208 = cgp_core_163 & cgp_core_197;
  assign cgp_core_209 = cgp_core_207 ^ cgp_core_206;
  assign cgp_core_210 = cgp_core_207 & cgp_core_206;
  assign cgp_core_211 = cgp_core_208 | cgp_core_210;
  assign cgp_core_212 = cgp_core_168 ^ cgp_core_202;
  assign cgp_core_213 = cgp_core_168 & cgp_core_202;
  assign cgp_core_214 = cgp_core_212 ^ cgp_core_211;
  assign cgp_core_215 = cgp_core_212 & cgp_core_211;
  assign cgp_core_216 = cgp_core_213 | cgp_core_215;
  assign cgp_core_219 = cgp_core_201 | cgp_core_216;
  assign cgp_core_220 = input_a[44] | input_a[53];
  assign cgp_core_221 = ~(input_a[56] & input_a[47]);
  assign cgp_core_222 = cgp_core_125 ^ cgp_core_205;
  assign cgp_core_223 = cgp_core_125 & cgp_core_205;
  assign cgp_core_224 = cgp_core_129 ^ cgp_core_209;
  assign cgp_core_225 = cgp_core_129 & cgp_core_209;
  assign cgp_core_226 = cgp_core_224 ^ cgp_core_223;
  assign cgp_core_227 = cgp_core_224 & cgp_core_223;
  assign cgp_core_228 = cgp_core_225 | cgp_core_227;
  assign cgp_core_229 = cgp_core_134 ^ cgp_core_214;
  assign cgp_core_230 = cgp_core_134 & cgp_core_214;
  assign cgp_core_231 = cgp_core_229 ^ cgp_core_228;
  assign cgp_core_232 = cgp_core_229 & cgp_core_228;
  assign cgp_core_233 = cgp_core_230 | cgp_core_232;
  assign cgp_core_234 = cgp_core_139 ^ cgp_core_219;
  assign cgp_core_235 = cgp_core_139 & cgp_core_219;
  assign cgp_core_236 = cgp_core_234 ^ cgp_core_233;
  assign cgp_core_237 = cgp_core_234 & cgp_core_233;
  assign cgp_core_238 = cgp_core_235 | cgp_core_237;
  assign cgp_core_240 = input_a[29] | input_a[48];
  assign cgp_core_242 = input_a[34] | input_a[57];
  assign cgp_core_243 = ~(input_a[4] & input_a[45]);
  assign cgp_core_244 = input_a[31] ^ input_a[32];
  assign cgp_core_245 = input_a[31] & input_a[32];
  assign cgp_core_246 = input_a[30] ^ cgp_core_244;
  assign cgp_core_247 = input_a[30] & cgp_core_244;
  assign cgp_core_248 = cgp_core_245 | cgp_core_247;
  assign cgp_core_250 = input_a[33] ^ input_a[34];
  assign cgp_core_251 = input_a[33] & input_a[34];
  assign cgp_core_252 = input_a[35] ^ input_a[36];
  assign cgp_core_253 = input_a[35] & input_a[36];
  assign cgp_core_254 = cgp_core_250 ^ cgp_core_252;
  assign cgp_core_255 = cgp_core_250 & cgp_core_252;
  assign cgp_core_256 = cgp_core_251 ^ cgp_core_253;
  assign cgp_core_257 = cgp_core_251 & cgp_core_253;
  assign cgp_core_258 = cgp_core_256 | cgp_core_255;
  assign cgp_core_261 = cgp_core_246 ^ cgp_core_254;
  assign cgp_core_262 = cgp_core_246 & cgp_core_254;
  assign cgp_core_263 = cgp_core_248 ^ cgp_core_258;
  assign cgp_core_264 = cgp_core_248 & cgp_core_258;
  assign cgp_core_265 = cgp_core_263 ^ cgp_core_262;
  assign cgp_core_266 = cgp_core_263 & cgp_core_262;
  assign cgp_core_267 = cgp_core_264 | cgp_core_266;
  assign cgp_core_269 = ~(input_a[46] & input_a[43]);
  assign cgp_core_270 = cgp_core_257 | cgp_core_267;
  assign cgp_core_271 = input_a[59] ^ input_a[5];
  assign cgp_core_273 = input_a[37] ^ input_a[38];
  assign cgp_core_274 = input_a[37] & input_a[38];
  assign cgp_core_275 = input_a[39] ^ input_a[40];
  assign cgp_core_276 = input_a[39] & input_a[40];
  assign cgp_core_277 = cgp_core_273 ^ cgp_core_275;
  assign cgp_core_278 = cgp_core_273 & cgp_core_275;
  assign cgp_core_279 = cgp_core_274 ^ cgp_core_276;
  assign cgp_core_280 = cgp_core_274 & cgp_core_276;
  assign cgp_core_281 = cgp_core_279 | cgp_core_278;
  assign cgp_core_282 = ~(input_a[8] ^ input_a[37]);
  assign cgp_core_284 = input_a[41] ^ input_a[42];
  assign cgp_core_285 = input_a[41] & input_a[42];
  assign cgp_core_286 = input_a[43] ^ input_a[44];
  assign cgp_core_287 = input_a[43] & input_a[44];
  assign cgp_core_288 = cgp_core_284 ^ cgp_core_286;
  assign cgp_core_289 = cgp_core_284 & cgp_core_286;
  assign cgp_core_290 = cgp_core_285 ^ cgp_core_287;
  assign cgp_core_291 = cgp_core_285 & cgp_core_287;
  assign cgp_core_292 = cgp_core_290 | cgp_core_289;
  assign cgp_core_293 = ~(input_a[14] | input_a[46]);
  assign cgp_core_295 = cgp_core_277 ^ cgp_core_288;
  assign cgp_core_296 = cgp_core_277 & cgp_core_288;
  assign cgp_core_297 = cgp_core_281 ^ cgp_core_292;
  assign cgp_core_298 = cgp_core_281 & cgp_core_292;
  assign cgp_core_299 = cgp_core_297 ^ cgp_core_296;
  assign cgp_core_300 = cgp_core_297 & cgp_core_296;
  assign cgp_core_301 = cgp_core_298 | cgp_core_300;
  assign cgp_core_302 = cgp_core_280 ^ cgp_core_291;
  assign cgp_core_303 = cgp_core_280 & cgp_core_291;
  assign cgp_core_304 = cgp_core_302 | cgp_core_301;
  assign cgp_core_307 = cgp_core_261 ^ cgp_core_295;
  assign cgp_core_308 = cgp_core_261 & cgp_core_295;
  assign cgp_core_309 = cgp_core_265 ^ cgp_core_299;
  assign cgp_core_310 = cgp_core_265 & cgp_core_299;
  assign cgp_core_311 = cgp_core_309 ^ cgp_core_308;
  assign cgp_core_312 = cgp_core_309 & cgp_core_308;
  assign cgp_core_313 = cgp_core_310 | cgp_core_312;
  assign cgp_core_314 = cgp_core_270 ^ cgp_core_304;
  assign cgp_core_315 = cgp_core_270 & cgp_core_304;
  assign cgp_core_316 = cgp_core_314 ^ cgp_core_313;
  assign cgp_core_317 = cgp_core_314 & cgp_core_313;
  assign cgp_core_318 = cgp_core_315 | cgp_core_317;
  assign cgp_core_320 = ~(input_a[53] & input_a[9]);
  assign cgp_core_321 = cgp_core_303 | cgp_core_318;
  assign cgp_core_323 = ~(input_a[33] | input_a[4]);
  assign cgp_core_324 = input_a[46] ^ input_a[47];
  assign cgp_core_325 = input_a[46] & input_a[47];
  assign cgp_core_326 = input_a[45] ^ cgp_core_324;
  assign cgp_core_327 = input_a[45] & cgp_core_324;
  assign cgp_core_328 = cgp_core_325 | cgp_core_327;
  assign cgp_core_330 = input_a[48] ^ input_a[49];
  assign cgp_core_331 = input_a[48] & input_a[49];
  assign cgp_core_332 = input_a[50] ^ input_a[51];
  assign cgp_core_333 = input_a[50] & input_a[51];
  assign cgp_core_334 = cgp_core_330 ^ cgp_core_332;
  assign cgp_core_335 = cgp_core_330 & cgp_core_332;
  assign cgp_core_336 = cgp_core_331 ^ cgp_core_333;
  assign cgp_core_337 = cgp_core_331 & cgp_core_333;
  assign cgp_core_338 = cgp_core_336 | cgp_core_335;
  assign cgp_core_341 = cgp_core_326 ^ cgp_core_334;
  assign cgp_core_342 = cgp_core_326 & cgp_core_334;
  assign cgp_core_343 = cgp_core_328 ^ cgp_core_338;
  assign cgp_core_344 = cgp_core_328 & cgp_core_338;
  assign cgp_core_345 = cgp_core_343 ^ cgp_core_342;
  assign cgp_core_346 = cgp_core_343 & cgp_core_342;
  assign cgp_core_347 = cgp_core_344 | cgp_core_346;
  assign cgp_core_349 = input_a[18] & input_a[27];
  assign cgp_core_350 = cgp_core_337 | cgp_core_347;
  assign cgp_core_353 = input_a[52] ^ input_a[53];
  assign cgp_core_354 = input_a[52] & input_a[53];
  assign cgp_core_355 = input_a[54] ^ input_a[55];
  assign cgp_core_356 = input_a[54] & input_a[55];
  assign cgp_core_357 = cgp_core_353 ^ cgp_core_355;
  assign cgp_core_358 = cgp_core_353 & cgp_core_355;
  assign cgp_core_359 = cgp_core_354 ^ cgp_core_356;
  assign cgp_core_360 = cgp_core_354 & cgp_core_356;
  assign cgp_core_361 = cgp_core_359 | cgp_core_358;
  assign cgp_core_362 = input_a[22] ^ input_a[59];
  assign cgp_core_364 = input_a[56] ^ input_a[57];
  assign cgp_core_365 = input_a[56] & input_a[57];
  assign cgp_core_366 = input_a[58] ^ input_a[59];
  assign cgp_core_367 = input_a[58] & input_a[59];
  assign cgp_core_368 = cgp_core_364 ^ cgp_core_366;
  assign cgp_core_369 = cgp_core_364 & cgp_core_366;
  assign cgp_core_370 = cgp_core_365 ^ cgp_core_367;
  assign cgp_core_371 = cgp_core_365 & cgp_core_367;
  assign cgp_core_372 = cgp_core_370 | cgp_core_369;
  assign cgp_core_373 = ~input_a[36];
  assign cgp_core_375 = cgp_core_357 ^ cgp_core_368;
  assign cgp_core_376 = cgp_core_357 & cgp_core_368;
  assign cgp_core_377 = cgp_core_361 ^ cgp_core_372;
  assign cgp_core_378 = cgp_core_361 & cgp_core_372;
  assign cgp_core_379 = cgp_core_377 ^ cgp_core_376;
  assign cgp_core_380 = cgp_core_377 & cgp_core_376;
  assign cgp_core_381 = cgp_core_378 | cgp_core_380;
  assign cgp_core_382 = cgp_core_360 ^ cgp_core_371;
  assign cgp_core_383 = cgp_core_360 & cgp_core_371;
  assign cgp_core_384 = cgp_core_382 | cgp_core_381;
  assign cgp_core_385 = input_a[53] & input_a[13];
  assign cgp_core_387 = cgp_core_341 ^ cgp_core_375;
  assign cgp_core_388 = cgp_core_341 & cgp_core_375;
  assign cgp_core_389 = cgp_core_345 ^ cgp_core_379;
  assign cgp_core_390 = cgp_core_345 & cgp_core_379;
  assign cgp_core_391 = cgp_core_389 ^ cgp_core_388;
  assign cgp_core_392 = cgp_core_389 & cgp_core_388;
  assign cgp_core_393 = cgp_core_390 | cgp_core_392;
  assign cgp_core_394 = cgp_core_350 ^ cgp_core_384;
  assign cgp_core_395 = cgp_core_350 & cgp_core_384;
  assign cgp_core_396 = cgp_core_394 ^ cgp_core_393;
  assign cgp_core_397 = cgp_core_394 & cgp_core_393;
  assign cgp_core_398 = cgp_core_395 | cgp_core_397;
  assign cgp_core_400 = ~input_a[0];
  assign cgp_core_401 = cgp_core_383 | cgp_core_398;
  assign cgp_core_403 = ~(input_a[19] ^ input_a[2]);
  assign cgp_core_404 = cgp_core_307 ^ cgp_core_387;
  assign cgp_core_405 = cgp_core_307 & cgp_core_387;
  assign cgp_core_406 = cgp_core_311 ^ cgp_core_391;
  assign cgp_core_407 = cgp_core_311 & cgp_core_391;
  assign cgp_core_408 = cgp_core_406 ^ cgp_core_405;
  assign cgp_core_409 = cgp_core_406 & cgp_core_405;
  assign cgp_core_410 = cgp_core_407 | cgp_core_409;
  assign cgp_core_411 = cgp_core_316 ^ cgp_core_396;
  assign cgp_core_412 = cgp_core_316 & cgp_core_396;
  assign cgp_core_413 = cgp_core_411 ^ cgp_core_410;
  assign cgp_core_414 = cgp_core_411 & cgp_core_410;
  assign cgp_core_415 = cgp_core_412 | cgp_core_414;
  assign cgp_core_416 = cgp_core_321 ^ cgp_core_401;
  assign cgp_core_417 = cgp_core_321 & cgp_core_401;
  assign cgp_core_418 = cgp_core_416 ^ cgp_core_415;
  assign cgp_core_419 = cgp_core_416 & cgp_core_415;
  assign cgp_core_420 = cgp_core_417 | cgp_core_419;
  assign cgp_core_422 = ~(input_a[59] | input_a[48]);
  assign cgp_core_424 = ~(input_a[32] & input_a[14]);
  assign cgp_core_426 = cgp_core_222 ^ cgp_core_404;
  assign cgp_core_427 = cgp_core_222 & cgp_core_404;
  assign cgp_core_428 = cgp_core_226 ^ cgp_core_408;
  assign cgp_core_429 = cgp_core_226 & cgp_core_408;
  assign cgp_core_430 = cgp_core_428 ^ cgp_core_427;
  assign cgp_core_431 = cgp_core_428 & cgp_core_427;
  assign cgp_core_432 = cgp_core_429 | cgp_core_431;
  assign cgp_core_433 = cgp_core_231 ^ cgp_core_413;
  assign cgp_core_434 = cgp_core_231 & cgp_core_413;
  assign cgp_core_435 = cgp_core_433 ^ cgp_core_432;
  assign cgp_core_436 = cgp_core_433 & cgp_core_432;
  assign cgp_core_437 = cgp_core_434 | cgp_core_436;
  assign cgp_core_438 = cgp_core_236 ^ cgp_core_418;
  assign cgp_core_439 = cgp_core_236 & cgp_core_418;
  assign cgp_core_440 = cgp_core_438 ^ cgp_core_437;
  assign cgp_core_441 = cgp_core_438 & cgp_core_437;
  assign cgp_core_442 = cgp_core_439 | cgp_core_441;
  assign cgp_core_443 = cgp_core_238 ^ cgp_core_420;
  assign cgp_core_444 = cgp_core_238 & cgp_core_420;
  assign cgp_core_445 = cgp_core_443 ^ cgp_core_442;
  assign cgp_core_446 = cgp_core_443 & cgp_core_442;
  assign cgp_core_447 = cgp_core_444 | cgp_core_446;
  assign cgp_core_448 = input_a[9] & input_a[50];
  assign cgp_core_449 = ~(input_a[17] | input_a[15]);
  assign cgp_core_450 = ~(input_a[22] ^ input_a[13]);
  assign cgp_core_452 = input_a[55] & input_a[28];

  assign cgp_out[0] = cgp_core_426;
  assign cgp_out[1] = cgp_core_430;
  assign cgp_out[2] = cgp_core_435;
  assign cgp_out[3] = cgp_core_440;
  assign cgp_out[4] = cgp_core_445;
  assign cgp_out[5] = cgp_core_447;
endmodule

module cmp_neg(input [28:0] input_a, output [4:0] cgp_out);
  wire cgp_core_031;
  wire cgp_core_032;
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_035;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_102;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_112;
  wire cgp_core_113;
  wire cgp_core_114;
  wire cgp_core_115;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_118;
  wire cgp_core_119;
  wire cgp_core_120;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_129;
  wire cgp_core_131;
  wire cgp_core_132;
  wire cgp_core_135;
  wire cgp_core_136;
  wire cgp_core_137;
  wire cgp_core_138;
  wire cgp_core_139;
  wire cgp_core_140;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_146;
  wire cgp_core_147;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_150;
  wire cgp_core_151;
  wire cgp_core_152;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_157;
  wire cgp_core_158;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_161;
  wire cgp_core_162;
  wire cgp_core_163;
  wire cgp_core_164;
  wire cgp_core_165;
  wire cgp_core_166;
  wire cgp_core_167;
  wire cgp_core_169;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_180;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_188;
  wire cgp_core_189;
  wire cgp_core_190;
  wire cgp_core_191;
  wire cgp_core_192;
  wire cgp_core_193;
  wire cgp_core_194;
  wire cgp_core_195;
  wire cgp_core_196;
  wire cgp_core_197;
  wire cgp_core_198;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_203;
  wire cgp_core_205;
  wire cgp_core_206;
  wire cgp_core_207;

  assign cgp_core_031 = input_a[1] ^ input_a[2];
  assign cgp_core_032 = input_a[1] & input_a[2];
  assign cgp_core_033 = input_a[0] ^ cgp_core_031;
  assign cgp_core_034 = input_a[0] & cgp_core_031;
  assign cgp_core_035 = cgp_core_032 | cgp_core_034;
  assign cgp_core_037 = input_a[3] ^ input_a[4];
  assign cgp_core_038 = input_a[3] & input_a[4];
  assign cgp_core_039 = input_a[5] ^ input_a[6];
  assign cgp_core_040 = input_a[5] & input_a[6];
  assign cgp_core_041 = cgp_core_037 ^ cgp_core_039;
  assign cgp_core_042 = cgp_core_037 & cgp_core_039;
  assign cgp_core_043 = cgp_core_038 ^ cgp_core_040;
  assign cgp_core_044 = cgp_core_038 & cgp_core_040;
  assign cgp_core_045 = cgp_core_043 | cgp_core_042;
  assign cgp_core_046 = input_a[5] ^ input_a[7];
  assign cgp_core_048 = cgp_core_033 ^ cgp_core_041;
  assign cgp_core_049 = cgp_core_033 & cgp_core_041;
  assign cgp_core_050 = cgp_core_035 ^ cgp_core_045;
  assign cgp_core_051 = cgp_core_035 & cgp_core_045;
  assign cgp_core_052 = cgp_core_050 ^ cgp_core_049;
  assign cgp_core_053 = cgp_core_050 & cgp_core_049;
  assign cgp_core_054 = cgp_core_051 | cgp_core_053;
  assign cgp_core_057 = cgp_core_044 | cgp_core_054;
  assign cgp_core_058 = ~input_a[19];
  assign cgp_core_060 = input_a[8] ^ input_a[9];
  assign cgp_core_061 = input_a[8] & input_a[9];
  assign cgp_core_062 = input_a[7] ^ cgp_core_060;
  assign cgp_core_063 = input_a[7] & cgp_core_060;
  assign cgp_core_064 = cgp_core_061 | cgp_core_063;
  assign cgp_core_066 = input_a[10] ^ input_a[11];
  assign cgp_core_067 = input_a[10] & input_a[11];
  assign cgp_core_068 = input_a[12] ^ input_a[13];
  assign cgp_core_069 = input_a[12] & input_a[13];
  assign cgp_core_070 = cgp_core_066 ^ cgp_core_068;
  assign cgp_core_071 = cgp_core_066 & cgp_core_068;
  assign cgp_core_072 = cgp_core_067 ^ cgp_core_069;
  assign cgp_core_073 = cgp_core_067 & cgp_core_069;
  assign cgp_core_074 = cgp_core_072 | cgp_core_071;
  assign cgp_core_075 = input_a[19] ^ input_a[10];
  assign cgp_core_077 = cgp_core_062 ^ cgp_core_070;
  assign cgp_core_078 = cgp_core_062 & cgp_core_070;
  assign cgp_core_079 = cgp_core_064 ^ cgp_core_074;
  assign cgp_core_080 = cgp_core_064 & cgp_core_074;
  assign cgp_core_081 = cgp_core_079 ^ cgp_core_078;
  assign cgp_core_082 = cgp_core_079 & cgp_core_078;
  assign cgp_core_083 = cgp_core_080 | cgp_core_082;
  assign cgp_core_085 = ~(input_a[27] & input_a[20]);
  assign cgp_core_086 = cgp_core_073 | cgp_core_083;
  assign cgp_core_087 = ~(input_a[13] ^ input_a[0]);
  assign cgp_core_088 = input_a[21] ^ input_a[18];
  assign cgp_core_089 = cgp_core_048 ^ cgp_core_077;
  assign cgp_core_090 = cgp_core_048 & cgp_core_077;
  assign cgp_core_091 = cgp_core_052 ^ cgp_core_081;
  assign cgp_core_092 = cgp_core_052 & cgp_core_081;
  assign cgp_core_093 = cgp_core_091 ^ cgp_core_090;
  assign cgp_core_094 = cgp_core_091 & cgp_core_090;
  assign cgp_core_095 = cgp_core_092 | cgp_core_094;
  assign cgp_core_096 = cgp_core_057 ^ cgp_core_086;
  assign cgp_core_097 = cgp_core_057 & cgp_core_086;
  assign cgp_core_098 = cgp_core_096 ^ cgp_core_095;
  assign cgp_core_099 = cgp_core_096 & cgp_core_095;
  assign cgp_core_100 = cgp_core_097 | cgp_core_099;
  assign cgp_core_102 = input_a[19] ^ input_a[7];
  assign cgp_core_106 = input_a[15] ^ input_a[16];
  assign cgp_core_107 = input_a[15] & input_a[16];
  assign cgp_core_108 = input_a[14] ^ cgp_core_106;
  assign cgp_core_109 = input_a[14] & cgp_core_106;
  assign cgp_core_110 = cgp_core_107 | cgp_core_109;
  assign cgp_core_112 = input_a[17] ^ input_a[18];
  assign cgp_core_113 = input_a[17] & input_a[18];
  assign cgp_core_114 = input_a[19] ^ input_a[20];
  assign cgp_core_115 = input_a[19] & input_a[20];
  assign cgp_core_116 = cgp_core_112 ^ cgp_core_114;
  assign cgp_core_117 = cgp_core_112 & cgp_core_114;
  assign cgp_core_118 = cgp_core_113 ^ cgp_core_115;
  assign cgp_core_119 = cgp_core_113 & cgp_core_115;
  assign cgp_core_120 = cgp_core_118 | cgp_core_117;
  assign cgp_core_123 = cgp_core_108 ^ cgp_core_116;
  assign cgp_core_124 = cgp_core_108 & cgp_core_116;
  assign cgp_core_125 = cgp_core_110 ^ cgp_core_120;
  assign cgp_core_126 = cgp_core_110 & cgp_core_120;
  assign cgp_core_127 = cgp_core_125 ^ cgp_core_124;
  assign cgp_core_128 = cgp_core_125 & cgp_core_124;
  assign cgp_core_129 = cgp_core_126 | cgp_core_128;
  assign cgp_core_131 = ~input_a[19];
  assign cgp_core_132 = cgp_core_119 | cgp_core_129;
  assign cgp_core_135 = input_a[21] ^ input_a[22];
  assign cgp_core_136 = input_a[21] & input_a[22];
  assign cgp_core_137 = input_a[23] ^ input_a[24];
  assign cgp_core_138 = input_a[23] & input_a[24];
  assign cgp_core_139 = cgp_core_135 ^ cgp_core_137;
  assign cgp_core_140 = cgp_core_135 & cgp_core_137;
  assign cgp_core_141 = cgp_core_136 ^ cgp_core_138;
  assign cgp_core_142 = cgp_core_136 & cgp_core_138;
  assign cgp_core_143 = cgp_core_141 | cgp_core_140;
  assign cgp_core_144 = ~(input_a[26] | input_a[27]);
  assign cgp_core_146 = input_a[25] ^ input_a[26];
  assign cgp_core_147 = input_a[25] & input_a[26];
  assign cgp_core_148 = input_a[27] ^ input_a[28];
  assign cgp_core_149 = input_a[27] & input_a[28];
  assign cgp_core_150 = cgp_core_146 ^ cgp_core_148;
  assign cgp_core_151 = cgp_core_146 & cgp_core_148;
  assign cgp_core_152 = cgp_core_147 ^ cgp_core_149;
  assign cgp_core_153 = cgp_core_147 & cgp_core_149;
  assign cgp_core_154 = cgp_core_152 | cgp_core_151;
  assign cgp_core_157 = cgp_core_139 ^ cgp_core_150;
  assign cgp_core_158 = cgp_core_139 & cgp_core_150;
  assign cgp_core_159 = cgp_core_143 ^ cgp_core_154;
  assign cgp_core_160 = cgp_core_143 & cgp_core_154;
  assign cgp_core_161 = cgp_core_159 ^ cgp_core_158;
  assign cgp_core_162 = cgp_core_159 & cgp_core_158;
  assign cgp_core_163 = cgp_core_160 | cgp_core_162;
  assign cgp_core_164 = cgp_core_142 ^ cgp_core_153;
  assign cgp_core_165 = cgp_core_142 & cgp_core_153;
  assign cgp_core_166 = cgp_core_164 | cgp_core_163;
  assign cgp_core_167 = input_a[16] ^ input_a[8];
  assign cgp_core_169 = cgp_core_123 ^ cgp_core_157;
  assign cgp_core_170 = cgp_core_123 & cgp_core_157;
  assign cgp_core_171 = cgp_core_127 ^ cgp_core_161;
  assign cgp_core_172 = cgp_core_127 & cgp_core_161;
  assign cgp_core_173 = cgp_core_171 ^ cgp_core_170;
  assign cgp_core_174 = cgp_core_171 & cgp_core_170;
  assign cgp_core_175 = cgp_core_172 | cgp_core_174;
  assign cgp_core_176 = cgp_core_132 ^ cgp_core_166;
  assign cgp_core_177 = cgp_core_132 & cgp_core_166;
  assign cgp_core_178 = cgp_core_176 ^ cgp_core_175;
  assign cgp_core_179 = cgp_core_176 & cgp_core_175;
  assign cgp_core_180 = cgp_core_177 | cgp_core_179;
  assign cgp_core_182 = ~(input_a[4] & input_a[25]);
  assign cgp_core_183 = cgp_core_165 | cgp_core_180;
  assign cgp_core_184 = ~(input_a[11] ^ input_a[26]);
  assign cgp_core_185 = input_a[2] ^ input_a[2];
  assign cgp_core_186 = cgp_core_089 ^ cgp_core_169;
  assign cgp_core_187 = cgp_core_089 & cgp_core_169;
  assign cgp_core_188 = cgp_core_093 ^ cgp_core_173;
  assign cgp_core_189 = cgp_core_093 & cgp_core_173;
  assign cgp_core_190 = cgp_core_188 ^ cgp_core_187;
  assign cgp_core_191 = cgp_core_188 & cgp_core_187;
  assign cgp_core_192 = cgp_core_189 | cgp_core_191;
  assign cgp_core_193 = cgp_core_098 ^ cgp_core_178;
  assign cgp_core_194 = cgp_core_098 & cgp_core_178;
  assign cgp_core_195 = cgp_core_193 ^ cgp_core_192;
  assign cgp_core_196 = cgp_core_193 & cgp_core_192;
  assign cgp_core_197 = cgp_core_194 | cgp_core_196;
  assign cgp_core_198 = cgp_core_100 ^ cgp_core_183;
  assign cgp_core_199 = cgp_core_100 & cgp_core_183;
  assign cgp_core_200 = cgp_core_198 ^ cgp_core_197;
  assign cgp_core_201 = cgp_core_198 & cgp_core_197;
  assign cgp_core_202 = cgp_core_199 | cgp_core_201;
  assign cgp_core_203 = ~(input_a[27] ^ input_a[17]);
  assign cgp_core_205 = ~input_a[10];
  assign cgp_core_206 = input_a[6] & input_a[22];
  assign cgp_core_207 = input_a[14] | input_a[10];

  assign cgp_out[0] = cgp_core_186;
  assign cgp_out[1] = cgp_core_190;
  assign cgp_out[2] = cgp_core_195;
  assign cgp_out[3] = cgp_core_200;
  assign cgp_out[4] = cgp_core_202;
endmodule
module pcc(input [59:0] pos, input [28:0] neg, output outval);
    wire [5:0] cnt_pos;
    wire [4:0] cnt_neg;

    cmp_pos ipos(pos, cnt_pos);
    cmp_neg ineg(neg, cnt_neg);

    assign outval = (cnt_pos >= cnt_neg);
endmodule
