// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.88865
// WCE=18.0
// EP=0.834026%
// Printed PDK parameters:
//  Area=62411156.0
//  Delay=69684504.0
//  Power=3092900.0

module popcount38_u38d(input [37:0] input_a, output [5:0] popcount38_u38d_out);
  wire popcount38_u38d_core_040;
  wire popcount38_u38d_core_042;
  wire popcount38_u38d_core_043;
  wire popcount38_u38d_core_047;
  wire popcount38_u38d_core_049;
  wire popcount38_u38d_core_051;
  wire popcount38_u38d_core_054;
  wire popcount38_u38d_core_057;
  wire popcount38_u38d_core_059;
  wire popcount38_u38d_core_060;
  wire popcount38_u38d_core_061;
  wire popcount38_u38d_core_063;
  wire popcount38_u38d_core_064;
  wire popcount38_u38d_core_067;
  wire popcount38_u38d_core_068;
  wire popcount38_u38d_core_070_not;
  wire popcount38_u38d_core_073;
  wire popcount38_u38d_core_077;
  wire popcount38_u38d_core_078;
  wire popcount38_u38d_core_082;
  wire popcount38_u38d_core_083;
  wire popcount38_u38d_core_084;
  wire popcount38_u38d_core_085;
  wire popcount38_u38d_core_090;
  wire popcount38_u38d_core_092;
  wire popcount38_u38d_core_093;
  wire popcount38_u38d_core_094;
  wire popcount38_u38d_core_095;
  wire popcount38_u38d_core_096;
  wire popcount38_u38d_core_100;
  wire popcount38_u38d_core_101;
  wire popcount38_u38d_core_102;
  wire popcount38_u38d_core_103;
  wire popcount38_u38d_core_104;
  wire popcount38_u38d_core_105;
  wire popcount38_u38d_core_107_not;
  wire popcount38_u38d_core_109;
  wire popcount38_u38d_core_110;
  wire popcount38_u38d_core_111;
  wire popcount38_u38d_core_112;
  wire popcount38_u38d_core_113;
  wire popcount38_u38d_core_115;
  wire popcount38_u38d_core_117;
  wire popcount38_u38d_core_118;
  wire popcount38_u38d_core_119;
  wire popcount38_u38d_core_120;
  wire popcount38_u38d_core_121;
  wire popcount38_u38d_core_122;
  wire popcount38_u38d_core_123;
  wire popcount38_u38d_core_124;
  wire popcount38_u38d_core_125;
  wire popcount38_u38d_core_126;
  wire popcount38_u38d_core_127;
  wire popcount38_u38d_core_129;
  wire popcount38_u38d_core_131;
  wire popcount38_u38d_core_132;
  wire popcount38_u38d_core_133;
  wire popcount38_u38d_core_135;
  wire popcount38_u38d_core_136;
  wire popcount38_u38d_core_140;
  wire popcount38_u38d_core_141;
  wire popcount38_u38d_core_142;
  wire popcount38_u38d_core_143;
  wire popcount38_u38d_core_144;
  wire popcount38_u38d_core_146;
  wire popcount38_u38d_core_147;
  wire popcount38_u38d_core_148;
  wire popcount38_u38d_core_149;
  wire popcount38_u38d_core_151;
  wire popcount38_u38d_core_153;
  wire popcount38_u38d_core_154;
  wire popcount38_u38d_core_155;
  wire popcount38_u38d_core_156;
  wire popcount38_u38d_core_157;
  wire popcount38_u38d_core_158;
  wire popcount38_u38d_core_159;
  wire popcount38_u38d_core_160;
  wire popcount38_u38d_core_161;
  wire popcount38_u38d_core_162;
  wire popcount38_u38d_core_163;
  wire popcount38_u38d_core_164;
  wire popcount38_u38d_core_167;
  wire popcount38_u38d_core_168;
  wire popcount38_u38d_core_169;
  wire popcount38_u38d_core_171;
  wire popcount38_u38d_core_172;
  wire popcount38_u38d_core_174;
  wire popcount38_u38d_core_176;
  wire popcount38_u38d_core_177;
  wire popcount38_u38d_core_180;
  wire popcount38_u38d_core_182;
  wire popcount38_u38d_core_183;
  wire popcount38_u38d_core_184_not;
  wire popcount38_u38d_core_185;
  wire popcount38_u38d_core_186;
  wire popcount38_u38d_core_188;
  wire popcount38_u38d_core_191;
  wire popcount38_u38d_core_192;
  wire popcount38_u38d_core_193;
  wire popcount38_u38d_core_194;
  wire popcount38_u38d_core_196;
  wire popcount38_u38d_core_197;
  wire popcount38_u38d_core_198;
  wire popcount38_u38d_core_200;
  wire popcount38_u38d_core_201_not;
  wire popcount38_u38d_core_203;
  wire popcount38_u38d_core_204;
  wire popcount38_u38d_core_205_not;
  wire popcount38_u38d_core_206;
  wire popcount38_u38d_core_207;
  wire popcount38_u38d_core_208;
  wire popcount38_u38d_core_209;
  wire popcount38_u38d_core_212;
  wire popcount38_u38d_core_213;
  wire popcount38_u38d_core_215;
  wire popcount38_u38d_core_216;
  wire popcount38_u38d_core_217;
  wire popcount38_u38d_core_219;
  wire popcount38_u38d_core_220;
  wire popcount38_u38d_core_221;
  wire popcount38_u38d_core_222;
  wire popcount38_u38d_core_223;
  wire popcount38_u38d_core_224;
  wire popcount38_u38d_core_225;
  wire popcount38_u38d_core_226;
  wire popcount38_u38d_core_227;
  wire popcount38_u38d_core_228;
  wire popcount38_u38d_core_229;
  wire popcount38_u38d_core_231;
  wire popcount38_u38d_core_232;
  wire popcount38_u38d_core_233;
  wire popcount38_u38d_core_234;
  wire popcount38_u38d_core_236;
  wire popcount38_u38d_core_238;
  wire popcount38_u38d_core_239;
  wire popcount38_u38d_core_240;
  wire popcount38_u38d_core_241;
  wire popcount38_u38d_core_242;
  wire popcount38_u38d_core_244;
  wire popcount38_u38d_core_246;
  wire popcount38_u38d_core_250;
  wire popcount38_u38d_core_251;
  wire popcount38_u38d_core_252;
  wire popcount38_u38d_core_255;
  wire popcount38_u38d_core_256;
  wire popcount38_u38d_core_257;
  wire popcount38_u38d_core_258;
  wire popcount38_u38d_core_259;
  wire popcount38_u38d_core_261;
  wire popcount38_u38d_core_262;
  wire popcount38_u38d_core_263;
  wire popcount38_u38d_core_265;
  wire popcount38_u38d_core_266;
  wire popcount38_u38d_core_268;
  wire popcount38_u38d_core_270_not;
  wire popcount38_u38d_core_272;
  wire popcount38_u38d_core_273;
  wire popcount38_u38d_core_274;
  wire popcount38_u38d_core_275;
  wire popcount38_u38d_core_276;
  wire popcount38_u38d_core_277;
  wire popcount38_u38d_core_278;
  wire popcount38_u38d_core_279;
  wire popcount38_u38d_core_280;
  wire popcount38_u38d_core_281;
  wire popcount38_u38d_core_282;
  wire popcount38_u38d_core_283;
  wire popcount38_u38d_core_284;
  wire popcount38_u38d_core_285;
  wire popcount38_u38d_core_286;
  wire popcount38_u38d_core_288;
  wire popcount38_u38d_core_290;
  wire popcount38_u38d_core_291;
  wire popcount38_u38d_core_292;
  wire popcount38_u38d_core_293_not;
  wire popcount38_u38d_core_295;

  assign popcount38_u38d_core_040 = ~input_a[5];
  assign popcount38_u38d_core_042 = input_a[30] | input_a[37];
  assign popcount38_u38d_core_043 = input_a[3] ^ input_a[34];
  assign popcount38_u38d_core_047 = input_a[15] | input_a[17];
  assign popcount38_u38d_core_049 = ~(input_a[14] ^ input_a[2]);
  assign popcount38_u38d_core_051 = input_a[28] ^ input_a[25];
  assign popcount38_u38d_core_054 = input_a[6] & input_a[4];
  assign popcount38_u38d_core_057 = popcount38_u38d_core_054 | input_a[32];
  assign popcount38_u38d_core_059 = input_a[23] ^ input_a[25];
  assign popcount38_u38d_core_060 = input_a[8] & input_a[25];
  assign popcount38_u38d_core_061 = input_a[32] | popcount38_u38d_core_057;
  assign popcount38_u38d_core_063 = popcount38_u38d_core_061 ^ popcount38_u38d_core_060;
  assign popcount38_u38d_core_064 = input_a[24] & popcount38_u38d_core_060;
  assign popcount38_u38d_core_067 = ~(input_a[27] ^ input_a[25]);
  assign popcount38_u38d_core_068 = ~input_a[32];
  assign popcount38_u38d_core_070_not = ~popcount38_u38d_core_063;
  assign popcount38_u38d_core_073 = input_a[15] | input_a[2];
  assign popcount38_u38d_core_077 = popcount38_u38d_core_064 | popcount38_u38d_core_063;
  assign popcount38_u38d_core_078 = ~(input_a[4] & input_a[18]);
  assign popcount38_u38d_core_082 = input_a[9] ^ input_a[10];
  assign popcount38_u38d_core_083 = input_a[9] & input_a[10];
  assign popcount38_u38d_core_084 = input_a[7] | input_a[24];
  assign popcount38_u38d_core_085 = input_a[34] | input_a[10];
  assign popcount38_u38d_core_090 = ~(input_a[8] & input_a[37]);
  assign popcount38_u38d_core_092 = popcount38_u38d_core_083 ^ input_a[37];
  assign popcount38_u38d_core_093 = input_a[10] & input_a[37];
  assign popcount38_u38d_core_094 = popcount38_u38d_core_092 ^ popcount38_u38d_core_082;
  assign popcount38_u38d_core_095 = popcount38_u38d_core_092 & popcount38_u38d_core_082;
  assign popcount38_u38d_core_096 = popcount38_u38d_core_093 | popcount38_u38d_core_095;
  assign popcount38_u38d_core_100 = input_a[23] & input_a[15];
  assign popcount38_u38d_core_101 = input_a[17] ^ input_a[18];
  assign popcount38_u38d_core_102 = input_a[17] & input_a[18];
  assign popcount38_u38d_core_103 = ~(input_a[16] & popcount38_u38d_core_101);
  assign popcount38_u38d_core_104 = input_a[16] & popcount38_u38d_core_101;
  assign popcount38_u38d_core_105 = popcount38_u38d_core_102 | popcount38_u38d_core_104;
  assign popcount38_u38d_core_107_not = ~popcount38_u38d_core_103;
  assign popcount38_u38d_core_109 = popcount38_u38d_core_100 ^ popcount38_u38d_core_105;
  assign popcount38_u38d_core_110 = popcount38_u38d_core_100 & popcount38_u38d_core_105;
  assign popcount38_u38d_core_111 = popcount38_u38d_core_109 ^ popcount38_u38d_core_103;
  assign popcount38_u38d_core_112 = popcount38_u38d_core_109 & popcount38_u38d_core_103;
  assign popcount38_u38d_core_113 = popcount38_u38d_core_110 | popcount38_u38d_core_112;
  assign popcount38_u38d_core_115 = ~(input_a[0] & input_a[11]);
  assign popcount38_u38d_core_117 = popcount38_u38d_core_090 & popcount38_u38d_core_107_not;
  assign popcount38_u38d_core_118 = popcount38_u38d_core_094 ^ popcount38_u38d_core_111;
  assign popcount38_u38d_core_119 = popcount38_u38d_core_094 & popcount38_u38d_core_111;
  assign popcount38_u38d_core_120 = popcount38_u38d_core_118 ^ popcount38_u38d_core_117;
  assign popcount38_u38d_core_121 = popcount38_u38d_core_118 & popcount38_u38d_core_117;
  assign popcount38_u38d_core_122 = popcount38_u38d_core_119 | popcount38_u38d_core_121;
  assign popcount38_u38d_core_123 = popcount38_u38d_core_096 ^ popcount38_u38d_core_113;
  assign popcount38_u38d_core_124 = popcount38_u38d_core_096 & popcount38_u38d_core_113;
  assign popcount38_u38d_core_125 = popcount38_u38d_core_123 ^ popcount38_u38d_core_122;
  assign popcount38_u38d_core_126 = popcount38_u38d_core_123 & popcount38_u38d_core_122;
  assign popcount38_u38d_core_127 = popcount38_u38d_core_124 | popcount38_u38d_core_126;
  assign popcount38_u38d_core_129 = input_a[10] ^ input_a[10];
  assign popcount38_u38d_core_131 = input_a[22] | input_a[32];
  assign popcount38_u38d_core_132 = ~input_a[20];
  assign popcount38_u38d_core_133 = input_a[0] & input_a[28];
  assign popcount38_u38d_core_135 = popcount38_u38d_core_070_not ^ popcount38_u38d_core_120;
  assign popcount38_u38d_core_136 = popcount38_u38d_core_070_not & popcount38_u38d_core_120;
  assign popcount38_u38d_core_140 = popcount38_u38d_core_077 ^ popcount38_u38d_core_125;
  assign popcount38_u38d_core_141 = popcount38_u38d_core_077 & popcount38_u38d_core_125;
  assign popcount38_u38d_core_142 = popcount38_u38d_core_140 ^ popcount38_u38d_core_136;
  assign popcount38_u38d_core_143 = popcount38_u38d_core_140 & popcount38_u38d_core_136;
  assign popcount38_u38d_core_144 = popcount38_u38d_core_141 | popcount38_u38d_core_143;
  assign popcount38_u38d_core_146 = ~(input_a[33] ^ input_a[3]);
  assign popcount38_u38d_core_147 = popcount38_u38d_core_127 | popcount38_u38d_core_144;
  assign popcount38_u38d_core_148 = input_a[14] & input_a[4];
  assign popcount38_u38d_core_149 = ~(input_a[16] | input_a[11]);
  assign popcount38_u38d_core_151 = ~(input_a[22] & input_a[20]);
  assign popcount38_u38d_core_153 = ~(input_a[29] & input_a[0]);
  assign popcount38_u38d_core_154 = input_a[35] | input_a[4];
  assign popcount38_u38d_core_155 = input_a[6] ^ input_a[12];
  assign popcount38_u38d_core_156 = input_a[0] & input_a[36];
  assign popcount38_u38d_core_157 = input_a[21] ^ input_a[22];
  assign popcount38_u38d_core_158 = input_a[21] & input_a[22];
  assign popcount38_u38d_core_159 = input_a[30] ^ input_a[6];
  assign popcount38_u38d_core_160 = input_a[19] & popcount38_u38d_core_157;
  assign popcount38_u38d_core_161 = popcount38_u38d_core_156 ^ popcount38_u38d_core_158;
  assign popcount38_u38d_core_162 = popcount38_u38d_core_156 & popcount38_u38d_core_158;
  assign popcount38_u38d_core_163 = popcount38_u38d_core_161 | popcount38_u38d_core_160;
  assign popcount38_u38d_core_164 = ~(input_a[22] & input_a[34]);
  assign popcount38_u38d_core_167 = ~input_a[34];
  assign popcount38_u38d_core_168 = input_a[26] ^ input_a[27];
  assign popcount38_u38d_core_169 = input_a[26] & input_a[27];
  assign popcount38_u38d_core_171 = input_a[25] & popcount38_u38d_core_168;
  assign popcount38_u38d_core_172 = popcount38_u38d_core_169 | popcount38_u38d_core_171;
  assign popcount38_u38d_core_174 = input_a[4] | input_a[33];
  assign popcount38_u38d_core_176 = input_a[8] | popcount38_u38d_core_172;
  assign popcount38_u38d_core_177 = input_a[12] | popcount38_u38d_core_172;
  assign popcount38_u38d_core_180 = input_a[1] | input_a[27];
  assign popcount38_u38d_core_182 = ~input_a[13];
  assign popcount38_u38d_core_183 = input_a[24] ^ input_a[13];
  assign popcount38_u38d_core_184_not = ~input_a[36];
  assign popcount38_u38d_core_185 = popcount38_u38d_core_163 ^ popcount38_u38d_core_176;
  assign popcount38_u38d_core_186 = popcount38_u38d_core_163 & popcount38_u38d_core_176;
  assign popcount38_u38d_core_188 = input_a[35] & input_a[32];
  assign popcount38_u38d_core_191 = ~(input_a[20] ^ input_a[4]);
  assign popcount38_u38d_core_192 = popcount38_u38d_core_162 | popcount38_u38d_core_186;
  assign popcount38_u38d_core_193 = ~(input_a[33] | input_a[0]);
  assign popcount38_u38d_core_194 = ~input_a[1];
  assign popcount38_u38d_core_196 = ~(input_a[23] & input_a[22]);
  assign popcount38_u38d_core_197 = input_a[28] ^ input_a[29];
  assign popcount38_u38d_core_198 = input_a[28] & input_a[29];
  assign popcount38_u38d_core_200 = input_a[3] & input_a[12];
  assign popcount38_u38d_core_201_not = ~input_a[30];
  assign popcount38_u38d_core_203 = popcount38_u38d_core_200 ^ input_a[30];
  assign popcount38_u38d_core_204 = popcount38_u38d_core_200 & input_a[30];
  assign popcount38_u38d_core_205_not = ~input_a[32];
  assign popcount38_u38d_core_206 = popcount38_u38d_core_197 & popcount38_u38d_core_201_not;
  assign popcount38_u38d_core_207 = popcount38_u38d_core_198 ^ popcount38_u38d_core_203;
  assign popcount38_u38d_core_208 = popcount38_u38d_core_198 & popcount38_u38d_core_203;
  assign popcount38_u38d_core_209 = popcount38_u38d_core_207 | popcount38_u38d_core_206;
  assign popcount38_u38d_core_212 = popcount38_u38d_core_204 | popcount38_u38d_core_208;
  assign popcount38_u38d_core_213 = ~(input_a[37] ^ input_a[34]);
  assign popcount38_u38d_core_215 = input_a[33] & input_a[20];
  assign popcount38_u38d_core_216 = ~(input_a[35] & input_a[37]);
  assign popcount38_u38d_core_217 = input_a[4] ^ input_a[12];
  assign popcount38_u38d_core_219 = input_a[35] & popcount38_u38d_core_216;
  assign popcount38_u38d_core_220 = input_a[13] | popcount38_u38d_core_219;
  assign popcount38_u38d_core_221 = input_a[37] & popcount38_u38d_core_219;
  assign popcount38_u38d_core_222 = input_a[36] | input_a[31];
  assign popcount38_u38d_core_223 = input_a[11] & input_a[31];
  assign popcount38_u38d_core_224 = popcount38_u38d_core_215 ^ popcount38_u38d_core_220;
  assign popcount38_u38d_core_225 = popcount38_u38d_core_215 & popcount38_u38d_core_220;
  assign popcount38_u38d_core_226 = popcount38_u38d_core_224 ^ popcount38_u38d_core_223;
  assign popcount38_u38d_core_227 = popcount38_u38d_core_224 & popcount38_u38d_core_223;
  assign popcount38_u38d_core_228 = popcount38_u38d_core_225 | popcount38_u38d_core_227;
  assign popcount38_u38d_core_229 = popcount38_u38d_core_221 | popcount38_u38d_core_228;
  assign popcount38_u38d_core_231 = ~input_a[27];
  assign popcount38_u38d_core_232 = ~(input_a[25] | input_a[0]);
  assign popcount38_u38d_core_233 = popcount38_u38d_core_209 ^ popcount38_u38d_core_226;
  assign popcount38_u38d_core_234 = popcount38_u38d_core_209 & popcount38_u38d_core_226;
  assign popcount38_u38d_core_236 = ~(input_a[20] | input_a[37]);
  assign popcount38_u38d_core_238 = popcount38_u38d_core_212 ^ popcount38_u38d_core_229;
  assign popcount38_u38d_core_239 = popcount38_u38d_core_212 & popcount38_u38d_core_229;
  assign popcount38_u38d_core_240 = popcount38_u38d_core_238 ^ popcount38_u38d_core_234;
  assign popcount38_u38d_core_241 = popcount38_u38d_core_238 & popcount38_u38d_core_234;
  assign popcount38_u38d_core_242 = popcount38_u38d_core_239 | popcount38_u38d_core_241;
  assign popcount38_u38d_core_244 = input_a[33] | input_a[32];
  assign popcount38_u38d_core_246 = input_a[6] & input_a[3];
  assign popcount38_u38d_core_250 = popcount38_u38d_core_185 ^ popcount38_u38d_core_233;
  assign popcount38_u38d_core_251 = popcount38_u38d_core_185 & popcount38_u38d_core_233;
  assign popcount38_u38d_core_252 = popcount38_u38d_core_250 | input_a[5];
  assign popcount38_u38d_core_255 = popcount38_u38d_core_192 ^ popcount38_u38d_core_240;
  assign popcount38_u38d_core_256 = popcount38_u38d_core_192 & popcount38_u38d_core_240;
  assign popcount38_u38d_core_257 = popcount38_u38d_core_255 ^ popcount38_u38d_core_251;
  assign popcount38_u38d_core_258 = popcount38_u38d_core_255 & popcount38_u38d_core_251;
  assign popcount38_u38d_core_259 = popcount38_u38d_core_256 | popcount38_u38d_core_258;
  assign popcount38_u38d_core_261 = input_a[15] & input_a[32];
  assign popcount38_u38d_core_262 = popcount38_u38d_core_242 | popcount38_u38d_core_259;
  assign popcount38_u38d_core_263 = input_a[23] | input_a[17];
  assign popcount38_u38d_core_265 = input_a[22] & input_a[4];
  assign popcount38_u38d_core_266 = ~(input_a[8] & input_a[3]);
  assign popcount38_u38d_core_268 = input_a[28] & input_a[11];
  assign popcount38_u38d_core_270_not = ~input_a[1];
  assign popcount38_u38d_core_272 = popcount38_u38d_core_135 ^ popcount38_u38d_core_252;
  assign popcount38_u38d_core_273 = popcount38_u38d_core_135 & popcount38_u38d_core_252;
  assign popcount38_u38d_core_274 = popcount38_u38d_core_272 ^ input_a[1];
  assign popcount38_u38d_core_275 = popcount38_u38d_core_272 & input_a[1];
  assign popcount38_u38d_core_276 = popcount38_u38d_core_273 | popcount38_u38d_core_275;
  assign popcount38_u38d_core_277 = popcount38_u38d_core_142 ^ popcount38_u38d_core_257;
  assign popcount38_u38d_core_278 = popcount38_u38d_core_142 & popcount38_u38d_core_257;
  assign popcount38_u38d_core_279 = popcount38_u38d_core_277 ^ popcount38_u38d_core_276;
  assign popcount38_u38d_core_280 = popcount38_u38d_core_277 & popcount38_u38d_core_276;
  assign popcount38_u38d_core_281 = popcount38_u38d_core_278 | popcount38_u38d_core_280;
  assign popcount38_u38d_core_282 = popcount38_u38d_core_147 ^ popcount38_u38d_core_262;
  assign popcount38_u38d_core_283 = popcount38_u38d_core_147 & popcount38_u38d_core_262;
  assign popcount38_u38d_core_284 = popcount38_u38d_core_282 ^ popcount38_u38d_core_281;
  assign popcount38_u38d_core_285 = popcount38_u38d_core_282 & popcount38_u38d_core_281;
  assign popcount38_u38d_core_286 = popcount38_u38d_core_283 | popcount38_u38d_core_285;
  assign popcount38_u38d_core_288 = ~(input_a[17] ^ input_a[32]);
  assign popcount38_u38d_core_290 = input_a[13] & input_a[1];
  assign popcount38_u38d_core_291 = ~(input_a[13] | input_a[4]);
  assign popcount38_u38d_core_292 = ~(input_a[27] | input_a[24]);
  assign popcount38_u38d_core_293_not = ~input_a[19];
  assign popcount38_u38d_core_295 = input_a[34] & input_a[15];

  assign popcount38_u38d_out[0] = popcount38_u38d_core_270_not;
  assign popcount38_u38d_out[1] = popcount38_u38d_core_274;
  assign popcount38_u38d_out[2] = popcount38_u38d_core_279;
  assign popcount38_u38d_out[3] = popcount38_u38d_core_284;
  assign popcount38_u38d_out[4] = popcount38_u38d_core_286;
  assign popcount38_u38d_out[5] = 1'b0;
endmodule