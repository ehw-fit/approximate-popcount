// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.00019
// WCE=12.0
// EP=0.917529%
// Printed PDK parameters:
//  Area=21124698.0
//  Delay=40196880.0
//  Power=920570.0

module popcount24_cnyw(input [23:0] input_a, output [4:0] popcount24_cnyw_out);
  wire popcount24_cnyw_core_027;
  wire popcount24_cnyw_core_028_not;
  wire popcount24_cnyw_core_029;
  wire popcount24_cnyw_core_030;
  wire popcount24_cnyw_core_031;
  wire popcount24_cnyw_core_033;
  wire popcount24_cnyw_core_034;
  wire popcount24_cnyw_core_035;
  wire popcount24_cnyw_core_037;
  wire popcount24_cnyw_core_038;
  wire popcount24_cnyw_core_040;
  wire popcount24_cnyw_core_041;
  wire popcount24_cnyw_core_046;
  wire popcount24_cnyw_core_048;
  wire popcount24_cnyw_core_052;
  wire popcount24_cnyw_core_053;
  wire popcount24_cnyw_core_056;
  wire popcount24_cnyw_core_057;
  wire popcount24_cnyw_core_058;
  wire popcount24_cnyw_core_059;
  wire popcount24_cnyw_core_060;
  wire popcount24_cnyw_core_061;
  wire popcount24_cnyw_core_062;
  wire popcount24_cnyw_core_063;
  wire popcount24_cnyw_core_064_not;
  wire popcount24_cnyw_core_066;
  wire popcount24_cnyw_core_067;
  wire popcount24_cnyw_core_068;
  wire popcount24_cnyw_core_070;
  wire popcount24_cnyw_core_072;
  wire popcount24_cnyw_core_075;
  wire popcount24_cnyw_core_076;
  wire popcount24_cnyw_core_077;
  wire popcount24_cnyw_core_079;
  wire popcount24_cnyw_core_080;
  wire popcount24_cnyw_core_081;
  wire popcount24_cnyw_core_082;
  wire popcount24_cnyw_core_083;
  wire popcount24_cnyw_core_084;
  wire popcount24_cnyw_core_085;
  wire popcount24_cnyw_core_088;
  wire popcount24_cnyw_core_091;
  wire popcount24_cnyw_core_092;
  wire popcount24_cnyw_core_093;
  wire popcount24_cnyw_core_094;
  wire popcount24_cnyw_core_097;
  wire popcount24_cnyw_core_098;
  wire popcount24_cnyw_core_100;
  wire popcount24_cnyw_core_101;
  wire popcount24_cnyw_core_104;
  wire popcount24_cnyw_core_105;
  wire popcount24_cnyw_core_106;
  wire popcount24_cnyw_core_107;
  wire popcount24_cnyw_core_108;
  wire popcount24_cnyw_core_109;
  wire popcount24_cnyw_core_111;
  wire popcount24_cnyw_core_114;
  wire popcount24_cnyw_core_115;
  wire popcount24_cnyw_core_116;
  wire popcount24_cnyw_core_117;
  wire popcount24_cnyw_core_119;
  wire popcount24_cnyw_core_120;
  wire popcount24_cnyw_core_121;
  wire popcount24_cnyw_core_122_not;
  wire popcount24_cnyw_core_123;
  wire popcount24_cnyw_core_124_not;
  wire popcount24_cnyw_core_126;
  wire popcount24_cnyw_core_127;
  wire popcount24_cnyw_core_129;
  wire popcount24_cnyw_core_132;
  wire popcount24_cnyw_core_133_not;
  wire popcount24_cnyw_core_134;
  wire popcount24_cnyw_core_135;
  wire popcount24_cnyw_core_136;
  wire popcount24_cnyw_core_137;
  wire popcount24_cnyw_core_138;
  wire popcount24_cnyw_core_141;
  wire popcount24_cnyw_core_143;
  wire popcount24_cnyw_core_144;
  wire popcount24_cnyw_core_148;
  wire popcount24_cnyw_core_149;
  wire popcount24_cnyw_core_152;
  wire popcount24_cnyw_core_154;
  wire popcount24_cnyw_core_155;
  wire popcount24_cnyw_core_156;
  wire popcount24_cnyw_core_157;
  wire popcount24_cnyw_core_158;
  wire popcount24_cnyw_core_159;
  wire popcount24_cnyw_core_161;
  wire popcount24_cnyw_core_163;
  wire popcount24_cnyw_core_164;
  wire popcount24_cnyw_core_165;
  wire popcount24_cnyw_core_166;
  wire popcount24_cnyw_core_169;
  wire popcount24_cnyw_core_174;
  wire popcount24_cnyw_core_175;
  wire popcount24_cnyw_core_177;

  assign popcount24_cnyw_core_027 = input_a[8] & input_a[13];
  assign popcount24_cnyw_core_028_not = ~input_a[9];
  assign popcount24_cnyw_core_029 = input_a[21] & input_a[19];
  assign popcount24_cnyw_core_030 = popcount24_cnyw_core_027 | popcount24_cnyw_core_029;
  assign popcount24_cnyw_core_031 = ~(input_a[5] ^ input_a[5]);
  assign popcount24_cnyw_core_033 = input_a[22] & input_a[16];
  assign popcount24_cnyw_core_034 = ~(input_a[10] ^ input_a[9]);
  assign popcount24_cnyw_core_035 = ~(input_a[11] & input_a[8]);
  assign popcount24_cnyw_core_037 = ~(input_a[12] | input_a[9]);
  assign popcount24_cnyw_core_038 = ~(input_a[16] | input_a[8]);
  assign popcount24_cnyw_core_040 = popcount24_cnyw_core_030 ^ popcount24_cnyw_core_033;
  assign popcount24_cnyw_core_041 = popcount24_cnyw_core_030 & popcount24_cnyw_core_033;
  assign popcount24_cnyw_core_046 = input_a[5] ^ input_a[17];
  assign popcount24_cnyw_core_048 = input_a[1] | input_a[19];
  assign popcount24_cnyw_core_052 = ~(input_a[16] | input_a[0]);
  assign popcount24_cnyw_core_053 = ~input_a[23];
  assign popcount24_cnyw_core_056 = input_a[10] ^ input_a[11];
  assign popcount24_cnyw_core_057 = input_a[10] & input_a[11];
  assign popcount24_cnyw_core_058 = input_a[9] ^ popcount24_cnyw_core_056;
  assign popcount24_cnyw_core_059 = input_a[9] & popcount24_cnyw_core_056;
  assign popcount24_cnyw_core_060 = popcount24_cnyw_core_057 | popcount24_cnyw_core_059;
  assign popcount24_cnyw_core_061 = input_a[21] | input_a[5];
  assign popcount24_cnyw_core_062 = input_a[6] ^ popcount24_cnyw_core_058;
  assign popcount24_cnyw_core_063 = input_a[6] & popcount24_cnyw_core_058;
  assign popcount24_cnyw_core_064_not = ~popcount24_cnyw_core_060;
  assign popcount24_cnyw_core_066 = popcount24_cnyw_core_064_not ^ popcount24_cnyw_core_063;
  assign popcount24_cnyw_core_067 = input_a[6] & popcount24_cnyw_core_063;
  assign popcount24_cnyw_core_068 = popcount24_cnyw_core_060 | popcount24_cnyw_core_067;
  assign popcount24_cnyw_core_070 = ~input_a[14];
  assign popcount24_cnyw_core_072 = ~input_a[17];
  assign popcount24_cnyw_core_075 = input_a[0] & popcount24_cnyw_core_062;
  assign popcount24_cnyw_core_076 = popcount24_cnyw_core_040 | popcount24_cnyw_core_066;
  assign popcount24_cnyw_core_077 = popcount24_cnyw_core_040 & popcount24_cnyw_core_066;
  assign popcount24_cnyw_core_079 = popcount24_cnyw_core_076 & popcount24_cnyw_core_075;
  assign popcount24_cnyw_core_080 = popcount24_cnyw_core_077 | popcount24_cnyw_core_079;
  assign popcount24_cnyw_core_081 = popcount24_cnyw_core_041 ^ popcount24_cnyw_core_068;
  assign popcount24_cnyw_core_082 = popcount24_cnyw_core_041 & popcount24_cnyw_core_068;
  assign popcount24_cnyw_core_083 = popcount24_cnyw_core_081 ^ popcount24_cnyw_core_080;
  assign popcount24_cnyw_core_084 = popcount24_cnyw_core_081 & popcount24_cnyw_core_080;
  assign popcount24_cnyw_core_085 = popcount24_cnyw_core_082 | popcount24_cnyw_core_084;
  assign popcount24_cnyw_core_088 = input_a[23] | input_a[4];
  assign popcount24_cnyw_core_091 = ~(input_a[11] & input_a[2]);
  assign popcount24_cnyw_core_092 = input_a[7] & input_a[18];
  assign popcount24_cnyw_core_093 = input_a[5] | input_a[18];
  assign popcount24_cnyw_core_094 = input_a[3] | input_a[11];
  assign popcount24_cnyw_core_097 = input_a[18] | input_a[0];
  assign popcount24_cnyw_core_098 = input_a[23] & input_a[4];
  assign popcount24_cnyw_core_100 = input_a[12] & input_a[17];
  assign popcount24_cnyw_core_101 = popcount24_cnyw_core_098 | popcount24_cnyw_core_100;
  assign popcount24_cnyw_core_104 = input_a[1] & input_a[15];
  assign popcount24_cnyw_core_105 = popcount24_cnyw_core_092 ^ popcount24_cnyw_core_101;
  assign popcount24_cnyw_core_106 = popcount24_cnyw_core_092 & popcount24_cnyw_core_101;
  assign popcount24_cnyw_core_107 = popcount24_cnyw_core_105 ^ popcount24_cnyw_core_104;
  assign popcount24_cnyw_core_108 = popcount24_cnyw_core_105 & input_a[1];
  assign popcount24_cnyw_core_109 = popcount24_cnyw_core_106 | popcount24_cnyw_core_108;
  assign popcount24_cnyw_core_111 = input_a[2] | input_a[17];
  assign popcount24_cnyw_core_114 = ~input_a[4];
  assign popcount24_cnyw_core_115 = ~(input_a[6] | input_a[18]);
  assign popcount24_cnyw_core_116 = input_a[12] & input_a[19];
  assign popcount24_cnyw_core_117 = ~(input_a[14] | input_a[15]);
  assign popcount24_cnyw_core_119 = ~(input_a[4] ^ input_a[8]);
  assign popcount24_cnyw_core_120 = ~(input_a[9] & input_a[22]);
  assign popcount24_cnyw_core_121 = ~(input_a[5] & input_a[10]);
  assign popcount24_cnyw_core_122_not = ~input_a[6];
  assign popcount24_cnyw_core_123 = ~(input_a[18] | input_a[1]);
  assign popcount24_cnyw_core_124_not = ~input_a[6];
  assign popcount24_cnyw_core_126 = ~(input_a[15] ^ input_a[15]);
  assign popcount24_cnyw_core_127 = input_a[1] ^ input_a[6];
  assign popcount24_cnyw_core_129 = ~input_a[15];
  assign popcount24_cnyw_core_132 = input_a[3] & input_a[19];
  assign popcount24_cnyw_core_133_not = ~input_a[6];
  assign popcount24_cnyw_core_134 = input_a[7] | input_a[5];
  assign popcount24_cnyw_core_135 = ~(input_a[18] | input_a[12]);
  assign popcount24_cnyw_core_136 = input_a[15] | input_a[0];
  assign popcount24_cnyw_core_137 = ~(input_a[22] | input_a[13]);
  assign popcount24_cnyw_core_138 = input_a[13] & input_a[22];
  assign popcount24_cnyw_core_141 = ~(input_a[8] ^ input_a[6]);
  assign popcount24_cnyw_core_143 = ~(input_a[15] & input_a[0]);
  assign popcount24_cnyw_core_144 = input_a[15] | input_a[5];
  assign popcount24_cnyw_core_148 = popcount24_cnyw_core_109 ^ popcount24_cnyw_core_107;
  assign popcount24_cnyw_core_149 = popcount24_cnyw_core_109 & popcount24_cnyw_core_107;
  assign popcount24_cnyw_core_152 = input_a[5] | input_a[15];
  assign popcount24_cnyw_core_154 = input_a[3] ^ input_a[11];
  assign popcount24_cnyw_core_155 = input_a[3] ^ input_a[6];
  assign popcount24_cnyw_core_156 = ~(input_a[7] | input_a[17]);
  assign popcount24_cnyw_core_157 = ~(input_a[22] ^ input_a[5]);
  assign popcount24_cnyw_core_158 = ~(input_a[4] ^ input_a[6]);
  assign popcount24_cnyw_core_159 = input_a[22] & input_a[2];
  assign popcount24_cnyw_core_161 = input_a[3] & input_a[17];
  assign popcount24_cnyw_core_163 = popcount24_cnyw_core_083 | popcount24_cnyw_core_148;
  assign popcount24_cnyw_core_164 = popcount24_cnyw_core_083 & popcount24_cnyw_core_148;
  assign popcount24_cnyw_core_165 = input_a[4] ^ input_a[13];
  assign popcount24_cnyw_core_166 = ~(input_a[5] & input_a[21]);
  assign popcount24_cnyw_core_169 = input_a[15] & popcount24_cnyw_core_149;
  assign popcount24_cnyw_core_174 = input_a[18] | input_a[2];
  assign popcount24_cnyw_core_175 = popcount24_cnyw_core_085 | popcount24_cnyw_core_169;
  assign popcount24_cnyw_core_177 = ~(input_a[1] | input_a[13]);

  assign popcount24_cnyw_out[0] = input_a[20];
  assign popcount24_cnyw_out[1] = popcount24_cnyw_core_108;
  assign popcount24_cnyw_out[2] = popcount24_cnyw_core_163;
  assign popcount24_cnyw_out[3] = popcount24_cnyw_core_164;
  assign popcount24_cnyw_out[4] = popcount24_cnyw_core_175;
endmodule