// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=18.0278
// WCE=54.0
// EP=0.991483%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_flsk(input [38:0] input_a, output [5:0] popcount39_flsk_out);
  wire popcount39_flsk_core_041;
  wire popcount39_flsk_core_042;
  wire popcount39_flsk_core_044_not;
  wire popcount39_flsk_core_045;
  wire popcount39_flsk_core_048;
  wire popcount39_flsk_core_049;
  wire popcount39_flsk_core_050;
  wire popcount39_flsk_core_051;
  wire popcount39_flsk_core_053;
  wire popcount39_flsk_core_054;
  wire popcount39_flsk_core_055;
  wire popcount39_flsk_core_056;
  wire popcount39_flsk_core_058;
  wire popcount39_flsk_core_059;
  wire popcount39_flsk_core_060;
  wire popcount39_flsk_core_063;
  wire popcount39_flsk_core_064;
  wire popcount39_flsk_core_066;
  wire popcount39_flsk_core_067;
  wire popcount39_flsk_core_068;
  wire popcount39_flsk_core_069;
  wire popcount39_flsk_core_072;
  wire popcount39_flsk_core_073;
  wire popcount39_flsk_core_074;
  wire popcount39_flsk_core_075;
  wire popcount39_flsk_core_078;
  wire popcount39_flsk_core_079;
  wire popcount39_flsk_core_080;
  wire popcount39_flsk_core_081;
  wire popcount39_flsk_core_082;
  wire popcount39_flsk_core_083;
  wire popcount39_flsk_core_084;
  wire popcount39_flsk_core_085;
  wire popcount39_flsk_core_086;
  wire popcount39_flsk_core_088;
  wire popcount39_flsk_core_089;
  wire popcount39_flsk_core_090;
  wire popcount39_flsk_core_091;
  wire popcount39_flsk_core_093;
  wire popcount39_flsk_core_097;
  wire popcount39_flsk_core_098;
  wire popcount39_flsk_core_099;
  wire popcount39_flsk_core_100;
  wire popcount39_flsk_core_101;
  wire popcount39_flsk_core_102;
  wire popcount39_flsk_core_103;
  wire popcount39_flsk_core_104;
  wire popcount39_flsk_core_105;
  wire popcount39_flsk_core_106;
  wire popcount39_flsk_core_107;
  wire popcount39_flsk_core_108;
  wire popcount39_flsk_core_109;
  wire popcount39_flsk_core_110;
  wire popcount39_flsk_core_111;
  wire popcount39_flsk_core_114;
  wire popcount39_flsk_core_118;
  wire popcount39_flsk_core_122;
  wire popcount39_flsk_core_123;
  wire popcount39_flsk_core_124;
  wire popcount39_flsk_core_125;
  wire popcount39_flsk_core_127;
  wire popcount39_flsk_core_129;
  wire popcount39_flsk_core_130;
  wire popcount39_flsk_core_132;
  wire popcount39_flsk_core_135;
  wire popcount39_flsk_core_136;
  wire popcount39_flsk_core_137;
  wire popcount39_flsk_core_138;
  wire popcount39_flsk_core_140;
  wire popcount39_flsk_core_141;
  wire popcount39_flsk_core_142;
  wire popcount39_flsk_core_143;
  wire popcount39_flsk_core_145;
  wire popcount39_flsk_core_146;
  wire popcount39_flsk_core_149;
  wire popcount39_flsk_core_150;
  wire popcount39_flsk_core_152;
  wire popcount39_flsk_core_153;
  wire popcount39_flsk_core_154;
  wire popcount39_flsk_core_155;
  wire popcount39_flsk_core_157;
  wire popcount39_flsk_core_158;
  wire popcount39_flsk_core_160_not;
  wire popcount39_flsk_core_161;
  wire popcount39_flsk_core_162;
  wire popcount39_flsk_core_163;
  wire popcount39_flsk_core_165;
  wire popcount39_flsk_core_166;
  wire popcount39_flsk_core_168;
  wire popcount39_flsk_core_170;
  wire popcount39_flsk_core_171;
  wire popcount39_flsk_core_172;
  wire popcount39_flsk_core_173;
  wire popcount39_flsk_core_174;
  wire popcount39_flsk_core_177;
  wire popcount39_flsk_core_179;
  wire popcount39_flsk_core_183;
  wire popcount39_flsk_core_185;
  wire popcount39_flsk_core_186;
  wire popcount39_flsk_core_187;
  wire popcount39_flsk_core_191;
  wire popcount39_flsk_core_192;
  wire popcount39_flsk_core_195;
  wire popcount39_flsk_core_196;
  wire popcount39_flsk_core_197;
  wire popcount39_flsk_core_200;
  wire popcount39_flsk_core_203;
  wire popcount39_flsk_core_204;
  wire popcount39_flsk_core_205;
  wire popcount39_flsk_core_207;
  wire popcount39_flsk_core_209;
  wire popcount39_flsk_core_210;
  wire popcount39_flsk_core_212;
  wire popcount39_flsk_core_215;
  wire popcount39_flsk_core_216;
  wire popcount39_flsk_core_218;
  wire popcount39_flsk_core_221;
  wire popcount39_flsk_core_222;
  wire popcount39_flsk_core_224;
  wire popcount39_flsk_core_225;
  wire popcount39_flsk_core_227;
  wire popcount39_flsk_core_229;
  wire popcount39_flsk_core_230;
  wire popcount39_flsk_core_231;
  wire popcount39_flsk_core_232;
  wire popcount39_flsk_core_233;
  wire popcount39_flsk_core_234;
  wire popcount39_flsk_core_235;
  wire popcount39_flsk_core_236;
  wire popcount39_flsk_core_238;
  wire popcount39_flsk_core_240;
  wire popcount39_flsk_core_242;
  wire popcount39_flsk_core_243;
  wire popcount39_flsk_core_245;
  wire popcount39_flsk_core_247;
  wire popcount39_flsk_core_248;
  wire popcount39_flsk_core_249;
  wire popcount39_flsk_core_252;
  wire popcount39_flsk_core_253;
  wire popcount39_flsk_core_254;
  wire popcount39_flsk_core_255;
  wire popcount39_flsk_core_256;
  wire popcount39_flsk_core_257;
  wire popcount39_flsk_core_258;
  wire popcount39_flsk_core_259;
  wire popcount39_flsk_core_260;
  wire popcount39_flsk_core_261;
  wire popcount39_flsk_core_263;
  wire popcount39_flsk_core_265;
  wire popcount39_flsk_core_269;
  wire popcount39_flsk_core_270;
  wire popcount39_flsk_core_271;
  wire popcount39_flsk_core_273;
  wire popcount39_flsk_core_274;
  wire popcount39_flsk_core_275;
  wire popcount39_flsk_core_276;
  wire popcount39_flsk_core_277;
  wire popcount39_flsk_core_279;
  wire popcount39_flsk_core_280;
  wire popcount39_flsk_core_281_not;
  wire popcount39_flsk_core_282;
  wire popcount39_flsk_core_283;
  wire popcount39_flsk_core_284;
  wire popcount39_flsk_core_285;
  wire popcount39_flsk_core_286;
  wire popcount39_flsk_core_288;
  wire popcount39_flsk_core_289;
  wire popcount39_flsk_core_292;
  wire popcount39_flsk_core_295;
  wire popcount39_flsk_core_296;
  wire popcount39_flsk_core_297;
  wire popcount39_flsk_core_299;
  wire popcount39_flsk_core_300;
  wire popcount39_flsk_core_301;
  wire popcount39_flsk_core_304;

  assign popcount39_flsk_core_041 = ~(input_a[1] ^ input_a[24]);
  assign popcount39_flsk_core_042 = ~(input_a[9] ^ input_a[15]);
  assign popcount39_flsk_core_044_not = ~input_a[18];
  assign popcount39_flsk_core_045 = ~(input_a[32] ^ input_a[16]);
  assign popcount39_flsk_core_048 = input_a[36] ^ input_a[26];
  assign popcount39_flsk_core_049 = ~(input_a[36] | input_a[17]);
  assign popcount39_flsk_core_050 = input_a[11] & input_a[9];
  assign popcount39_flsk_core_051 = input_a[30] ^ input_a[18];
  assign popcount39_flsk_core_053 = input_a[37] ^ input_a[33];
  assign popcount39_flsk_core_054 = ~input_a[26];
  assign popcount39_flsk_core_055 = input_a[11] ^ input_a[34];
  assign popcount39_flsk_core_056 = input_a[38] | input_a[34];
  assign popcount39_flsk_core_058 = input_a[4] ^ input_a[35];
  assign popcount39_flsk_core_059 = input_a[34] & input_a[16];
  assign popcount39_flsk_core_060 = input_a[2] & input_a[2];
  assign popcount39_flsk_core_063 = input_a[21] ^ input_a[32];
  assign popcount39_flsk_core_064 = input_a[27] | input_a[11];
  assign popcount39_flsk_core_066 = input_a[0] ^ input_a[7];
  assign popcount39_flsk_core_067 = ~input_a[34];
  assign popcount39_flsk_core_068 = ~(input_a[9] & input_a[10]);
  assign popcount39_flsk_core_069 = ~input_a[24];
  assign popcount39_flsk_core_072 = ~(input_a[5] | input_a[7]);
  assign popcount39_flsk_core_073 = input_a[20] | input_a[19];
  assign popcount39_flsk_core_074 = input_a[16] ^ input_a[3];
  assign popcount39_flsk_core_075 = ~(input_a[6] | input_a[13]);
  assign popcount39_flsk_core_078 = ~(input_a[12] ^ input_a[34]);
  assign popcount39_flsk_core_079 = input_a[34] & input_a[33];
  assign popcount39_flsk_core_080 = input_a[22] | input_a[27];
  assign popcount39_flsk_core_081 = ~(input_a[38] | input_a[36]);
  assign popcount39_flsk_core_082 = ~(input_a[31] | input_a[5]);
  assign popcount39_flsk_core_083 = input_a[28] ^ input_a[31];
  assign popcount39_flsk_core_084 = ~(input_a[22] | input_a[3]);
  assign popcount39_flsk_core_085 = ~input_a[15];
  assign popcount39_flsk_core_086 = ~(input_a[38] ^ input_a[6]);
  assign popcount39_flsk_core_088 = ~(input_a[34] & input_a[25]);
  assign popcount39_flsk_core_089 = ~input_a[21];
  assign popcount39_flsk_core_090 = ~input_a[12];
  assign popcount39_flsk_core_091 = input_a[22] | input_a[18];
  assign popcount39_flsk_core_093 = ~(input_a[12] ^ input_a[37]);
  assign popcount39_flsk_core_097 = input_a[17] ^ input_a[21];
  assign popcount39_flsk_core_098 = ~(input_a[17] ^ input_a[1]);
  assign popcount39_flsk_core_099 = ~input_a[7];
  assign popcount39_flsk_core_100 = input_a[9] ^ input_a[4];
  assign popcount39_flsk_core_101 = ~(input_a[10] | input_a[14]);
  assign popcount39_flsk_core_102 = input_a[18] | input_a[18];
  assign popcount39_flsk_core_103 = input_a[37] & input_a[30];
  assign popcount39_flsk_core_104 = input_a[17] | input_a[33];
  assign popcount39_flsk_core_105 = input_a[17] & input_a[7];
  assign popcount39_flsk_core_106 = input_a[14] ^ input_a[1];
  assign popcount39_flsk_core_107 = input_a[11] & input_a[9];
  assign popcount39_flsk_core_108 = ~(input_a[13] | input_a[15]);
  assign popcount39_flsk_core_109 = ~(input_a[19] | input_a[10]);
  assign popcount39_flsk_core_110 = input_a[37] ^ input_a[1];
  assign popcount39_flsk_core_111 = ~input_a[4];
  assign popcount39_flsk_core_114 = input_a[32] | input_a[19];
  assign popcount39_flsk_core_118 = ~input_a[10];
  assign popcount39_flsk_core_122 = ~(input_a[26] & input_a[16]);
  assign popcount39_flsk_core_123 = ~(input_a[3] | input_a[15]);
  assign popcount39_flsk_core_124 = ~(input_a[29] | input_a[36]);
  assign popcount39_flsk_core_125 = input_a[16] & input_a[17];
  assign popcount39_flsk_core_127 = ~(input_a[35] | input_a[23]);
  assign popcount39_flsk_core_129 = ~(input_a[26] ^ input_a[14]);
  assign popcount39_flsk_core_130 = input_a[32] & input_a[3];
  assign popcount39_flsk_core_132 = input_a[30] ^ input_a[16];
  assign popcount39_flsk_core_135 = ~input_a[29];
  assign popcount39_flsk_core_136 = input_a[29] | input_a[3];
  assign popcount39_flsk_core_137 = ~(input_a[35] | input_a[32]);
  assign popcount39_flsk_core_138 = input_a[28] & input_a[28];
  assign popcount39_flsk_core_140 = ~(input_a[30] & input_a[6]);
  assign popcount39_flsk_core_141 = ~(input_a[4] & input_a[18]);
  assign popcount39_flsk_core_142 = ~(input_a[35] | input_a[10]);
  assign popcount39_flsk_core_143 = ~(input_a[38] | input_a[11]);
  assign popcount39_flsk_core_145 = ~(input_a[33] | input_a[32]);
  assign popcount39_flsk_core_146 = ~(input_a[26] & input_a[4]);
  assign popcount39_flsk_core_149 = ~input_a[28];
  assign popcount39_flsk_core_150 = input_a[24] | input_a[29];
  assign popcount39_flsk_core_152 = input_a[16] | input_a[21];
  assign popcount39_flsk_core_153 = ~(input_a[38] ^ input_a[12]);
  assign popcount39_flsk_core_154 = ~(input_a[33] | input_a[0]);
  assign popcount39_flsk_core_155 = ~(input_a[29] | input_a[38]);
  assign popcount39_flsk_core_157 = input_a[1] ^ input_a[13];
  assign popcount39_flsk_core_158 = input_a[21] ^ input_a[10];
  assign popcount39_flsk_core_160_not = ~input_a[19];
  assign popcount39_flsk_core_161 = ~input_a[13];
  assign popcount39_flsk_core_162 = ~input_a[19];
  assign popcount39_flsk_core_163 = ~(input_a[8] & input_a[37]);
  assign popcount39_flsk_core_165 = ~(input_a[29] & input_a[11]);
  assign popcount39_flsk_core_166 = input_a[31] | input_a[19];
  assign popcount39_flsk_core_168 = ~(input_a[27] & input_a[37]);
  assign popcount39_flsk_core_170 = ~(input_a[19] & input_a[30]);
  assign popcount39_flsk_core_171 = input_a[29] ^ input_a[25];
  assign popcount39_flsk_core_172 = input_a[34] & input_a[7];
  assign popcount39_flsk_core_173 = ~(input_a[18] & input_a[7]);
  assign popcount39_flsk_core_174 = input_a[36] & input_a[32];
  assign popcount39_flsk_core_177 = ~(input_a[15] | input_a[5]);
  assign popcount39_flsk_core_179 = input_a[21] ^ input_a[14];
  assign popcount39_flsk_core_183 = ~(input_a[15] & input_a[15]);
  assign popcount39_flsk_core_185 = ~(input_a[19] ^ input_a[23]);
  assign popcount39_flsk_core_186 = input_a[25] | input_a[14];
  assign popcount39_flsk_core_187 = ~(input_a[9] ^ input_a[20]);
  assign popcount39_flsk_core_191 = ~(input_a[13] | input_a[31]);
  assign popcount39_flsk_core_192 = input_a[5] | input_a[9];
  assign popcount39_flsk_core_195 = ~(input_a[28] ^ input_a[32]);
  assign popcount39_flsk_core_196 = input_a[22] | input_a[37];
  assign popcount39_flsk_core_197 = ~(input_a[15] | input_a[10]);
  assign popcount39_flsk_core_200 = input_a[15] | input_a[12];
  assign popcount39_flsk_core_203 = input_a[37] | input_a[37];
  assign popcount39_flsk_core_204 = ~(input_a[25] & input_a[13]);
  assign popcount39_flsk_core_205 = ~(input_a[30] & input_a[7]);
  assign popcount39_flsk_core_207 = ~input_a[20];
  assign popcount39_flsk_core_209 = input_a[20] | input_a[21];
  assign popcount39_flsk_core_210 = ~(input_a[32] ^ input_a[17]);
  assign popcount39_flsk_core_212 = ~(input_a[33] ^ input_a[17]);
  assign popcount39_flsk_core_215 = input_a[14] ^ input_a[22];
  assign popcount39_flsk_core_216 = input_a[23] | input_a[34];
  assign popcount39_flsk_core_218 = ~input_a[34];
  assign popcount39_flsk_core_221 = ~(input_a[30] & input_a[16]);
  assign popcount39_flsk_core_222 = input_a[14] ^ input_a[15];
  assign popcount39_flsk_core_224 = ~(input_a[9] & input_a[17]);
  assign popcount39_flsk_core_225 = ~input_a[16];
  assign popcount39_flsk_core_227 = input_a[36] ^ input_a[3];
  assign popcount39_flsk_core_229 = input_a[5] ^ input_a[17];
  assign popcount39_flsk_core_230 = ~(input_a[5] | input_a[7]);
  assign popcount39_flsk_core_231 = ~(input_a[0] & input_a[38]);
  assign popcount39_flsk_core_232 = ~(input_a[28] & input_a[14]);
  assign popcount39_flsk_core_233 = input_a[27] & input_a[25];
  assign popcount39_flsk_core_234 = ~input_a[27];
  assign popcount39_flsk_core_235 = input_a[28] ^ input_a[20];
  assign popcount39_flsk_core_236 = input_a[29] | input_a[18];
  assign popcount39_flsk_core_238 = input_a[5] ^ input_a[37];
  assign popcount39_flsk_core_240 = ~input_a[32];
  assign popcount39_flsk_core_242 = ~(input_a[33] | input_a[29]);
  assign popcount39_flsk_core_243 = input_a[28] & input_a[34];
  assign popcount39_flsk_core_245 = ~input_a[0];
  assign popcount39_flsk_core_247 = input_a[4] ^ input_a[5];
  assign popcount39_flsk_core_248 = input_a[20] ^ input_a[27];
  assign popcount39_flsk_core_249 = input_a[2] & input_a[4];
  assign popcount39_flsk_core_252 = input_a[6] | input_a[23];
  assign popcount39_flsk_core_253 = input_a[0] ^ input_a[33];
  assign popcount39_flsk_core_254 = input_a[6] | input_a[22];
  assign popcount39_flsk_core_255 = input_a[6] | input_a[4];
  assign popcount39_flsk_core_256 = input_a[14] & input_a[8];
  assign popcount39_flsk_core_257 = ~(input_a[26] ^ input_a[5]);
  assign popcount39_flsk_core_258 = ~(input_a[14] & input_a[8]);
  assign popcount39_flsk_core_259 = ~(input_a[17] & input_a[0]);
  assign popcount39_flsk_core_260 = ~(input_a[31] & input_a[8]);
  assign popcount39_flsk_core_261 = input_a[6] | input_a[25];
  assign popcount39_flsk_core_263 = ~input_a[10];
  assign popcount39_flsk_core_265 = ~input_a[31];
  assign popcount39_flsk_core_269 = input_a[28] ^ input_a[27];
  assign popcount39_flsk_core_270 = ~(input_a[33] & input_a[32]);
  assign popcount39_flsk_core_271 = ~(input_a[32] | input_a[3]);
  assign popcount39_flsk_core_273 = input_a[18] ^ input_a[23];
  assign popcount39_flsk_core_274 = input_a[14] & input_a[24];
  assign popcount39_flsk_core_275 = ~(input_a[4] ^ input_a[36]);
  assign popcount39_flsk_core_276 = input_a[24] ^ input_a[3];
  assign popcount39_flsk_core_277 = ~(input_a[23] | input_a[6]);
  assign popcount39_flsk_core_279 = ~(input_a[29] ^ input_a[33]);
  assign popcount39_flsk_core_280 = ~(input_a[23] ^ input_a[27]);
  assign popcount39_flsk_core_281_not = ~input_a[3];
  assign popcount39_flsk_core_282 = input_a[38] ^ input_a[7];
  assign popcount39_flsk_core_283 = ~(input_a[31] ^ input_a[29]);
  assign popcount39_flsk_core_284 = ~input_a[35];
  assign popcount39_flsk_core_285 = ~(input_a[0] | input_a[25]);
  assign popcount39_flsk_core_286 = ~(input_a[4] ^ input_a[35]);
  assign popcount39_flsk_core_288 = input_a[9] | input_a[6];
  assign popcount39_flsk_core_289 = input_a[22] | input_a[17];
  assign popcount39_flsk_core_292 = ~(input_a[25] ^ input_a[31]);
  assign popcount39_flsk_core_295 = ~(input_a[30] & input_a[34]);
  assign popcount39_flsk_core_296 = ~(input_a[21] & input_a[27]);
  assign popcount39_flsk_core_297 = input_a[17] | input_a[0];
  assign popcount39_flsk_core_299 = ~(input_a[18] & input_a[24]);
  assign popcount39_flsk_core_300 = ~input_a[14];
  assign popcount39_flsk_core_301 = ~(input_a[26] | input_a[25]);
  assign popcount39_flsk_core_304 = input_a[31] ^ input_a[4];

  assign popcount39_flsk_out[0] = input_a[9];
  assign popcount39_flsk_out[1] = 1'b0;
  assign popcount39_flsk_out[2] = 1'b0;
  assign popcount39_flsk_out[3] = 1'b1;
  assign popcount39_flsk_out[4] = input_a[29];
  assign popcount39_flsk_out[5] = input_a[28];
endmodule