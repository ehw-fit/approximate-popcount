// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.84216
// WCE=31.0
// EP=0.967491%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount36_9tg7(input [35:0] input_a, output [5:0] popcount36_9tg7_out);
  wire popcount36_9tg7_core_038;
  wire popcount36_9tg7_core_039_not;
  wire popcount36_9tg7_core_040;
  wire popcount36_9tg7_core_041;
  wire popcount36_9tg7_core_043;
  wire popcount36_9tg7_core_046;
  wire popcount36_9tg7_core_047;
  wire popcount36_9tg7_core_048;
  wire popcount36_9tg7_core_050;
  wire popcount36_9tg7_core_051;
  wire popcount36_9tg7_core_053;
  wire popcount36_9tg7_core_054;
  wire popcount36_9tg7_core_055;
  wire popcount36_9tg7_core_056;
  wire popcount36_9tg7_core_057;
  wire popcount36_9tg7_core_058;
  wire popcount36_9tg7_core_059;
  wire popcount36_9tg7_core_065;
  wire popcount36_9tg7_core_066;
  wire popcount36_9tg7_core_067;
  wire popcount36_9tg7_core_071;
  wire popcount36_9tg7_core_072;
  wire popcount36_9tg7_core_075;
  wire popcount36_9tg7_core_076;
  wire popcount36_9tg7_core_077;
  wire popcount36_9tg7_core_079;
  wire popcount36_9tg7_core_080;
  wire popcount36_9tg7_core_084;
  wire popcount36_9tg7_core_085;
  wire popcount36_9tg7_core_087;
  wire popcount36_9tg7_core_089;
  wire popcount36_9tg7_core_090;
  wire popcount36_9tg7_core_091;
  wire popcount36_9tg7_core_092;
  wire popcount36_9tg7_core_093;
  wire popcount36_9tg7_core_098;
  wire popcount36_9tg7_core_100;
  wire popcount36_9tg7_core_103;
  wire popcount36_9tg7_core_104;
  wire popcount36_9tg7_core_105_not;
  wire popcount36_9tg7_core_107;
  wire popcount36_9tg7_core_108;
  wire popcount36_9tg7_core_110;
  wire popcount36_9tg7_core_111;
  wire popcount36_9tg7_core_112;
  wire popcount36_9tg7_core_113;
  wire popcount36_9tg7_core_114;
  wire popcount36_9tg7_core_115;
  wire popcount36_9tg7_core_118;
  wire popcount36_9tg7_core_120;
  wire popcount36_9tg7_core_121;
  wire popcount36_9tg7_core_123;
  wire popcount36_9tg7_core_125;
  wire popcount36_9tg7_core_126;
  wire popcount36_9tg7_core_127;
  wire popcount36_9tg7_core_128;
  wire popcount36_9tg7_core_129;
  wire popcount36_9tg7_core_130;
  wire popcount36_9tg7_core_132;
  wire popcount36_9tg7_core_133;
  wire popcount36_9tg7_core_135;
  wire popcount36_9tg7_core_136;
  wire popcount36_9tg7_core_139;
  wire popcount36_9tg7_core_140;
  wire popcount36_9tg7_core_142;
  wire popcount36_9tg7_core_143;
  wire popcount36_9tg7_core_144;
  wire popcount36_9tg7_core_147_not;
  wire popcount36_9tg7_core_148;
  wire popcount36_9tg7_core_151;
  wire popcount36_9tg7_core_152;
  wire popcount36_9tg7_core_153;
  wire popcount36_9tg7_core_154;
  wire popcount36_9tg7_core_155;
  wire popcount36_9tg7_core_156;
  wire popcount36_9tg7_core_157;
  wire popcount36_9tg7_core_158;
  wire popcount36_9tg7_core_159;
  wire popcount36_9tg7_core_160;
  wire popcount36_9tg7_core_161;
  wire popcount36_9tg7_core_162;
  wire popcount36_9tg7_core_163;
  wire popcount36_9tg7_core_164;
  wire popcount36_9tg7_core_165;
  wire popcount36_9tg7_core_167_not;
  wire popcount36_9tg7_core_168;
  wire popcount36_9tg7_core_169;
  wire popcount36_9tg7_core_170;
  wire popcount36_9tg7_core_172;
  wire popcount36_9tg7_core_175;
  wire popcount36_9tg7_core_176;
  wire popcount36_9tg7_core_177;
  wire popcount36_9tg7_core_178_not;
  wire popcount36_9tg7_core_181;
  wire popcount36_9tg7_core_182;
  wire popcount36_9tg7_core_183;
  wire popcount36_9tg7_core_184;
  wire popcount36_9tg7_core_185;
  wire popcount36_9tg7_core_186;
  wire popcount36_9tg7_core_189;
  wire popcount36_9tg7_core_190_not;
  wire popcount36_9tg7_core_192;
  wire popcount36_9tg7_core_193;
  wire popcount36_9tg7_core_194;
  wire popcount36_9tg7_core_195;
  wire popcount36_9tg7_core_196;
  wire popcount36_9tg7_core_197;
  wire popcount36_9tg7_core_199;
  wire popcount36_9tg7_core_200;
  wire popcount36_9tg7_core_201;
  wire popcount36_9tg7_core_202;
  wire popcount36_9tg7_core_203;
  wire popcount36_9tg7_core_204;
  wire popcount36_9tg7_core_205;
  wire popcount36_9tg7_core_206;
  wire popcount36_9tg7_core_208;
  wire popcount36_9tg7_core_210;
  wire popcount36_9tg7_core_212;
  wire popcount36_9tg7_core_214;
  wire popcount36_9tg7_core_216;
  wire popcount36_9tg7_core_218;
  wire popcount36_9tg7_core_220;
  wire popcount36_9tg7_core_221;
  wire popcount36_9tg7_core_222;
  wire popcount36_9tg7_core_224;
  wire popcount36_9tg7_core_225;
  wire popcount36_9tg7_core_227;
  wire popcount36_9tg7_core_230;
  wire popcount36_9tg7_core_232;
  wire popcount36_9tg7_core_234;
  wire popcount36_9tg7_core_236;
  wire popcount36_9tg7_core_237;
  wire popcount36_9tg7_core_238;
  wire popcount36_9tg7_core_239;
  wire popcount36_9tg7_core_244;
  wire popcount36_9tg7_core_245;
  wire popcount36_9tg7_core_246;
  wire popcount36_9tg7_core_249;
  wire popcount36_9tg7_core_251;
  wire popcount36_9tg7_core_256;
  wire popcount36_9tg7_core_258;
  wire popcount36_9tg7_core_259;
  wire popcount36_9tg7_core_261;
  wire popcount36_9tg7_core_262;
  wire popcount36_9tg7_core_263_not;
  wire popcount36_9tg7_core_264;
  wire popcount36_9tg7_core_265;
  wire popcount36_9tg7_core_267;
  wire popcount36_9tg7_core_268;
  wire popcount36_9tg7_core_270;
  wire popcount36_9tg7_core_272;
  wire popcount36_9tg7_core_273;
  wire popcount36_9tg7_core_274;
  wire popcount36_9tg7_core_275;
  wire popcount36_9tg7_core_276;

  assign popcount36_9tg7_core_038 = ~(input_a[21] & input_a[0]);
  assign popcount36_9tg7_core_039_not = ~input_a[9];
  assign popcount36_9tg7_core_040 = input_a[18] | input_a[7];
  assign popcount36_9tg7_core_041 = ~(input_a[16] | input_a[4]);
  assign popcount36_9tg7_core_043 = input_a[26] & input_a[9];
  assign popcount36_9tg7_core_046 = ~(input_a[35] & input_a[16]);
  assign popcount36_9tg7_core_047 = input_a[18] ^ input_a[16];
  assign popcount36_9tg7_core_048 = ~(input_a[27] & input_a[18]);
  assign popcount36_9tg7_core_050 = input_a[10] ^ input_a[31];
  assign popcount36_9tg7_core_051 = ~(input_a[10] ^ input_a[31]);
  assign popcount36_9tg7_core_053 = ~(input_a[29] ^ input_a[24]);
  assign popcount36_9tg7_core_054 = input_a[5] | input_a[22];
  assign popcount36_9tg7_core_055 = input_a[3] | input_a[19];
  assign popcount36_9tg7_core_056 = ~(input_a[34] | input_a[0]);
  assign popcount36_9tg7_core_057 = input_a[22] ^ input_a[31];
  assign popcount36_9tg7_core_058 = input_a[2] ^ input_a[33];
  assign popcount36_9tg7_core_059 = input_a[34] ^ input_a[1];
  assign popcount36_9tg7_core_065 = input_a[11] ^ input_a[16];
  assign popcount36_9tg7_core_066 = ~(input_a[16] & input_a[2]);
  assign popcount36_9tg7_core_067 = input_a[13] ^ input_a[14];
  assign popcount36_9tg7_core_071 = input_a[4] & input_a[15];
  assign popcount36_9tg7_core_072 = input_a[17] & input_a[20];
  assign popcount36_9tg7_core_075 = input_a[30] | input_a[18];
  assign popcount36_9tg7_core_076 = ~(input_a[35] & input_a[14]);
  assign popcount36_9tg7_core_077 = ~(input_a[9] & input_a[5]);
  assign popcount36_9tg7_core_079 = input_a[24] ^ input_a[24];
  assign popcount36_9tg7_core_080 = input_a[22] & input_a[16];
  assign popcount36_9tg7_core_084 = ~(input_a[7] | input_a[8]);
  assign popcount36_9tg7_core_085 = ~(input_a[11] & input_a[22]);
  assign popcount36_9tg7_core_087 = input_a[34] & input_a[26];
  assign popcount36_9tg7_core_089 = ~input_a[13];
  assign popcount36_9tg7_core_090 = ~(input_a[19] | input_a[3]);
  assign popcount36_9tg7_core_091 = input_a[11] ^ input_a[4];
  assign popcount36_9tg7_core_092 = input_a[2] | input_a[3];
  assign popcount36_9tg7_core_093 = input_a[33] ^ input_a[4];
  assign popcount36_9tg7_core_098 = input_a[14] | input_a[26];
  assign popcount36_9tg7_core_100 = ~(input_a[24] & input_a[21]);
  assign popcount36_9tg7_core_103 = input_a[4] & input_a[26];
  assign popcount36_9tg7_core_104 = ~(input_a[26] | input_a[4]);
  assign popcount36_9tg7_core_105_not = ~input_a[12];
  assign popcount36_9tg7_core_107 = ~input_a[32];
  assign popcount36_9tg7_core_108 = ~(input_a[17] ^ input_a[13]);
  assign popcount36_9tg7_core_110 = ~(input_a[17] & input_a[26]);
  assign popcount36_9tg7_core_111 = ~(input_a[27] & input_a[16]);
  assign popcount36_9tg7_core_112 = input_a[19] ^ input_a[20];
  assign popcount36_9tg7_core_113 = ~(input_a[3] | input_a[31]);
  assign popcount36_9tg7_core_114 = ~input_a[4];
  assign popcount36_9tg7_core_115 = input_a[4] | input_a[23];
  assign popcount36_9tg7_core_118 = ~(input_a[25] & input_a[9]);
  assign popcount36_9tg7_core_120 = input_a[15] ^ input_a[8];
  assign popcount36_9tg7_core_121 = ~input_a[11];
  assign popcount36_9tg7_core_123 = input_a[21] & input_a[6];
  assign popcount36_9tg7_core_125 = input_a[17] ^ input_a[34];
  assign popcount36_9tg7_core_126 = ~(input_a[18] & input_a[18]);
  assign popcount36_9tg7_core_127 = ~(input_a[1] | input_a[12]);
  assign popcount36_9tg7_core_128 = input_a[34] & input_a[9];
  assign popcount36_9tg7_core_129 = input_a[9] | input_a[31];
  assign popcount36_9tg7_core_130 = ~(input_a[15] & input_a[8]);
  assign popcount36_9tg7_core_132 = input_a[10] | input_a[14];
  assign popcount36_9tg7_core_133 = input_a[33] & input_a[12];
  assign popcount36_9tg7_core_135 = ~(input_a[5] ^ input_a[15]);
  assign popcount36_9tg7_core_136 = ~(input_a[13] | input_a[10]);
  assign popcount36_9tg7_core_139 = input_a[1] & input_a[6];
  assign popcount36_9tg7_core_140 = ~(input_a[20] & input_a[31]);
  assign popcount36_9tg7_core_142 = input_a[29] | input_a[33];
  assign popcount36_9tg7_core_143 = ~(input_a[34] & input_a[11]);
  assign popcount36_9tg7_core_144 = input_a[14] & input_a[5];
  assign popcount36_9tg7_core_147_not = ~input_a[28];
  assign popcount36_9tg7_core_148 = input_a[35] & input_a[0];
  assign popcount36_9tg7_core_151 = input_a[5] | input_a[7];
  assign popcount36_9tg7_core_152 = input_a[23] ^ input_a[9];
  assign popcount36_9tg7_core_153 = input_a[9] ^ input_a[19];
  assign popcount36_9tg7_core_154 = ~(input_a[1] ^ input_a[1]);
  assign popcount36_9tg7_core_155 = ~input_a[29];
  assign popcount36_9tg7_core_156 = input_a[30] ^ input_a[11];
  assign popcount36_9tg7_core_157 = input_a[9] ^ input_a[10];
  assign popcount36_9tg7_core_158 = input_a[31] ^ input_a[33];
  assign popcount36_9tg7_core_159 = input_a[22] ^ input_a[29];
  assign popcount36_9tg7_core_160 = ~(input_a[2] ^ input_a[26]);
  assign popcount36_9tg7_core_161 = ~(input_a[25] ^ input_a[1]);
  assign popcount36_9tg7_core_162 = input_a[3] & input_a[18];
  assign popcount36_9tg7_core_163 = ~input_a[16];
  assign popcount36_9tg7_core_164 = ~input_a[6];
  assign popcount36_9tg7_core_165 = ~(input_a[11] & input_a[7]);
  assign popcount36_9tg7_core_167_not = ~input_a[21];
  assign popcount36_9tg7_core_168 = ~input_a[19];
  assign popcount36_9tg7_core_169 = ~input_a[24];
  assign popcount36_9tg7_core_170 = ~(input_a[16] ^ input_a[34]);
  assign popcount36_9tg7_core_172 = ~(input_a[16] & input_a[28]);
  assign popcount36_9tg7_core_175 = ~(input_a[8] ^ input_a[7]);
  assign popcount36_9tg7_core_176 = input_a[20] ^ input_a[7];
  assign popcount36_9tg7_core_177 = ~(input_a[16] ^ input_a[17]);
  assign popcount36_9tg7_core_178_not = ~input_a[18];
  assign popcount36_9tg7_core_181 = ~(input_a[2] | input_a[4]);
  assign popcount36_9tg7_core_182 = input_a[29] ^ input_a[11];
  assign popcount36_9tg7_core_183 = input_a[5] ^ input_a[14];
  assign popcount36_9tg7_core_184 = input_a[30] | input_a[23];
  assign popcount36_9tg7_core_185 = ~(input_a[11] ^ input_a[31]);
  assign popcount36_9tg7_core_186 = ~(input_a[0] | input_a[8]);
  assign popcount36_9tg7_core_189 = ~input_a[31];
  assign popcount36_9tg7_core_190_not = ~input_a[27];
  assign popcount36_9tg7_core_192 = input_a[12] & input_a[9];
  assign popcount36_9tg7_core_193 = ~(input_a[15] ^ input_a[3]);
  assign popcount36_9tg7_core_194 = input_a[20] | input_a[23];
  assign popcount36_9tg7_core_195 = input_a[1] & input_a[31];
  assign popcount36_9tg7_core_196 = ~(input_a[8] | input_a[32]);
  assign popcount36_9tg7_core_197 = ~(input_a[2] | input_a[35]);
  assign popcount36_9tg7_core_199 = ~input_a[19];
  assign popcount36_9tg7_core_200 = ~(input_a[31] & input_a[29]);
  assign popcount36_9tg7_core_201 = input_a[4] | input_a[9];
  assign popcount36_9tg7_core_202 = input_a[22] ^ input_a[27];
  assign popcount36_9tg7_core_203 = ~(input_a[5] & input_a[23]);
  assign popcount36_9tg7_core_204 = ~(input_a[18] ^ input_a[0]);
  assign popcount36_9tg7_core_205 = ~(input_a[29] & input_a[17]);
  assign popcount36_9tg7_core_206 = ~(input_a[15] | input_a[4]);
  assign popcount36_9tg7_core_208 = input_a[35] & input_a[22];
  assign popcount36_9tg7_core_210 = ~(input_a[33] & input_a[21]);
  assign popcount36_9tg7_core_212 = ~(input_a[16] | input_a[15]);
  assign popcount36_9tg7_core_214 = ~(input_a[9] ^ input_a[2]);
  assign popcount36_9tg7_core_216 = input_a[0] ^ input_a[20];
  assign popcount36_9tg7_core_218 = input_a[32] & input_a[20];
  assign popcount36_9tg7_core_220 = ~(input_a[18] & input_a[27]);
  assign popcount36_9tg7_core_221 = ~(input_a[34] & input_a[34]);
  assign popcount36_9tg7_core_222 = ~(input_a[30] & input_a[32]);
  assign popcount36_9tg7_core_224 = input_a[28] | input_a[3];
  assign popcount36_9tg7_core_225 = ~(input_a[1] & input_a[4]);
  assign popcount36_9tg7_core_227 = input_a[20] ^ input_a[19];
  assign popcount36_9tg7_core_230 = input_a[15] | input_a[31];
  assign popcount36_9tg7_core_232 = ~input_a[34];
  assign popcount36_9tg7_core_234 = input_a[20] | input_a[12];
  assign popcount36_9tg7_core_236 = ~(input_a[31] ^ input_a[15]);
  assign popcount36_9tg7_core_237 = input_a[14] ^ input_a[25];
  assign popcount36_9tg7_core_238 = ~(input_a[10] | input_a[34]);
  assign popcount36_9tg7_core_239 = input_a[35] ^ input_a[30];
  assign popcount36_9tg7_core_244 = ~(input_a[7] ^ input_a[6]);
  assign popcount36_9tg7_core_245 = ~(input_a[28] & input_a[0]);
  assign popcount36_9tg7_core_246 = input_a[10] & input_a[30];
  assign popcount36_9tg7_core_249 = ~input_a[20];
  assign popcount36_9tg7_core_251 = input_a[29] & input_a[16];
  assign popcount36_9tg7_core_256 = input_a[3] & input_a[0];
  assign popcount36_9tg7_core_258 = input_a[24] | input_a[12];
  assign popcount36_9tg7_core_259 = ~(input_a[4] & input_a[8]);
  assign popcount36_9tg7_core_261 = input_a[15] | input_a[23];
  assign popcount36_9tg7_core_262 = input_a[7] & input_a[6];
  assign popcount36_9tg7_core_263_not = ~input_a[23];
  assign popcount36_9tg7_core_264 = ~input_a[35];
  assign popcount36_9tg7_core_265 = ~(input_a[27] ^ input_a[2]);
  assign popcount36_9tg7_core_267 = ~(input_a[30] | input_a[12]);
  assign popcount36_9tg7_core_268 = input_a[31] & input_a[23];
  assign popcount36_9tg7_core_270 = ~(input_a[27] | input_a[21]);
  assign popcount36_9tg7_core_272 = ~(input_a[16] ^ input_a[11]);
  assign popcount36_9tg7_core_273 = input_a[4] & input_a[1];
  assign popcount36_9tg7_core_274 = input_a[24] & input_a[14];
  assign popcount36_9tg7_core_275 = input_a[31] & input_a[0];
  assign popcount36_9tg7_core_276 = input_a[15] | input_a[1];

  assign popcount36_9tg7_out[0] = input_a[15];
  assign popcount36_9tg7_out[1] = input_a[1];
  assign popcount36_9tg7_out[2] = input_a[24];
  assign popcount36_9tg7_out[3] = input_a[7];
  assign popcount36_9tg7_out[4] = input_a[2];
  assign popcount36_9tg7_out[5] = 1'b0;
endmodule