// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=8.31678
// WCE=35.0
// EP=0.965255%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_go6i(input [38:0] input_a, output [5:0] popcount39_go6i_out);
  wire popcount39_go6i_core_041;
  wire popcount39_go6i_core_042;
  wire popcount39_go6i_core_043;
  wire popcount39_go6i_core_044;
  wire popcount39_go6i_core_045;
  wire popcount39_go6i_core_047;
  wire popcount39_go6i_core_049_not;
  wire popcount39_go6i_core_051;
  wire popcount39_go6i_core_053;
  wire popcount39_go6i_core_056;
  wire popcount39_go6i_core_057;
  wire popcount39_go6i_core_058_not;
  wire popcount39_go6i_core_060;
  wire popcount39_go6i_core_063;
  wire popcount39_go6i_core_066;
  wire popcount39_go6i_core_067;
  wire popcount39_go6i_core_068;
  wire popcount39_go6i_core_069;
  wire popcount39_go6i_core_070;
  wire popcount39_go6i_core_071;
  wire popcount39_go6i_core_072;
  wire popcount39_go6i_core_073;
  wire popcount39_go6i_core_074;
  wire popcount39_go6i_core_076;
  wire popcount39_go6i_core_077;
  wire popcount39_go6i_core_079;
  wire popcount39_go6i_core_080;
  wire popcount39_go6i_core_083;
  wire popcount39_go6i_core_084;
  wire popcount39_go6i_core_085;
  wire popcount39_go6i_core_086;
  wire popcount39_go6i_core_087;
  wire popcount39_go6i_core_089;
  wire popcount39_go6i_core_091;
  wire popcount39_go6i_core_092;
  wire popcount39_go6i_core_093;
  wire popcount39_go6i_core_095;
  wire popcount39_go6i_core_096;
  wire popcount39_go6i_core_097;
  wire popcount39_go6i_core_098;
  wire popcount39_go6i_core_099;
  wire popcount39_go6i_core_100;
  wire popcount39_go6i_core_101;
  wire popcount39_go6i_core_103;
  wire popcount39_go6i_core_106;
  wire popcount39_go6i_core_108;
  wire popcount39_go6i_core_109;
  wire popcount39_go6i_core_110;
  wire popcount39_go6i_core_111;
  wire popcount39_go6i_core_113;
  wire popcount39_go6i_core_114;
  wire popcount39_go6i_core_115;
  wire popcount39_go6i_core_116;
  wire popcount39_go6i_core_117;
  wire popcount39_go6i_core_119;
  wire popcount39_go6i_core_120;
  wire popcount39_go6i_core_121;
  wire popcount39_go6i_core_122;
  wire popcount39_go6i_core_126;
  wire popcount39_go6i_core_127;
  wire popcount39_go6i_core_130;
  wire popcount39_go6i_core_132;
  wire popcount39_go6i_core_133;
  wire popcount39_go6i_core_134;
  wire popcount39_go6i_core_136;
  wire popcount39_go6i_core_137;
  wire popcount39_go6i_core_138;
  wire popcount39_go6i_core_139;
  wire popcount39_go6i_core_140;
  wire popcount39_go6i_core_141;
  wire popcount39_go6i_core_142;
  wire popcount39_go6i_core_143;
  wire popcount39_go6i_core_144;
  wire popcount39_go6i_core_145;
  wire popcount39_go6i_core_146;
  wire popcount39_go6i_core_147;
  wire popcount39_go6i_core_149;
  wire popcount39_go6i_core_150;
  wire popcount39_go6i_core_151;
  wire popcount39_go6i_core_152;
  wire popcount39_go6i_core_155;
  wire popcount39_go6i_core_156;
  wire popcount39_go6i_core_158;
  wire popcount39_go6i_core_159;
  wire popcount39_go6i_core_160;
  wire popcount39_go6i_core_162;
  wire popcount39_go6i_core_163_not;
  wire popcount39_go6i_core_164;
  wire popcount39_go6i_core_166;
  wire popcount39_go6i_core_167;
  wire popcount39_go6i_core_168;
  wire popcount39_go6i_core_170;
  wire popcount39_go6i_core_171;
  wire popcount39_go6i_core_172;
  wire popcount39_go6i_core_173;
  wire popcount39_go6i_core_174;
  wire popcount39_go6i_core_176;
  wire popcount39_go6i_core_177;
  wire popcount39_go6i_core_178;
  wire popcount39_go6i_core_179;
  wire popcount39_go6i_core_183;
  wire popcount39_go6i_core_186;
  wire popcount39_go6i_core_187;
  wire popcount39_go6i_core_188;
  wire popcount39_go6i_core_190;
  wire popcount39_go6i_core_191;
  wire popcount39_go6i_core_192;
  wire popcount39_go6i_core_193;
  wire popcount39_go6i_core_194;
  wire popcount39_go6i_core_198;
  wire popcount39_go6i_core_199;
  wire popcount39_go6i_core_204;
  wire popcount39_go6i_core_206;
  wire popcount39_go6i_core_207;
  wire popcount39_go6i_core_208;
  wire popcount39_go6i_core_209;
  wire popcount39_go6i_core_210;
  wire popcount39_go6i_core_211;
  wire popcount39_go6i_core_213;
  wire popcount39_go6i_core_214_not;
  wire popcount39_go6i_core_216;
  wire popcount39_go6i_core_217;
  wire popcount39_go6i_core_220;
  wire popcount39_go6i_core_221;
  wire popcount39_go6i_core_222;
  wire popcount39_go6i_core_223;
  wire popcount39_go6i_core_225;
  wire popcount39_go6i_core_226;
  wire popcount39_go6i_core_227;
  wire popcount39_go6i_core_228;
  wire popcount39_go6i_core_229;
  wire popcount39_go6i_core_231;
  wire popcount39_go6i_core_232;
  wire popcount39_go6i_core_234;
  wire popcount39_go6i_core_235;
  wire popcount39_go6i_core_237;
  wire popcount39_go6i_core_238;
  wire popcount39_go6i_core_239;
  wire popcount39_go6i_core_240;
  wire popcount39_go6i_core_241;
  wire popcount39_go6i_core_243;
  wire popcount39_go6i_core_245;
  wire popcount39_go6i_core_246;
  wire popcount39_go6i_core_248;
  wire popcount39_go6i_core_252;
  wire popcount39_go6i_core_254;
  wire popcount39_go6i_core_255;
  wire popcount39_go6i_core_256;
  wire popcount39_go6i_core_257;
  wire popcount39_go6i_core_258;
  wire popcount39_go6i_core_259;
  wire popcount39_go6i_core_260;
  wire popcount39_go6i_core_261;
  wire popcount39_go6i_core_262;
  wire popcount39_go6i_core_263;
  wire popcount39_go6i_core_266;
  wire popcount39_go6i_core_267;
  wire popcount39_go6i_core_268;
  wire popcount39_go6i_core_270;
  wire popcount39_go6i_core_271;
  wire popcount39_go6i_core_273;
  wire popcount39_go6i_core_274;
  wire popcount39_go6i_core_275;
  wire popcount39_go6i_core_276;
  wire popcount39_go6i_core_277;
  wire popcount39_go6i_core_278;
  wire popcount39_go6i_core_279;
  wire popcount39_go6i_core_280;
  wire popcount39_go6i_core_281;
  wire popcount39_go6i_core_282;
  wire popcount39_go6i_core_283;
  wire popcount39_go6i_core_284;
  wire popcount39_go6i_core_286;
  wire popcount39_go6i_core_287;
  wire popcount39_go6i_core_291;
  wire popcount39_go6i_core_292;
  wire popcount39_go6i_core_293;
  wire popcount39_go6i_core_294;
  wire popcount39_go6i_core_295;
  wire popcount39_go6i_core_297;
  wire popcount39_go6i_core_299;
  wire popcount39_go6i_core_300;
  wire popcount39_go6i_core_301;
  wire popcount39_go6i_core_302_not;
  wire popcount39_go6i_core_304_not;

  assign popcount39_go6i_core_041 = input_a[34] ^ input_a[31];
  assign popcount39_go6i_core_042 = input_a[24] & input_a[16];
  assign popcount39_go6i_core_043 = input_a[34] & input_a[25];
  assign popcount39_go6i_core_044 = ~(input_a[26] | input_a[23]);
  assign popcount39_go6i_core_045 = ~(input_a[21] | input_a[14]);
  assign popcount39_go6i_core_047 = ~(input_a[37] ^ input_a[3]);
  assign popcount39_go6i_core_049_not = ~input_a[24];
  assign popcount39_go6i_core_051 = ~input_a[4];
  assign popcount39_go6i_core_053 = ~input_a[24];
  assign popcount39_go6i_core_056 = ~(input_a[8] ^ input_a[34]);
  assign popcount39_go6i_core_057 = input_a[26] | input_a[2];
  assign popcount39_go6i_core_058_not = ~input_a[17];
  assign popcount39_go6i_core_060 = ~(input_a[10] | input_a[11]);
  assign popcount39_go6i_core_063 = input_a[26] ^ input_a[29];
  assign popcount39_go6i_core_066 = input_a[18] ^ input_a[21];
  assign popcount39_go6i_core_067 = ~input_a[28];
  assign popcount39_go6i_core_068 = ~(input_a[20] | input_a[1]);
  assign popcount39_go6i_core_069 = input_a[8] ^ input_a[22];
  assign popcount39_go6i_core_070 = ~input_a[7];
  assign popcount39_go6i_core_071 = ~input_a[17];
  assign popcount39_go6i_core_072 = ~input_a[29];
  assign popcount39_go6i_core_073 = input_a[28] ^ input_a[10];
  assign popcount39_go6i_core_074 = ~(input_a[10] | input_a[7]);
  assign popcount39_go6i_core_076 = ~(input_a[10] & input_a[0]);
  assign popcount39_go6i_core_077 = input_a[2] & input_a[24];
  assign popcount39_go6i_core_079 = ~input_a[13];
  assign popcount39_go6i_core_080 = ~(input_a[27] | input_a[11]);
  assign popcount39_go6i_core_083 = ~(input_a[7] ^ input_a[29]);
  assign popcount39_go6i_core_084 = ~input_a[18];
  assign popcount39_go6i_core_085 = input_a[34] | input_a[37];
  assign popcount39_go6i_core_086 = ~(input_a[10] & input_a[10]);
  assign popcount39_go6i_core_087 = ~(input_a[30] & input_a[35]);
  assign popcount39_go6i_core_089 = input_a[22] ^ input_a[27];
  assign popcount39_go6i_core_091 = input_a[1] | input_a[28];
  assign popcount39_go6i_core_092 = input_a[3] & input_a[5];
  assign popcount39_go6i_core_093 = input_a[5] ^ input_a[27];
  assign popcount39_go6i_core_095 = input_a[37] | input_a[4];
  assign popcount39_go6i_core_096 = ~(input_a[14] & input_a[29]);
  assign popcount39_go6i_core_097 = ~(input_a[5] ^ input_a[32]);
  assign popcount39_go6i_core_098 = input_a[17] | input_a[21];
  assign popcount39_go6i_core_099 = ~(input_a[7] | input_a[15]);
  assign popcount39_go6i_core_100 = input_a[20] | input_a[33];
  assign popcount39_go6i_core_101 = input_a[34] | input_a[12];
  assign popcount39_go6i_core_103 = ~(input_a[2] & input_a[36]);
  assign popcount39_go6i_core_106 = input_a[18] & input_a[21];
  assign popcount39_go6i_core_108 = input_a[18] | input_a[8];
  assign popcount39_go6i_core_109 = ~(input_a[6] ^ input_a[27]);
  assign popcount39_go6i_core_110 = ~input_a[8];
  assign popcount39_go6i_core_111 = input_a[17] ^ input_a[37];
  assign popcount39_go6i_core_113 = input_a[1] ^ input_a[14];
  assign popcount39_go6i_core_114 = input_a[6] ^ input_a[20];
  assign popcount39_go6i_core_115 = input_a[5] | input_a[1];
  assign popcount39_go6i_core_116 = ~(input_a[1] ^ input_a[21]);
  assign popcount39_go6i_core_117 = input_a[14] ^ input_a[2];
  assign popcount39_go6i_core_119 = ~(input_a[35] & input_a[9]);
  assign popcount39_go6i_core_120 = ~(input_a[16] & input_a[34]);
  assign popcount39_go6i_core_121 = input_a[37] | input_a[24];
  assign popcount39_go6i_core_122 = input_a[7] | input_a[12];
  assign popcount39_go6i_core_126 = ~(input_a[13] ^ input_a[27]);
  assign popcount39_go6i_core_127 = ~input_a[6];
  assign popcount39_go6i_core_130 = ~(input_a[5] ^ input_a[34]);
  assign popcount39_go6i_core_132 = ~(input_a[26] | input_a[25]);
  assign popcount39_go6i_core_133 = input_a[1] | input_a[16];
  assign popcount39_go6i_core_134 = ~(input_a[8] ^ input_a[34]);
  assign popcount39_go6i_core_136 = input_a[9] | input_a[36];
  assign popcount39_go6i_core_137 = ~(input_a[17] | input_a[8]);
  assign popcount39_go6i_core_138 = input_a[24] ^ input_a[26];
  assign popcount39_go6i_core_139 = input_a[20] | input_a[36];
  assign popcount39_go6i_core_140 = input_a[2] & input_a[33];
  assign popcount39_go6i_core_141 = ~(input_a[26] ^ input_a[26]);
  assign popcount39_go6i_core_142 = ~(input_a[4] & input_a[15]);
  assign popcount39_go6i_core_143 = input_a[8] & input_a[6];
  assign popcount39_go6i_core_144 = input_a[31] | input_a[19];
  assign popcount39_go6i_core_145 = ~(input_a[18] ^ input_a[6]);
  assign popcount39_go6i_core_146 = input_a[21] | input_a[9];
  assign popcount39_go6i_core_147 = ~(input_a[34] | input_a[32]);
  assign popcount39_go6i_core_149 = ~(input_a[17] | input_a[36]);
  assign popcount39_go6i_core_150 = input_a[33] & input_a[33];
  assign popcount39_go6i_core_151 = ~(input_a[8] ^ input_a[25]);
  assign popcount39_go6i_core_152 = input_a[37] ^ input_a[21];
  assign popcount39_go6i_core_155 = input_a[5] ^ input_a[15];
  assign popcount39_go6i_core_156 = input_a[11] ^ input_a[33];
  assign popcount39_go6i_core_158 = ~(input_a[9] | input_a[22]);
  assign popcount39_go6i_core_159 = input_a[11] ^ input_a[24];
  assign popcount39_go6i_core_160 = input_a[10] ^ input_a[3];
  assign popcount39_go6i_core_162 = ~(input_a[36] | input_a[31]);
  assign popcount39_go6i_core_163_not = ~input_a[0];
  assign popcount39_go6i_core_164 = ~(input_a[5] | input_a[13]);
  assign popcount39_go6i_core_166 = input_a[21] | input_a[15];
  assign popcount39_go6i_core_167 = input_a[21] ^ input_a[21];
  assign popcount39_go6i_core_168 = input_a[36] ^ input_a[19];
  assign popcount39_go6i_core_170 = input_a[7] ^ input_a[36];
  assign popcount39_go6i_core_171 = ~(input_a[13] ^ input_a[8]);
  assign popcount39_go6i_core_172 = input_a[19] & input_a[26];
  assign popcount39_go6i_core_173 = input_a[19] & input_a[28];
  assign popcount39_go6i_core_174 = input_a[13] & input_a[38];
  assign popcount39_go6i_core_176 = input_a[32] ^ input_a[12];
  assign popcount39_go6i_core_177 = input_a[17] ^ input_a[3];
  assign popcount39_go6i_core_178 = input_a[32] & input_a[28];
  assign popcount39_go6i_core_179 = ~(input_a[15] & input_a[9]);
  assign popcount39_go6i_core_183 = ~input_a[5];
  assign popcount39_go6i_core_186 = ~(input_a[13] ^ input_a[13]);
  assign popcount39_go6i_core_187 = ~(input_a[18] | input_a[34]);
  assign popcount39_go6i_core_188 = ~(input_a[20] ^ input_a[3]);
  assign popcount39_go6i_core_190 = input_a[1] & input_a[23];
  assign popcount39_go6i_core_191 = input_a[15] & input_a[26];
  assign popcount39_go6i_core_192 = input_a[24] & input_a[34];
  assign popcount39_go6i_core_193 = ~(input_a[17] & input_a[28]);
  assign popcount39_go6i_core_194 = ~(input_a[12] ^ input_a[29]);
  assign popcount39_go6i_core_198 = input_a[11] | input_a[9];
  assign popcount39_go6i_core_199 = ~(input_a[14] | input_a[6]);
  assign popcount39_go6i_core_204 = input_a[24] ^ input_a[30];
  assign popcount39_go6i_core_206 = input_a[30] | input_a[5];
  assign popcount39_go6i_core_207 = ~(input_a[13] & input_a[9]);
  assign popcount39_go6i_core_208 = ~(input_a[28] | input_a[16]);
  assign popcount39_go6i_core_209 = ~input_a[27];
  assign popcount39_go6i_core_210 = input_a[31] | input_a[23];
  assign popcount39_go6i_core_211 = ~(input_a[17] ^ input_a[13]);
  assign popcount39_go6i_core_213 = input_a[16] ^ input_a[11];
  assign popcount39_go6i_core_214_not = ~input_a[25];
  assign popcount39_go6i_core_216 = input_a[28] | input_a[9];
  assign popcount39_go6i_core_217 = ~(input_a[21] & input_a[34]);
  assign popcount39_go6i_core_220 = input_a[7] | input_a[32];
  assign popcount39_go6i_core_221 = ~(input_a[19] & input_a[24]);
  assign popcount39_go6i_core_222 = input_a[25] & input_a[36];
  assign popcount39_go6i_core_223 = input_a[8] & input_a[13];
  assign popcount39_go6i_core_225 = ~(input_a[3] ^ input_a[7]);
  assign popcount39_go6i_core_226 = ~(input_a[23] ^ input_a[35]);
  assign popcount39_go6i_core_227 = input_a[3] ^ input_a[10];
  assign popcount39_go6i_core_228 = ~(input_a[13] ^ input_a[13]);
  assign popcount39_go6i_core_229 = input_a[8] & input_a[20];
  assign popcount39_go6i_core_231 = input_a[37] ^ input_a[26];
  assign popcount39_go6i_core_232 = ~input_a[12];
  assign popcount39_go6i_core_234 = ~(input_a[1] | input_a[17]);
  assign popcount39_go6i_core_235 = ~(input_a[21] ^ input_a[29]);
  assign popcount39_go6i_core_237 = ~(input_a[36] | input_a[21]);
  assign popcount39_go6i_core_238 = ~(input_a[13] | input_a[12]);
  assign popcount39_go6i_core_239 = ~input_a[20];
  assign popcount39_go6i_core_240 = input_a[20] ^ input_a[7];
  assign popcount39_go6i_core_241 = ~(input_a[28] & input_a[35]);
  assign popcount39_go6i_core_243 = ~input_a[3];
  assign popcount39_go6i_core_245 = ~(input_a[10] ^ input_a[14]);
  assign popcount39_go6i_core_246 = input_a[31] & input_a[28];
  assign popcount39_go6i_core_248 = ~input_a[12];
  assign popcount39_go6i_core_252 = input_a[23] & input_a[7];
  assign popcount39_go6i_core_254 = ~(input_a[25] ^ input_a[10]);
  assign popcount39_go6i_core_255 = input_a[2] | input_a[23];
  assign popcount39_go6i_core_256 = input_a[21] & input_a[36];
  assign popcount39_go6i_core_257 = input_a[26] & input_a[26];
  assign popcount39_go6i_core_258 = input_a[4] | input_a[10];
  assign popcount39_go6i_core_259 = input_a[16] | input_a[26];
  assign popcount39_go6i_core_260 = input_a[34] ^ input_a[0];
  assign popcount39_go6i_core_261 = ~(input_a[2] ^ input_a[24]);
  assign popcount39_go6i_core_262 = input_a[32] ^ input_a[31];
  assign popcount39_go6i_core_263 = input_a[2] ^ input_a[28];
  assign popcount39_go6i_core_266 = input_a[13] ^ input_a[15];
  assign popcount39_go6i_core_267 = ~(input_a[30] ^ input_a[12]);
  assign popcount39_go6i_core_268 = ~(input_a[33] & input_a[13]);
  assign popcount39_go6i_core_270 = ~(input_a[21] | input_a[24]);
  assign popcount39_go6i_core_271 = ~(input_a[7] ^ input_a[12]);
  assign popcount39_go6i_core_273 = ~input_a[23];
  assign popcount39_go6i_core_274 = ~(input_a[11] ^ input_a[34]);
  assign popcount39_go6i_core_275 = ~(input_a[36] & input_a[38]);
  assign popcount39_go6i_core_276 = input_a[32] ^ input_a[26];
  assign popcount39_go6i_core_277 = input_a[5] | input_a[33];
  assign popcount39_go6i_core_278 = ~(input_a[0] & input_a[24]);
  assign popcount39_go6i_core_279 = ~(input_a[24] & input_a[9]);
  assign popcount39_go6i_core_280 = ~(input_a[17] | input_a[4]);
  assign popcount39_go6i_core_281 = input_a[3] & input_a[35];
  assign popcount39_go6i_core_282 = input_a[20] | input_a[31];
  assign popcount39_go6i_core_283 = input_a[2] ^ input_a[26];
  assign popcount39_go6i_core_284 = input_a[21] ^ input_a[3];
  assign popcount39_go6i_core_286 = input_a[9] & input_a[10];
  assign popcount39_go6i_core_287 = ~input_a[11];
  assign popcount39_go6i_core_291 = ~(input_a[12] & input_a[14]);
  assign popcount39_go6i_core_292 = ~(input_a[25] ^ input_a[21]);
  assign popcount39_go6i_core_293 = ~input_a[31];
  assign popcount39_go6i_core_294 = ~(input_a[22] & input_a[30]);
  assign popcount39_go6i_core_295 = ~(input_a[14] | input_a[0]);
  assign popcount39_go6i_core_297 = input_a[17] | input_a[5];
  assign popcount39_go6i_core_299 = input_a[13] | input_a[30];
  assign popcount39_go6i_core_300 = input_a[1] | input_a[27];
  assign popcount39_go6i_core_301 = input_a[36] & input_a[36];
  assign popcount39_go6i_core_302_not = ~input_a[19];
  assign popcount39_go6i_core_304_not = ~input_a[22];

  assign popcount39_go6i_out[0] = 1'b0;
  assign popcount39_go6i_out[1] = input_a[21];
  assign popcount39_go6i_out[2] = input_a[32];
  assign popcount39_go6i_out[3] = input_a[30];
  assign popcount39_go6i_out[4] = input_a[8];
  assign popcount39_go6i_out[5] = 1'b0;
endmodule