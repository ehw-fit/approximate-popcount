// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.96135
// WCE=16.0
// EP=0.927611%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount21_x30l(input [20:0] input_a, output [4:0] popcount21_x30l_out);
  wire popcount21_x30l_core_023;
  wire popcount21_x30l_core_024;
  wire popcount21_x30l_core_027;
  wire popcount21_x30l_core_028;
  wire popcount21_x30l_core_030;
  wire popcount21_x30l_core_031;
  wire popcount21_x30l_core_033;
  wire popcount21_x30l_core_034;
  wire popcount21_x30l_core_036;
  wire popcount21_x30l_core_039;
  wire popcount21_x30l_core_043;
  wire popcount21_x30l_core_046;
  wire popcount21_x30l_core_047;
  wire popcount21_x30l_core_048;
  wire popcount21_x30l_core_049;
  wire popcount21_x30l_core_050_not;
  wire popcount21_x30l_core_052;
  wire popcount21_x30l_core_053;
  wire popcount21_x30l_core_054;
  wire popcount21_x30l_core_055;
  wire popcount21_x30l_core_056;
  wire popcount21_x30l_core_057;
  wire popcount21_x30l_core_058_not;
  wire popcount21_x30l_core_060_not;
  wire popcount21_x30l_core_062;
  wire popcount21_x30l_core_063;
  wire popcount21_x30l_core_064;
  wire popcount21_x30l_core_065;
  wire popcount21_x30l_core_067;
  wire popcount21_x30l_core_068;
  wire popcount21_x30l_core_070;
  wire popcount21_x30l_core_074;
  wire popcount21_x30l_core_075;
  wire popcount21_x30l_core_076;
  wire popcount21_x30l_core_077;
  wire popcount21_x30l_core_078;
  wire popcount21_x30l_core_079;
  wire popcount21_x30l_core_083;
  wire popcount21_x30l_core_085;
  wire popcount21_x30l_core_086;
  wire popcount21_x30l_core_088;
  wire popcount21_x30l_core_089;
  wire popcount21_x30l_core_095;
  wire popcount21_x30l_core_102;
  wire popcount21_x30l_core_105;
  wire popcount21_x30l_core_106;
  wire popcount21_x30l_core_107;
  wire popcount21_x30l_core_108;
  wire popcount21_x30l_core_109;
  wire popcount21_x30l_core_111;
  wire popcount21_x30l_core_112;
  wire popcount21_x30l_core_114;
  wire popcount21_x30l_core_115;
  wire popcount21_x30l_core_116;
  wire popcount21_x30l_core_117;
  wire popcount21_x30l_core_120;
  wire popcount21_x30l_core_121;
  wire popcount21_x30l_core_122;
  wire popcount21_x30l_core_123;
  wire popcount21_x30l_core_125;
  wire popcount21_x30l_core_126;
  wire popcount21_x30l_core_127;
  wire popcount21_x30l_core_128;
  wire popcount21_x30l_core_130;
  wire popcount21_x30l_core_131;
  wire popcount21_x30l_core_132;
  wire popcount21_x30l_core_133;
  wire popcount21_x30l_core_136;
  wire popcount21_x30l_core_139;
  wire popcount21_x30l_core_140_not;
  wire popcount21_x30l_core_141;
  wire popcount21_x30l_core_142_not;
  wire popcount21_x30l_core_144;
  wire popcount21_x30l_core_145;
  wire popcount21_x30l_core_146;
  wire popcount21_x30l_core_147;
  wire popcount21_x30l_core_148;
  wire popcount21_x30l_core_151;
  wire popcount21_x30l_core_152;
  wire popcount21_x30l_core_153;

  assign popcount21_x30l_core_023 = ~(input_a[3] | input_a[7]);
  assign popcount21_x30l_core_024 = ~input_a[12];
  assign popcount21_x30l_core_027 = input_a[4] ^ input_a[9];
  assign popcount21_x30l_core_028 = input_a[15] | input_a[10];
  assign popcount21_x30l_core_030 = input_a[10] ^ input_a[18];
  assign popcount21_x30l_core_031 = input_a[20] | input_a[3];
  assign popcount21_x30l_core_033 = input_a[2] | input_a[12];
  assign popcount21_x30l_core_034 = ~input_a[14];
  assign popcount21_x30l_core_036 = ~input_a[20];
  assign popcount21_x30l_core_039 = input_a[16] ^ input_a[0];
  assign popcount21_x30l_core_043 = input_a[18] & input_a[20];
  assign popcount21_x30l_core_046 = ~(input_a[14] | input_a[7]);
  assign popcount21_x30l_core_047 = ~(input_a[12] | input_a[9]);
  assign popcount21_x30l_core_048 = input_a[17] ^ input_a[2];
  assign popcount21_x30l_core_049 = ~input_a[3];
  assign popcount21_x30l_core_050_not = ~input_a[9];
  assign popcount21_x30l_core_052 = ~input_a[17];
  assign popcount21_x30l_core_053 = ~(input_a[10] ^ input_a[12]);
  assign popcount21_x30l_core_054 = ~input_a[18];
  assign popcount21_x30l_core_055 = ~(input_a[20] & input_a[2]);
  assign popcount21_x30l_core_056 = input_a[4] | input_a[13];
  assign popcount21_x30l_core_057 = input_a[13] | input_a[5];
  assign popcount21_x30l_core_058_not = ~input_a[5];
  assign popcount21_x30l_core_060_not = ~input_a[17];
  assign popcount21_x30l_core_062 = ~input_a[11];
  assign popcount21_x30l_core_063 = ~(input_a[11] & input_a[1]);
  assign popcount21_x30l_core_064 = input_a[14] | input_a[7];
  assign popcount21_x30l_core_065 = ~input_a[16];
  assign popcount21_x30l_core_067 = input_a[7] | input_a[2];
  assign popcount21_x30l_core_068 = input_a[19] ^ input_a[19];
  assign popcount21_x30l_core_070 = ~(input_a[3] | input_a[1]);
  assign popcount21_x30l_core_074 = input_a[18] | input_a[16];
  assign popcount21_x30l_core_075 = ~input_a[13];
  assign popcount21_x30l_core_076 = input_a[6] ^ input_a[17];
  assign popcount21_x30l_core_077 = input_a[10] ^ input_a[4];
  assign popcount21_x30l_core_078 = ~(input_a[8] & input_a[0]);
  assign popcount21_x30l_core_079 = input_a[10] | input_a[14];
  assign popcount21_x30l_core_083 = ~input_a[15];
  assign popcount21_x30l_core_085 = input_a[10] & input_a[20];
  assign popcount21_x30l_core_086 = input_a[9] ^ input_a[17];
  assign popcount21_x30l_core_088 = input_a[13] ^ input_a[17];
  assign popcount21_x30l_core_089 = ~input_a[19];
  assign popcount21_x30l_core_095 = input_a[5] | input_a[9];
  assign popcount21_x30l_core_102 = input_a[20] & input_a[15];
  assign popcount21_x30l_core_105 = ~(input_a[12] | input_a[19]);
  assign popcount21_x30l_core_106 = ~(input_a[20] ^ input_a[20]);
  assign popcount21_x30l_core_107 = ~(input_a[2] ^ input_a[0]);
  assign popcount21_x30l_core_108 = input_a[5] & input_a[7];
  assign popcount21_x30l_core_109 = input_a[6] | input_a[19];
  assign popcount21_x30l_core_111 = ~(input_a[9] & input_a[7]);
  assign popcount21_x30l_core_112 = ~(input_a[1] & input_a[11]);
  assign popcount21_x30l_core_114 = input_a[4] & input_a[15];
  assign popcount21_x30l_core_115 = ~input_a[0];
  assign popcount21_x30l_core_116 = ~input_a[14];
  assign popcount21_x30l_core_117 = input_a[4] ^ input_a[4];
  assign popcount21_x30l_core_120 = ~(input_a[3] ^ input_a[10]);
  assign popcount21_x30l_core_121 = ~(input_a[7] | input_a[3]);
  assign popcount21_x30l_core_122 = ~(input_a[0] ^ input_a[19]);
  assign popcount21_x30l_core_123 = ~(input_a[18] ^ input_a[12]);
  assign popcount21_x30l_core_125 = ~(input_a[14] | input_a[8]);
  assign popcount21_x30l_core_126 = input_a[14] | input_a[10];
  assign popcount21_x30l_core_127 = ~(input_a[12] | input_a[2]);
  assign popcount21_x30l_core_128 = ~input_a[7];
  assign popcount21_x30l_core_130 = ~(input_a[4] & input_a[1]);
  assign popcount21_x30l_core_131 = ~(input_a[4] ^ input_a[15]);
  assign popcount21_x30l_core_132 = input_a[7] ^ input_a[3];
  assign popcount21_x30l_core_133 = ~(input_a[2] | input_a[13]);
  assign popcount21_x30l_core_136 = ~(input_a[20] & input_a[11]);
  assign popcount21_x30l_core_139 = input_a[0] & input_a[15];
  assign popcount21_x30l_core_140_not = ~input_a[17];
  assign popcount21_x30l_core_141 = ~(input_a[7] & input_a[17]);
  assign popcount21_x30l_core_142_not = ~input_a[10];
  assign popcount21_x30l_core_144 = ~(input_a[2] | input_a[5]);
  assign popcount21_x30l_core_145 = input_a[9] & input_a[10];
  assign popcount21_x30l_core_146 = input_a[7] | input_a[1];
  assign popcount21_x30l_core_147 = input_a[6] & input_a[4];
  assign popcount21_x30l_core_148 = ~(input_a[19] | input_a[0]);
  assign popcount21_x30l_core_151 = input_a[1] ^ input_a[5];
  assign popcount21_x30l_core_152 = input_a[8] & input_a[18];
  assign popcount21_x30l_core_153 = input_a[1] | input_a[18];

  assign popcount21_x30l_out[0] = input_a[7];
  assign popcount21_x30l_out[1] = 1'b1;
  assign popcount21_x30l_out[2] = input_a[14];
  assign popcount21_x30l_out[3] = input_a[13];
  assign popcount21_x30l_out[4] = 1'b0;
endmodule