// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.70128
// WCE=17.0
// EP=0.937145%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount27_j1oh(input [26:0] input_a, output [4:0] popcount27_j1oh_out);
  wire popcount27_j1oh_core_029;
  wire popcount27_j1oh_core_033;
  wire popcount27_j1oh_core_034;
  wire popcount27_j1oh_core_036;
  wire popcount27_j1oh_core_038_not;
  wire popcount27_j1oh_core_039;
  wire popcount27_j1oh_core_040;
  wire popcount27_j1oh_core_044;
  wire popcount27_j1oh_core_046;
  wire popcount27_j1oh_core_047;
  wire popcount27_j1oh_core_049;
  wire popcount27_j1oh_core_051;
  wire popcount27_j1oh_core_052;
  wire popcount27_j1oh_core_055;
  wire popcount27_j1oh_core_057;
  wire popcount27_j1oh_core_058;
  wire popcount27_j1oh_core_059;
  wire popcount27_j1oh_core_060;
  wire popcount27_j1oh_core_061;
  wire popcount27_j1oh_core_063;
  wire popcount27_j1oh_core_065;
  wire popcount27_j1oh_core_068;
  wire popcount27_j1oh_core_070;
  wire popcount27_j1oh_core_072;
  wire popcount27_j1oh_core_073;
  wire popcount27_j1oh_core_074;
  wire popcount27_j1oh_core_075;
  wire popcount27_j1oh_core_076;
  wire popcount27_j1oh_core_077;
  wire popcount27_j1oh_core_078;
  wire popcount27_j1oh_core_080;
  wire popcount27_j1oh_core_081;
  wire popcount27_j1oh_core_083;
  wire popcount27_j1oh_core_086;
  wire popcount27_j1oh_core_087;
  wire popcount27_j1oh_core_090;
  wire popcount27_j1oh_core_093;
  wire popcount27_j1oh_core_094;
  wire popcount27_j1oh_core_095;
  wire popcount27_j1oh_core_096;
  wire popcount27_j1oh_core_098;
  wire popcount27_j1oh_core_100;
  wire popcount27_j1oh_core_101;
  wire popcount27_j1oh_core_103;
  wire popcount27_j1oh_core_104;
  wire popcount27_j1oh_core_106;
  wire popcount27_j1oh_core_107;
  wire popcount27_j1oh_core_108;
  wire popcount27_j1oh_core_109;
  wire popcount27_j1oh_core_111;
  wire popcount27_j1oh_core_112;
  wire popcount27_j1oh_core_113;
  wire popcount27_j1oh_core_115;
  wire popcount27_j1oh_core_118;
  wire popcount27_j1oh_core_119;
  wire popcount27_j1oh_core_121;
  wire popcount27_j1oh_core_122;
  wire popcount27_j1oh_core_123;
  wire popcount27_j1oh_core_124;
  wire popcount27_j1oh_core_125;
  wire popcount27_j1oh_core_126;
  wire popcount27_j1oh_core_127;
  wire popcount27_j1oh_core_128;
  wire popcount27_j1oh_core_129;
  wire popcount27_j1oh_core_132;
  wire popcount27_j1oh_core_133;
  wire popcount27_j1oh_core_134_not;
  wire popcount27_j1oh_core_136;
  wire popcount27_j1oh_core_138;
  wire popcount27_j1oh_core_139;
  wire popcount27_j1oh_core_140;
  wire popcount27_j1oh_core_141;
  wire popcount27_j1oh_core_142;
  wire popcount27_j1oh_core_143;
  wire popcount27_j1oh_core_144_not;
  wire popcount27_j1oh_core_145;
  wire popcount27_j1oh_core_146;
  wire popcount27_j1oh_core_147;
  wire popcount27_j1oh_core_148;
  wire popcount27_j1oh_core_151;
  wire popcount27_j1oh_core_152;
  wire popcount27_j1oh_core_155;
  wire popcount27_j1oh_core_156;
  wire popcount27_j1oh_core_157;
  wire popcount27_j1oh_core_158;
  wire popcount27_j1oh_core_160;
  wire popcount27_j1oh_core_162;
  wire popcount27_j1oh_core_163;
  wire popcount27_j1oh_core_164_not;
  wire popcount27_j1oh_core_165;
  wire popcount27_j1oh_core_166;
  wire popcount27_j1oh_core_168;
  wire popcount27_j1oh_core_169;
  wire popcount27_j1oh_core_170;
  wire popcount27_j1oh_core_172;
  wire popcount27_j1oh_core_173;
  wire popcount27_j1oh_core_174;
  wire popcount27_j1oh_core_178;
  wire popcount27_j1oh_core_179;
  wire popcount27_j1oh_core_180;
  wire popcount27_j1oh_core_181;
  wire popcount27_j1oh_core_182;
  wire popcount27_j1oh_core_184;
  wire popcount27_j1oh_core_187;
  wire popcount27_j1oh_core_190;
  wire popcount27_j1oh_core_191;
  wire popcount27_j1oh_core_193;
  wire popcount27_j1oh_core_194;

  assign popcount27_j1oh_core_029 = ~input_a[26];
  assign popcount27_j1oh_core_033 = input_a[4] & input_a[8];
  assign popcount27_j1oh_core_034 = input_a[17] ^ input_a[25];
  assign popcount27_j1oh_core_036 = input_a[5] ^ input_a[18];
  assign popcount27_j1oh_core_038_not = ~input_a[7];
  assign popcount27_j1oh_core_039 = ~input_a[14];
  assign popcount27_j1oh_core_040 = ~(input_a[4] ^ input_a[3]);
  assign popcount27_j1oh_core_044 = ~(input_a[21] | input_a[1]);
  assign popcount27_j1oh_core_046 = ~(input_a[24] | input_a[24]);
  assign popcount27_j1oh_core_047 = input_a[2] | input_a[9];
  assign popcount27_j1oh_core_049 = ~input_a[6];
  assign popcount27_j1oh_core_051 = ~input_a[17];
  assign popcount27_j1oh_core_052 = ~(input_a[1] | input_a[26]);
  assign popcount27_j1oh_core_055 = ~(input_a[19] & input_a[9]);
  assign popcount27_j1oh_core_057 = ~(input_a[3] & input_a[9]);
  assign popcount27_j1oh_core_058 = input_a[24] | input_a[19];
  assign popcount27_j1oh_core_059 = ~input_a[25];
  assign popcount27_j1oh_core_060 = ~(input_a[10] & input_a[22]);
  assign popcount27_j1oh_core_061 = ~(input_a[1] | input_a[10]);
  assign popcount27_j1oh_core_063 = input_a[15] & input_a[24];
  assign popcount27_j1oh_core_065 = ~(input_a[9] | input_a[16]);
  assign popcount27_j1oh_core_068 = input_a[8] ^ input_a[26];
  assign popcount27_j1oh_core_070 = ~(input_a[21] | input_a[23]);
  assign popcount27_j1oh_core_072 = ~(input_a[7] | input_a[2]);
  assign popcount27_j1oh_core_073 = input_a[10] & input_a[25];
  assign popcount27_j1oh_core_074 = ~(input_a[9] ^ input_a[21]);
  assign popcount27_j1oh_core_075 = input_a[2] & input_a[7];
  assign popcount27_j1oh_core_076 = ~(input_a[23] | input_a[17]);
  assign popcount27_j1oh_core_077 = ~(input_a[19] ^ input_a[9]);
  assign popcount27_j1oh_core_078 = ~(input_a[9] ^ input_a[1]);
  assign popcount27_j1oh_core_080 = ~(input_a[7] & input_a[9]);
  assign popcount27_j1oh_core_081 = ~(input_a[26] | input_a[0]);
  assign popcount27_j1oh_core_083 = input_a[24] ^ input_a[3];
  assign popcount27_j1oh_core_086 = ~(input_a[14] & input_a[18]);
  assign popcount27_j1oh_core_087 = ~(input_a[6] ^ input_a[3]);
  assign popcount27_j1oh_core_090 = input_a[11] ^ input_a[3];
  assign popcount27_j1oh_core_093 = ~input_a[11];
  assign popcount27_j1oh_core_094 = ~(input_a[16] | input_a[11]);
  assign popcount27_j1oh_core_095 = ~input_a[11];
  assign popcount27_j1oh_core_096 = input_a[14] ^ input_a[13];
  assign popcount27_j1oh_core_098 = ~input_a[15];
  assign popcount27_j1oh_core_100 = ~(input_a[7] | input_a[26]);
  assign popcount27_j1oh_core_101 = ~(input_a[16] & input_a[14]);
  assign popcount27_j1oh_core_103 = ~(input_a[11] & input_a[25]);
  assign popcount27_j1oh_core_104 = ~(input_a[22] ^ input_a[17]);
  assign popcount27_j1oh_core_106 = input_a[7] & input_a[16];
  assign popcount27_j1oh_core_107 = ~(input_a[15] & input_a[26]);
  assign popcount27_j1oh_core_108 = ~(input_a[2] | input_a[26]);
  assign popcount27_j1oh_core_109 = ~(input_a[3] & input_a[19]);
  assign popcount27_j1oh_core_111 = input_a[26] | input_a[2];
  assign popcount27_j1oh_core_112 = ~(input_a[10] & input_a[12]);
  assign popcount27_j1oh_core_113 = ~(input_a[21] & input_a[3]);
  assign popcount27_j1oh_core_115 = ~(input_a[1] ^ input_a[14]);
  assign popcount27_j1oh_core_118 = input_a[9] & input_a[26];
  assign popcount27_j1oh_core_119 = ~input_a[3];
  assign popcount27_j1oh_core_121 = ~(input_a[24] & input_a[17]);
  assign popcount27_j1oh_core_122 = ~input_a[19];
  assign popcount27_j1oh_core_123 = input_a[25] | input_a[16];
  assign popcount27_j1oh_core_124 = input_a[22] | input_a[26];
  assign popcount27_j1oh_core_125 = input_a[26] ^ input_a[5];
  assign popcount27_j1oh_core_126 = input_a[14] | input_a[20];
  assign popcount27_j1oh_core_127 = input_a[6] & input_a[1];
  assign popcount27_j1oh_core_128 = ~(input_a[2] | input_a[3]);
  assign popcount27_j1oh_core_129 = ~input_a[22];
  assign popcount27_j1oh_core_132 = input_a[3] & input_a[19];
  assign popcount27_j1oh_core_133 = ~(input_a[14] | input_a[18]);
  assign popcount27_j1oh_core_134_not = ~input_a[22];
  assign popcount27_j1oh_core_136 = ~(input_a[19] & input_a[21]);
  assign popcount27_j1oh_core_138 = input_a[13] | input_a[21];
  assign popcount27_j1oh_core_139 = ~(input_a[8] | input_a[12]);
  assign popcount27_j1oh_core_140 = input_a[8] ^ input_a[18];
  assign popcount27_j1oh_core_141 = input_a[23] & input_a[3];
  assign popcount27_j1oh_core_142 = input_a[8] ^ input_a[5];
  assign popcount27_j1oh_core_143 = input_a[15] ^ input_a[12];
  assign popcount27_j1oh_core_144_not = ~input_a[6];
  assign popcount27_j1oh_core_145 = ~input_a[13];
  assign popcount27_j1oh_core_146 = input_a[23] & input_a[19];
  assign popcount27_j1oh_core_147 = ~input_a[18];
  assign popcount27_j1oh_core_148 = input_a[22] | input_a[11];
  assign popcount27_j1oh_core_151 = ~input_a[17];
  assign popcount27_j1oh_core_152 = input_a[15] | input_a[12];
  assign popcount27_j1oh_core_155 = input_a[25] | input_a[13];
  assign popcount27_j1oh_core_156 = ~(input_a[15] | input_a[20]);
  assign popcount27_j1oh_core_157 = ~(input_a[1] | input_a[25]);
  assign popcount27_j1oh_core_158 = input_a[7] & input_a[10];
  assign popcount27_j1oh_core_160 = input_a[12] & input_a[24];
  assign popcount27_j1oh_core_162 = input_a[19] & input_a[26];
  assign popcount27_j1oh_core_163 = input_a[23] | input_a[3];
  assign popcount27_j1oh_core_164_not = ~input_a[22];
  assign popcount27_j1oh_core_165 = input_a[10] ^ input_a[15];
  assign popcount27_j1oh_core_166 = input_a[13] | input_a[11];
  assign popcount27_j1oh_core_168 = input_a[16] ^ input_a[22];
  assign popcount27_j1oh_core_169 = ~(input_a[25] ^ input_a[15]);
  assign popcount27_j1oh_core_170 = ~(input_a[25] ^ input_a[22]);
  assign popcount27_j1oh_core_172 = ~(input_a[13] ^ input_a[23]);
  assign popcount27_j1oh_core_173 = ~(input_a[14] | input_a[18]);
  assign popcount27_j1oh_core_174 = ~(input_a[26] & input_a[15]);
  assign popcount27_j1oh_core_178 = ~input_a[17];
  assign popcount27_j1oh_core_179 = input_a[17] & input_a[6];
  assign popcount27_j1oh_core_180 = ~input_a[2];
  assign popcount27_j1oh_core_181 = ~(input_a[21] | input_a[13]);
  assign popcount27_j1oh_core_182 = ~(input_a[25] & input_a[1]);
  assign popcount27_j1oh_core_184 = input_a[9] ^ input_a[3];
  assign popcount27_j1oh_core_187 = input_a[10] ^ input_a[4];
  assign popcount27_j1oh_core_190 = input_a[6] & input_a[12];
  assign popcount27_j1oh_core_191 = input_a[18] & input_a[14];
  assign popcount27_j1oh_core_193 = ~(input_a[0] & input_a[26]);
  assign popcount27_j1oh_core_194 = input_a[21] | input_a[3];

  assign popcount27_j1oh_out[0] = 1'b1;
  assign popcount27_j1oh_out[1] = input_a[25];
  assign popcount27_j1oh_out[2] = 1'b0;
  assign popcount27_j1oh_out[3] = 1'b1;
  assign popcount27_j1oh_out[4] = 1'b0;
endmodule