// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.39291
// WCE=14.0
// EP=0.870702%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount25_1aj0(input [24:0] input_a, output [4:0] popcount25_1aj0_out);
  wire popcount25_1aj0_core_027;
  wire popcount25_1aj0_core_030;
  wire popcount25_1aj0_core_032;
  wire popcount25_1aj0_core_035;
  wire popcount25_1aj0_core_037;
  wire popcount25_1aj0_core_038;
  wire popcount25_1aj0_core_040;
  wire popcount25_1aj0_core_041;
  wire popcount25_1aj0_core_044;
  wire popcount25_1aj0_core_046;
  wire popcount25_1aj0_core_047;
  wire popcount25_1aj0_core_048;
  wire popcount25_1aj0_core_049;
  wire popcount25_1aj0_core_051;
  wire popcount25_1aj0_core_052;
  wire popcount25_1aj0_core_055;
  wire popcount25_1aj0_core_056_not;
  wire popcount25_1aj0_core_058;
  wire popcount25_1aj0_core_059;
  wire popcount25_1aj0_core_061;
  wire popcount25_1aj0_core_062;
  wire popcount25_1aj0_core_063_not;
  wire popcount25_1aj0_core_064;
  wire popcount25_1aj0_core_066;
  wire popcount25_1aj0_core_067;
  wire popcount25_1aj0_core_070;
  wire popcount25_1aj0_core_072;
  wire popcount25_1aj0_core_073;
  wire popcount25_1aj0_core_074;
  wire popcount25_1aj0_core_075;
  wire popcount25_1aj0_core_076;
  wire popcount25_1aj0_core_077;
  wire popcount25_1aj0_core_080_not;
  wire popcount25_1aj0_core_081;
  wire popcount25_1aj0_core_082;
  wire popcount25_1aj0_core_083;
  wire popcount25_1aj0_core_084;
  wire popcount25_1aj0_core_085;
  wire popcount25_1aj0_core_089;
  wire popcount25_1aj0_core_090;
  wire popcount25_1aj0_core_091;
  wire popcount25_1aj0_core_092;
  wire popcount25_1aj0_core_093;
  wire popcount25_1aj0_core_095;
  wire popcount25_1aj0_core_096;
  wire popcount25_1aj0_core_098;
  wire popcount25_1aj0_core_101;
  wire popcount25_1aj0_core_102;
  wire popcount25_1aj0_core_103;
  wire popcount25_1aj0_core_104;
  wire popcount25_1aj0_core_105;
  wire popcount25_1aj0_core_106;
  wire popcount25_1aj0_core_108;
  wire popcount25_1aj0_core_109;
  wire popcount25_1aj0_core_110;
  wire popcount25_1aj0_core_111;
  wire popcount25_1aj0_core_112;
  wire popcount25_1aj0_core_114;
  wire popcount25_1aj0_core_115_not;
  wire popcount25_1aj0_core_122;
  wire popcount25_1aj0_core_123;
  wire popcount25_1aj0_core_125;
  wire popcount25_1aj0_core_126;
  wire popcount25_1aj0_core_128;
  wire popcount25_1aj0_core_130;
  wire popcount25_1aj0_core_131;
  wire popcount25_1aj0_core_132;
  wire popcount25_1aj0_core_134;
  wire popcount25_1aj0_core_135;
  wire popcount25_1aj0_core_136;
  wire popcount25_1aj0_core_137;
  wire popcount25_1aj0_core_138;
  wire popcount25_1aj0_core_139;
  wire popcount25_1aj0_core_141;
  wire popcount25_1aj0_core_142;
  wire popcount25_1aj0_core_143;
  wire popcount25_1aj0_core_144;
  wire popcount25_1aj0_core_145;
  wire popcount25_1aj0_core_148;
  wire popcount25_1aj0_core_149;
  wire popcount25_1aj0_core_151;
  wire popcount25_1aj0_core_152;
  wire popcount25_1aj0_core_154;
  wire popcount25_1aj0_core_155;
  wire popcount25_1aj0_core_156;
  wire popcount25_1aj0_core_157_not;
  wire popcount25_1aj0_core_158;
  wire popcount25_1aj0_core_159;
  wire popcount25_1aj0_core_160;
  wire popcount25_1aj0_core_163;
  wire popcount25_1aj0_core_164;
  wire popcount25_1aj0_core_165_not;
  wire popcount25_1aj0_core_168;
  wire popcount25_1aj0_core_169;
  wire popcount25_1aj0_core_171;
  wire popcount25_1aj0_core_172;
  wire popcount25_1aj0_core_173;
  wire popcount25_1aj0_core_174;
  wire popcount25_1aj0_core_176;
  wire popcount25_1aj0_core_177;
  wire popcount25_1aj0_core_178;
  wire popcount25_1aj0_core_179;
  wire popcount25_1aj0_core_180;
  wire popcount25_1aj0_core_181;
  wire popcount25_1aj0_core_182;
  wire popcount25_1aj0_core_183;

  assign popcount25_1aj0_core_027 = input_a[8] & input_a[11];
  assign popcount25_1aj0_core_030 = input_a[5] ^ input_a[7];
  assign popcount25_1aj0_core_032 = ~input_a[4];
  assign popcount25_1aj0_core_035 = ~(input_a[7] & input_a[21]);
  assign popcount25_1aj0_core_037 = ~(input_a[2] & input_a[11]);
  assign popcount25_1aj0_core_038 = ~(input_a[24] & input_a[18]);
  assign popcount25_1aj0_core_040 = input_a[6] | input_a[9];
  assign popcount25_1aj0_core_041 = ~(input_a[9] ^ input_a[9]);
  assign popcount25_1aj0_core_044 = ~input_a[1];
  assign popcount25_1aj0_core_046 = ~(input_a[16] ^ input_a[6]);
  assign popcount25_1aj0_core_047 = input_a[5] & input_a[2];
  assign popcount25_1aj0_core_048 = input_a[8] | input_a[13];
  assign popcount25_1aj0_core_049 = input_a[1] | input_a[9];
  assign popcount25_1aj0_core_051 = ~(input_a[7] ^ input_a[1]);
  assign popcount25_1aj0_core_052 = input_a[9] ^ input_a[3];
  assign popcount25_1aj0_core_055 = input_a[24] | input_a[7];
  assign popcount25_1aj0_core_056_not = ~input_a[15];
  assign popcount25_1aj0_core_058 = ~input_a[9];
  assign popcount25_1aj0_core_059 = input_a[1] | input_a[0];
  assign popcount25_1aj0_core_061 = ~(input_a[18] & input_a[13]);
  assign popcount25_1aj0_core_062 = input_a[17] ^ input_a[10];
  assign popcount25_1aj0_core_063_not = ~input_a[19];
  assign popcount25_1aj0_core_064 = input_a[12] & input_a[24];
  assign popcount25_1aj0_core_066 = input_a[4] | input_a[23];
  assign popcount25_1aj0_core_067 = ~(input_a[3] & input_a[1]);
  assign popcount25_1aj0_core_070 = ~(input_a[23] ^ input_a[18]);
  assign popcount25_1aj0_core_072 = input_a[16] ^ input_a[1];
  assign popcount25_1aj0_core_073 = ~(input_a[7] & input_a[17]);
  assign popcount25_1aj0_core_074 = ~(input_a[19] ^ input_a[18]);
  assign popcount25_1aj0_core_075 = ~(input_a[12] & input_a[11]);
  assign popcount25_1aj0_core_076 = ~(input_a[16] | input_a[16]);
  assign popcount25_1aj0_core_077 = input_a[14] | input_a[9];
  assign popcount25_1aj0_core_080_not = ~input_a[7];
  assign popcount25_1aj0_core_081 = input_a[1] ^ input_a[24];
  assign popcount25_1aj0_core_082 = ~input_a[2];
  assign popcount25_1aj0_core_083 = input_a[5] ^ input_a[20];
  assign popcount25_1aj0_core_084 = ~(input_a[2] | input_a[17]);
  assign popcount25_1aj0_core_085 = ~(input_a[9] & input_a[9]);
  assign popcount25_1aj0_core_089 = ~(input_a[21] & input_a[15]);
  assign popcount25_1aj0_core_090 = input_a[5] | input_a[19];
  assign popcount25_1aj0_core_091 = input_a[23] | input_a[17];
  assign popcount25_1aj0_core_092 = input_a[24] ^ input_a[21];
  assign popcount25_1aj0_core_093 = ~(input_a[21] ^ input_a[4]);
  assign popcount25_1aj0_core_095 = input_a[21] | input_a[2];
  assign popcount25_1aj0_core_096 = input_a[18] ^ input_a[17];
  assign popcount25_1aj0_core_098 = input_a[19] ^ input_a[11];
  assign popcount25_1aj0_core_101 = ~(input_a[7] | input_a[22]);
  assign popcount25_1aj0_core_102 = ~(input_a[6] | input_a[24]);
  assign popcount25_1aj0_core_103 = ~(input_a[7] & input_a[3]);
  assign popcount25_1aj0_core_104 = input_a[11] | input_a[19];
  assign popcount25_1aj0_core_105 = input_a[9] ^ input_a[12];
  assign popcount25_1aj0_core_106 = ~(input_a[3] | input_a[1]);
  assign popcount25_1aj0_core_108 = ~(input_a[13] | input_a[23]);
  assign popcount25_1aj0_core_109 = ~(input_a[14] | input_a[17]);
  assign popcount25_1aj0_core_110 = ~(input_a[11] & input_a[12]);
  assign popcount25_1aj0_core_111 = ~(input_a[10] & input_a[21]);
  assign popcount25_1aj0_core_112 = ~input_a[20];
  assign popcount25_1aj0_core_114 = ~(input_a[15] | input_a[23]);
  assign popcount25_1aj0_core_115_not = ~input_a[5];
  assign popcount25_1aj0_core_122 = ~(input_a[14] | input_a[23]);
  assign popcount25_1aj0_core_123 = input_a[24] & input_a[4];
  assign popcount25_1aj0_core_125 = ~(input_a[1] | input_a[7]);
  assign popcount25_1aj0_core_126 = input_a[14] ^ input_a[10];
  assign popcount25_1aj0_core_128 = ~(input_a[24] | input_a[15]);
  assign popcount25_1aj0_core_130 = ~(input_a[0] | input_a[0]);
  assign popcount25_1aj0_core_131 = input_a[9] | input_a[19];
  assign popcount25_1aj0_core_132 = input_a[8] & input_a[21];
  assign popcount25_1aj0_core_134 = ~(input_a[8] & input_a[20]);
  assign popcount25_1aj0_core_135 = input_a[22] & input_a[12];
  assign popcount25_1aj0_core_136 = input_a[9] | input_a[18];
  assign popcount25_1aj0_core_137 = ~(input_a[9] | input_a[4]);
  assign popcount25_1aj0_core_138 = input_a[23] & input_a[13];
  assign popcount25_1aj0_core_139 = input_a[0] | input_a[15];
  assign popcount25_1aj0_core_141 = ~input_a[13];
  assign popcount25_1aj0_core_142 = input_a[9] & input_a[9];
  assign popcount25_1aj0_core_143 = input_a[16] ^ input_a[2];
  assign popcount25_1aj0_core_144 = input_a[2] & input_a[10];
  assign popcount25_1aj0_core_145 = input_a[17] & input_a[4];
  assign popcount25_1aj0_core_148 = ~(input_a[9] ^ input_a[6]);
  assign popcount25_1aj0_core_149 = ~(input_a[9] | input_a[10]);
  assign popcount25_1aj0_core_151 = input_a[24] & input_a[8];
  assign popcount25_1aj0_core_152 = ~(input_a[3] & input_a[2]);
  assign popcount25_1aj0_core_154 = input_a[14] | input_a[22];
  assign popcount25_1aj0_core_155 = ~input_a[5];
  assign popcount25_1aj0_core_156 = input_a[7] | input_a[10];
  assign popcount25_1aj0_core_157_not = ~input_a[11];
  assign popcount25_1aj0_core_158 = input_a[10] ^ input_a[18];
  assign popcount25_1aj0_core_159 = input_a[2] & input_a[6];
  assign popcount25_1aj0_core_160 = input_a[16] ^ input_a[18];
  assign popcount25_1aj0_core_163 = ~(input_a[7] | input_a[23]);
  assign popcount25_1aj0_core_164 = input_a[5] ^ input_a[6];
  assign popcount25_1aj0_core_165_not = ~input_a[16];
  assign popcount25_1aj0_core_168 = ~input_a[11];
  assign popcount25_1aj0_core_169 = ~(input_a[16] & input_a[2]);
  assign popcount25_1aj0_core_171 = ~(input_a[12] ^ input_a[11]);
  assign popcount25_1aj0_core_172 = ~(input_a[2] & input_a[12]);
  assign popcount25_1aj0_core_173 = input_a[14] | input_a[4];
  assign popcount25_1aj0_core_174 = ~(input_a[24] ^ input_a[4]);
  assign popcount25_1aj0_core_176 = input_a[23] & input_a[24];
  assign popcount25_1aj0_core_177 = ~input_a[4];
  assign popcount25_1aj0_core_178 = input_a[23] | input_a[23];
  assign popcount25_1aj0_core_179 = ~input_a[14];
  assign popcount25_1aj0_core_180 = input_a[9] & input_a[12];
  assign popcount25_1aj0_core_181 = ~(input_a[13] ^ input_a[18]);
  assign popcount25_1aj0_core_182 = input_a[2] & input_a[3];
  assign popcount25_1aj0_core_183 = input_a[20] | input_a[10];

  assign popcount25_1aj0_out[0] = input_a[2];
  assign popcount25_1aj0_out[1] = input_a[19];
  assign popcount25_1aj0_out[2] = input_a[12];
  assign popcount25_1aj0_out[3] = 1'b1;
  assign popcount25_1aj0_out[4] = 1'b0;
endmodule