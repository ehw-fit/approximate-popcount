// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.66647
// WCE=7.0
// EP=0.816452%
// Printed PDK parameters:
//  Area=70111209.0
//  Delay=83817832.0
//  Power=3370000.0

module popcount34_3vkq(input [33:0] input_a, output [5:0] popcount34_3vkq_out);
  wire popcount34_3vkq_core_036;
  wire popcount34_3vkq_core_037;
  wire popcount34_3vkq_core_040;
  wire popcount34_3vkq_core_041;
  wire popcount34_3vkq_core_042;
  wire popcount34_3vkq_core_043;
  wire popcount34_3vkq_core_047;
  wire popcount34_3vkq_core_048;
  wire popcount34_3vkq_core_049;
  wire popcount34_3vkq_core_051_not;
  wire popcount34_3vkq_core_052;
  wire popcount34_3vkq_core_054;
  wire popcount34_3vkq_core_056;
  wire popcount34_3vkq_core_057;
  wire popcount34_3vkq_core_058;
  wire popcount34_3vkq_core_059;
  wire popcount34_3vkq_core_061;
  wire popcount34_3vkq_core_062;
  wire popcount34_3vkq_core_063;
  wire popcount34_3vkq_core_065;
  wire popcount34_3vkq_core_066;
  wire popcount34_3vkq_core_068;
  wire popcount34_3vkq_core_070;
  wire popcount34_3vkq_core_071;
  wire popcount34_3vkq_core_072;
  wire popcount34_3vkq_core_073;
  wire popcount34_3vkq_core_074;
  wire popcount34_3vkq_core_075;
  wire popcount34_3vkq_core_076;
  wire popcount34_3vkq_core_077;
  wire popcount34_3vkq_core_078;
  wire popcount34_3vkq_core_081;
  wire popcount34_3vkq_core_083;
  wire popcount34_3vkq_core_085;
  wire popcount34_3vkq_core_086;
  wire popcount34_3vkq_core_087;
  wire popcount34_3vkq_core_088;
  wire popcount34_3vkq_core_089;
  wire popcount34_3vkq_core_090;
  wire popcount34_3vkq_core_092;
  wire popcount34_3vkq_core_093;
  wire popcount34_3vkq_core_094;
  wire popcount34_3vkq_core_096;
  wire popcount34_3vkq_core_098;
  wire popcount34_3vkq_core_102;
  wire popcount34_3vkq_core_103;
  wire popcount34_3vkq_core_106_not;
  wire popcount34_3vkq_core_107;
  wire popcount34_3vkq_core_108;
  wire popcount34_3vkq_core_109;
  wire popcount34_3vkq_core_110;
  wire popcount34_3vkq_core_112;
  wire popcount34_3vkq_core_113;
  wire popcount34_3vkq_core_114;
  wire popcount34_3vkq_core_115;
  wire popcount34_3vkq_core_116;
  wire popcount34_3vkq_core_117;
  wire popcount34_3vkq_core_118;
  wire popcount34_3vkq_core_119;
  wire popcount34_3vkq_core_120;
  wire popcount34_3vkq_core_121;
  wire popcount34_3vkq_core_122;
  wire popcount34_3vkq_core_123;
  wire popcount34_3vkq_core_126;
  wire popcount34_3vkq_core_127;
  wire popcount34_3vkq_core_130;
  wire popcount34_3vkq_core_131;
  wire popcount34_3vkq_core_132;
  wire popcount34_3vkq_core_133;
  wire popcount34_3vkq_core_134;
  wire popcount34_3vkq_core_135;
  wire popcount34_3vkq_core_136;
  wire popcount34_3vkq_core_137;
  wire popcount34_3vkq_core_138;
  wire popcount34_3vkq_core_139;
  wire popcount34_3vkq_core_140;
  wire popcount34_3vkq_core_143;
  wire popcount34_3vkq_core_144;
  wire popcount34_3vkq_core_145;
  wire popcount34_3vkq_core_147;
  wire popcount34_3vkq_core_148;
  wire popcount34_3vkq_core_149;
  wire popcount34_3vkq_core_153;
  wire popcount34_3vkq_core_154;
  wire popcount34_3vkq_core_155;
  wire popcount34_3vkq_core_156;
  wire popcount34_3vkq_core_157;
  wire popcount34_3vkq_core_158;
  wire popcount34_3vkq_core_159;
  wire popcount34_3vkq_core_160;
  wire popcount34_3vkq_core_161;
  wire popcount34_3vkq_core_162;
  wire popcount34_3vkq_core_163;
  wire popcount34_3vkq_core_166;
  wire popcount34_3vkq_core_167;
  wire popcount34_3vkq_core_168;
  wire popcount34_3vkq_core_169;
  wire popcount34_3vkq_core_170;
  wire popcount34_3vkq_core_171;
  wire popcount34_3vkq_core_172;
  wire popcount34_3vkq_core_176;
  wire popcount34_3vkq_core_177;
  wire popcount34_3vkq_core_178;
  wire popcount34_3vkq_core_179;
  wire popcount34_3vkq_core_180;
  wire popcount34_3vkq_core_181;
  wire popcount34_3vkq_core_182;
  wire popcount34_3vkq_core_184;
  wire popcount34_3vkq_core_185;
  wire popcount34_3vkq_core_186;
  wire popcount34_3vkq_core_187;
  wire popcount34_3vkq_core_188;
  wire popcount34_3vkq_core_189;
  wire popcount34_3vkq_core_190;
  wire popcount34_3vkq_core_193;
  wire popcount34_3vkq_core_194;
  wire popcount34_3vkq_core_195;
  wire popcount34_3vkq_core_196;
  wire popcount34_3vkq_core_198;
  wire popcount34_3vkq_core_199;
  wire popcount34_3vkq_core_200;
  wire popcount34_3vkq_core_201;
  wire popcount34_3vkq_core_202;
  wire popcount34_3vkq_core_203;
  wire popcount34_3vkq_core_204;
  wire popcount34_3vkq_core_208;
  wire popcount34_3vkq_core_209;
  wire popcount34_3vkq_core_211;
  wire popcount34_3vkq_core_212;
  wire popcount34_3vkq_core_213;
  wire popcount34_3vkq_core_214;
  wire popcount34_3vkq_core_215;
  wire popcount34_3vkq_core_216;
  wire popcount34_3vkq_core_217;
  wire popcount34_3vkq_core_218;
  wire popcount34_3vkq_core_219;
  wire popcount34_3vkq_core_220;
  wire popcount34_3vkq_core_221;
  wire popcount34_3vkq_core_222;
  wire popcount34_3vkq_core_223;
  wire popcount34_3vkq_core_225;
  wire popcount34_3vkq_core_226;
  wire popcount34_3vkq_core_227;
  wire popcount34_3vkq_core_228;
  wire popcount34_3vkq_core_229;
  wire popcount34_3vkq_core_230;
  wire popcount34_3vkq_core_231;
  wire popcount34_3vkq_core_233;
  wire popcount34_3vkq_core_234;
  wire popcount34_3vkq_core_235;
  wire popcount34_3vkq_core_236;
  wire popcount34_3vkq_core_237;
  wire popcount34_3vkq_core_238;
  wire popcount34_3vkq_core_239;
  wire popcount34_3vkq_core_240;
  wire popcount34_3vkq_core_241;
  wire popcount34_3vkq_core_242;
  wire popcount34_3vkq_core_243;
  wire popcount34_3vkq_core_244;
  wire popcount34_3vkq_core_245;
  wire popcount34_3vkq_core_246;
  wire popcount34_3vkq_core_247;
  wire popcount34_3vkq_core_248;
  wire popcount34_3vkq_core_249;
  wire popcount34_3vkq_core_250;
  wire popcount34_3vkq_core_251;

  assign popcount34_3vkq_core_036 = ~(input_a[33] | input_a[22]);
  assign popcount34_3vkq_core_037 = input_a[0] & input_a[1];
  assign popcount34_3vkq_core_040 = input_a[11] | input_a[9];
  assign popcount34_3vkq_core_041 = ~input_a[19];
  assign popcount34_3vkq_core_042 = ~input_a[33];
  assign popcount34_3vkq_core_043 = popcount34_3vkq_core_037 & input_a[4];
  assign popcount34_3vkq_core_047 = ~(input_a[27] | input_a[13]);
  assign popcount34_3vkq_core_048 = ~(input_a[25] & input_a[22]);
  assign popcount34_3vkq_core_049 = input_a[18] ^ input_a[14];
  assign popcount34_3vkq_core_051_not = ~input_a[8];
  assign popcount34_3vkq_core_052 = input_a[5] & input_a[22];
  assign popcount34_3vkq_core_054 = input_a[33] & input_a[14];
  assign popcount34_3vkq_core_056 = input_a[11] ^ input_a[14];
  assign popcount34_3vkq_core_057 = ~input_a[14];
  assign popcount34_3vkq_core_058 = ~(input_a[24] ^ input_a[18]);
  assign popcount34_3vkq_core_059 = input_a[12] & input_a[14];
  assign popcount34_3vkq_core_061 = ~input_a[25];
  assign popcount34_3vkq_core_062 = popcount34_3vkq_core_052 | popcount34_3vkq_core_059;
  assign popcount34_3vkq_core_063 = ~(input_a[3] | input_a[5]);
  assign popcount34_3vkq_core_065 = ~(popcount34_3vkq_core_043 & input_a[3]);
  assign popcount34_3vkq_core_066 = popcount34_3vkq_core_043 & input_a[3];
  assign popcount34_3vkq_core_068 = input_a[32] ^ input_a[17];
  assign popcount34_3vkq_core_070 = input_a[8] ^ input_a[9];
  assign popcount34_3vkq_core_071 = input_a[8] & input_a[9];
  assign popcount34_3vkq_core_072 = input_a[10] ^ input_a[11];
  assign popcount34_3vkq_core_073 = input_a[10] & input_a[11];
  assign popcount34_3vkq_core_074 = popcount34_3vkq_core_070 ^ popcount34_3vkq_core_072;
  assign popcount34_3vkq_core_075 = popcount34_3vkq_core_070 & popcount34_3vkq_core_072;
  assign popcount34_3vkq_core_076 = popcount34_3vkq_core_071 ^ popcount34_3vkq_core_073;
  assign popcount34_3vkq_core_077 = popcount34_3vkq_core_071 & input_a[10];
  assign popcount34_3vkq_core_078 = popcount34_3vkq_core_076 | popcount34_3vkq_core_075;
  assign popcount34_3vkq_core_081 = ~input_a[16];
  assign popcount34_3vkq_core_083 = ~(input_a[4] | input_a[30]);
  assign popcount34_3vkq_core_085 = input_a[28] | input_a[17];
  assign popcount34_3vkq_core_086 = ~(input_a[17] & input_a[26]);
  assign popcount34_3vkq_core_087 = input_a[10] ^ input_a[30];
  assign popcount34_3vkq_core_088 = ~(input_a[7] ^ input_a[22]);
  assign popcount34_3vkq_core_089 = input_a[31] ^ input_a[30];
  assign popcount34_3vkq_core_090 = input_a[11] | input_a[24];
  assign popcount34_3vkq_core_092 = input_a[25] ^ input_a[16];
  assign popcount34_3vkq_core_093 = ~(input_a[18] | input_a[5]);
  assign popcount34_3vkq_core_094 = input_a[17] & input_a[6];
  assign popcount34_3vkq_core_096 = input_a[14] | input_a[24];
  assign popcount34_3vkq_core_098 = ~popcount34_3vkq_core_074;
  assign popcount34_3vkq_core_102 = popcount34_3vkq_core_078 ^ popcount34_3vkq_core_074;
  assign popcount34_3vkq_core_103 = popcount34_3vkq_core_078 & popcount34_3vkq_core_074;
  assign popcount34_3vkq_core_106_not = ~input_a[16];
  assign popcount34_3vkq_core_107 = popcount34_3vkq_core_077 | popcount34_3vkq_core_103;
  assign popcount34_3vkq_core_108 = ~(input_a[33] ^ input_a[7]);
  assign popcount34_3vkq_core_109 = input_a[3] | input_a[23];
  assign popcount34_3vkq_core_110 = ~input_a[9];
  assign popcount34_3vkq_core_112 = ~(input_a[15] | input_a[16]);
  assign popcount34_3vkq_core_113 = input_a[15] & popcount34_3vkq_core_098;
  assign popcount34_3vkq_core_114 = popcount34_3vkq_core_062 ^ popcount34_3vkq_core_102;
  assign popcount34_3vkq_core_115 = popcount34_3vkq_core_062 & popcount34_3vkq_core_102;
  assign popcount34_3vkq_core_116 = popcount34_3vkq_core_114 ^ popcount34_3vkq_core_113;
  assign popcount34_3vkq_core_117 = popcount34_3vkq_core_114 & popcount34_3vkq_core_113;
  assign popcount34_3vkq_core_118 = popcount34_3vkq_core_115 | popcount34_3vkq_core_117;
  assign popcount34_3vkq_core_119 = popcount34_3vkq_core_065 ^ popcount34_3vkq_core_107;
  assign popcount34_3vkq_core_120 = popcount34_3vkq_core_065 & popcount34_3vkq_core_107;
  assign popcount34_3vkq_core_121 = popcount34_3vkq_core_119 ^ popcount34_3vkq_core_118;
  assign popcount34_3vkq_core_122 = popcount34_3vkq_core_119 & popcount34_3vkq_core_118;
  assign popcount34_3vkq_core_123 = popcount34_3vkq_core_120 | popcount34_3vkq_core_122;
  assign popcount34_3vkq_core_126 = popcount34_3vkq_core_066 ^ popcount34_3vkq_core_123;
  assign popcount34_3vkq_core_127 = popcount34_3vkq_core_066 & popcount34_3vkq_core_123;
  assign popcount34_3vkq_core_130 = ~(input_a[11] ^ input_a[5]);
  assign popcount34_3vkq_core_131 = input_a[17] ^ input_a[18];
  assign popcount34_3vkq_core_132 = input_a[17] & input_a[18];
  assign popcount34_3vkq_core_133 = input_a[19] ^ input_a[20];
  assign popcount34_3vkq_core_134 = input_a[19] & input_a[20];
  assign popcount34_3vkq_core_135 = popcount34_3vkq_core_131 ^ popcount34_3vkq_core_133;
  assign popcount34_3vkq_core_136 = popcount34_3vkq_core_131 & popcount34_3vkq_core_133;
  assign popcount34_3vkq_core_137 = popcount34_3vkq_core_132 ^ popcount34_3vkq_core_134;
  assign popcount34_3vkq_core_138 = popcount34_3vkq_core_132 & popcount34_3vkq_core_134;
  assign popcount34_3vkq_core_139 = popcount34_3vkq_core_137 | popcount34_3vkq_core_136;
  assign popcount34_3vkq_core_140 = input_a[16] ^ input_a[14];
  assign popcount34_3vkq_core_143 = input_a[21] & input_a[6];
  assign popcount34_3vkq_core_144 = input_a[23] ^ input_a[24];
  assign popcount34_3vkq_core_145 = input_a[23] & input_a[24];
  assign popcount34_3vkq_core_147 = input_a[13] ^ input_a[33];
  assign popcount34_3vkq_core_148 = popcount34_3vkq_core_143 ^ popcount34_3vkq_core_145;
  assign popcount34_3vkq_core_149 = popcount34_3vkq_core_143 & popcount34_3vkq_core_145;
  assign popcount34_3vkq_core_153 = input_a[5] & input_a[9];
  assign popcount34_3vkq_core_154 = popcount34_3vkq_core_135 & popcount34_3vkq_core_144;
  assign popcount34_3vkq_core_155 = popcount34_3vkq_core_139 ^ popcount34_3vkq_core_148;
  assign popcount34_3vkq_core_156 = popcount34_3vkq_core_139 & popcount34_3vkq_core_148;
  assign popcount34_3vkq_core_157 = popcount34_3vkq_core_155 ^ popcount34_3vkq_core_154;
  assign popcount34_3vkq_core_158 = popcount34_3vkq_core_155 & popcount34_3vkq_core_154;
  assign popcount34_3vkq_core_159 = popcount34_3vkq_core_156 | popcount34_3vkq_core_158;
  assign popcount34_3vkq_core_160 = popcount34_3vkq_core_138 ^ popcount34_3vkq_core_149;
  assign popcount34_3vkq_core_161 = popcount34_3vkq_core_138 & popcount34_3vkq_core_149;
  assign popcount34_3vkq_core_162 = popcount34_3vkq_core_160 | popcount34_3vkq_core_159;
  assign popcount34_3vkq_core_163 = input_a[12] ^ input_a[23];
  assign popcount34_3vkq_core_166 = input_a[27] & input_a[2];
  assign popcount34_3vkq_core_167 = input_a[30] ^ input_a[19];
  assign popcount34_3vkq_core_168 = input_a[26] & input_a[28];
  assign popcount34_3vkq_core_169 = input_a[33] ^ input_a[22];
  assign popcount34_3vkq_core_170 = input_a[24] & input_a[0];
  assign popcount34_3vkq_core_171 = popcount34_3vkq_core_166 ^ popcount34_3vkq_core_168;
  assign popcount34_3vkq_core_172 = popcount34_3vkq_core_166 & popcount34_3vkq_core_168;
  assign popcount34_3vkq_core_176 = input_a[29] ^ input_a[30];
  assign popcount34_3vkq_core_177 = input_a[29] & input_a[30];
  assign popcount34_3vkq_core_178 = input_a[32] ^ input_a[33];
  assign popcount34_3vkq_core_179 = input_a[32] & input_a[33];
  assign popcount34_3vkq_core_180 = input_a[31] ^ popcount34_3vkq_core_178;
  assign popcount34_3vkq_core_181 = input_a[31] & popcount34_3vkq_core_178;
  assign popcount34_3vkq_core_182 = popcount34_3vkq_core_179 | popcount34_3vkq_core_181;
  assign popcount34_3vkq_core_184 = popcount34_3vkq_core_176 ^ popcount34_3vkq_core_180;
  assign popcount34_3vkq_core_185 = popcount34_3vkq_core_176 & popcount34_3vkq_core_180;
  assign popcount34_3vkq_core_186 = popcount34_3vkq_core_177 ^ popcount34_3vkq_core_182;
  assign popcount34_3vkq_core_187 = popcount34_3vkq_core_177 & popcount34_3vkq_core_182;
  assign popcount34_3vkq_core_188 = popcount34_3vkq_core_186 ^ popcount34_3vkq_core_185;
  assign popcount34_3vkq_core_189 = popcount34_3vkq_core_186 & popcount34_3vkq_core_185;
  assign popcount34_3vkq_core_190 = popcount34_3vkq_core_187 | popcount34_3vkq_core_189;
  assign popcount34_3vkq_core_193 = ~(input_a[21] ^ input_a[11]);
  assign popcount34_3vkq_core_194 = input_a[16] & popcount34_3vkq_core_184;
  assign popcount34_3vkq_core_195 = popcount34_3vkq_core_171 | popcount34_3vkq_core_188;
  assign popcount34_3vkq_core_196 = popcount34_3vkq_core_171 & popcount34_3vkq_core_188;
  assign popcount34_3vkq_core_198 = popcount34_3vkq_core_195 & popcount34_3vkq_core_194;
  assign popcount34_3vkq_core_199 = popcount34_3vkq_core_196 | popcount34_3vkq_core_198;
  assign popcount34_3vkq_core_200 = popcount34_3vkq_core_172 ^ popcount34_3vkq_core_190;
  assign popcount34_3vkq_core_201 = popcount34_3vkq_core_172 & popcount34_3vkq_core_190;
  assign popcount34_3vkq_core_202 = popcount34_3vkq_core_200 ^ popcount34_3vkq_core_199;
  assign popcount34_3vkq_core_203 = popcount34_3vkq_core_200 & popcount34_3vkq_core_199;
  assign popcount34_3vkq_core_204 = popcount34_3vkq_core_201 | popcount34_3vkq_core_203;
  assign popcount34_3vkq_core_208 = input_a[7] & input_a[25];
  assign popcount34_3vkq_core_209 = ~popcount34_3vkq_core_157;
  assign popcount34_3vkq_core_211 = popcount34_3vkq_core_209 ^ popcount34_3vkq_core_208;
  assign popcount34_3vkq_core_212 = input_a[7] & input_a[25];
  assign popcount34_3vkq_core_213 = popcount34_3vkq_core_157 | popcount34_3vkq_core_212;
  assign popcount34_3vkq_core_214 = popcount34_3vkq_core_162 ^ popcount34_3vkq_core_202;
  assign popcount34_3vkq_core_215 = popcount34_3vkq_core_162 & popcount34_3vkq_core_202;
  assign popcount34_3vkq_core_216 = popcount34_3vkq_core_214 ^ popcount34_3vkq_core_213;
  assign popcount34_3vkq_core_217 = popcount34_3vkq_core_214 & popcount34_3vkq_core_213;
  assign popcount34_3vkq_core_218 = popcount34_3vkq_core_215 | popcount34_3vkq_core_217;
  assign popcount34_3vkq_core_219 = popcount34_3vkq_core_161 ^ popcount34_3vkq_core_204;
  assign popcount34_3vkq_core_220 = popcount34_3vkq_core_161 & popcount34_3vkq_core_204;
  assign popcount34_3vkq_core_221 = popcount34_3vkq_core_219 ^ popcount34_3vkq_core_218;
  assign popcount34_3vkq_core_222 = popcount34_3vkq_core_219 & popcount34_3vkq_core_218;
  assign popcount34_3vkq_core_223 = popcount34_3vkq_core_220 | popcount34_3vkq_core_222;
  assign popcount34_3vkq_core_225 = ~(input_a[4] & input_a[23]);
  assign popcount34_3vkq_core_226 = input_a[11] | input_a[3];
  assign popcount34_3vkq_core_227 = ~(input_a[18] | input_a[2]);
  assign popcount34_3vkq_core_228 = popcount34_3vkq_core_116 ^ popcount34_3vkq_core_211;
  assign popcount34_3vkq_core_229 = popcount34_3vkq_core_116 & popcount34_3vkq_core_211;
  assign popcount34_3vkq_core_230 = ~(input_a[25] ^ input_a[24]);
  assign popcount34_3vkq_core_231 = ~(input_a[22] & input_a[33]);
  assign popcount34_3vkq_core_233 = popcount34_3vkq_core_121 ^ popcount34_3vkq_core_216;
  assign popcount34_3vkq_core_234 = popcount34_3vkq_core_121 & popcount34_3vkq_core_216;
  assign popcount34_3vkq_core_235 = popcount34_3vkq_core_233 ^ popcount34_3vkq_core_229;
  assign popcount34_3vkq_core_236 = popcount34_3vkq_core_233 & popcount34_3vkq_core_229;
  assign popcount34_3vkq_core_237 = popcount34_3vkq_core_234 | popcount34_3vkq_core_236;
  assign popcount34_3vkq_core_238 = popcount34_3vkq_core_126 ^ popcount34_3vkq_core_221;
  assign popcount34_3vkq_core_239 = popcount34_3vkq_core_126 & popcount34_3vkq_core_221;
  assign popcount34_3vkq_core_240 = popcount34_3vkq_core_238 ^ popcount34_3vkq_core_237;
  assign popcount34_3vkq_core_241 = popcount34_3vkq_core_238 & popcount34_3vkq_core_237;
  assign popcount34_3vkq_core_242 = popcount34_3vkq_core_239 | popcount34_3vkq_core_241;
  assign popcount34_3vkq_core_243 = popcount34_3vkq_core_127 ^ popcount34_3vkq_core_223;
  assign popcount34_3vkq_core_244 = popcount34_3vkq_core_127 & popcount34_3vkq_core_223;
  assign popcount34_3vkq_core_245 = popcount34_3vkq_core_243 ^ popcount34_3vkq_core_242;
  assign popcount34_3vkq_core_246 = popcount34_3vkq_core_243 & popcount34_3vkq_core_242;
  assign popcount34_3vkq_core_247 = popcount34_3vkq_core_244 | popcount34_3vkq_core_246;
  assign popcount34_3vkq_core_248 = ~input_a[31];
  assign popcount34_3vkq_core_249 = input_a[8] & input_a[15];
  assign popcount34_3vkq_core_250 = input_a[30] & input_a[9];
  assign popcount34_3vkq_core_251 = ~input_a[2];

  assign popcount34_3vkq_out[0] = input_a[13];
  assign popcount34_3vkq_out[1] = popcount34_3vkq_core_228;
  assign popcount34_3vkq_out[2] = popcount34_3vkq_core_235;
  assign popcount34_3vkq_out[3] = popcount34_3vkq_core_240;
  assign popcount34_3vkq_out[4] = popcount34_3vkq_core_245;
  assign popcount34_3vkq_out[5] = popcount34_3vkq_core_247;
endmodule