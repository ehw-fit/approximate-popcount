// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.72677
// WCE=17.0
// EP=0.888465%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_s2ta(input [28:0] input_a, output [4:0] popcount29_s2ta_out);
  wire popcount29_s2ta_core_031;
  wire popcount29_s2ta_core_032;
  wire popcount29_s2ta_core_035;
  wire popcount29_s2ta_core_036;
  wire popcount29_s2ta_core_038;
  wire popcount29_s2ta_core_039;
  wire popcount29_s2ta_core_040;
  wire popcount29_s2ta_core_042_not;
  wire popcount29_s2ta_core_044;
  wire popcount29_s2ta_core_045;
  wire popcount29_s2ta_core_047;
  wire popcount29_s2ta_core_051;
  wire popcount29_s2ta_core_052;
  wire popcount29_s2ta_core_053;
  wire popcount29_s2ta_core_055;
  wire popcount29_s2ta_core_056;
  wire popcount29_s2ta_core_057;
  wire popcount29_s2ta_core_058;
  wire popcount29_s2ta_core_059;
  wire popcount29_s2ta_core_060;
  wire popcount29_s2ta_core_061;
  wire popcount29_s2ta_core_062;
  wire popcount29_s2ta_core_063;
  wire popcount29_s2ta_core_064;
  wire popcount29_s2ta_core_065;
  wire popcount29_s2ta_core_066;
  wire popcount29_s2ta_core_067;
  wire popcount29_s2ta_core_068;
  wire popcount29_s2ta_core_069;
  wire popcount29_s2ta_core_070;
  wire popcount29_s2ta_core_074;
  wire popcount29_s2ta_core_075;
  wire popcount29_s2ta_core_076;
  wire popcount29_s2ta_core_077;
  wire popcount29_s2ta_core_078;
  wire popcount29_s2ta_core_079;
  wire popcount29_s2ta_core_080;
  wire popcount29_s2ta_core_081;
  wire popcount29_s2ta_core_083;
  wire popcount29_s2ta_core_084;
  wire popcount29_s2ta_core_085;
  wire popcount29_s2ta_core_086;
  wire popcount29_s2ta_core_089;
  wire popcount29_s2ta_core_092;
  wire popcount29_s2ta_core_094;
  wire popcount29_s2ta_core_095;
  wire popcount29_s2ta_core_099;
  wire popcount29_s2ta_core_100;
  wire popcount29_s2ta_core_101;
  wire popcount29_s2ta_core_104;
  wire popcount29_s2ta_core_106;
  wire popcount29_s2ta_core_107;
  wire popcount29_s2ta_core_109;
  wire popcount29_s2ta_core_110;
  wire popcount29_s2ta_core_111;
  wire popcount29_s2ta_core_112;
  wire popcount29_s2ta_core_113;
  wire popcount29_s2ta_core_114;
  wire popcount29_s2ta_core_115;
  wire popcount29_s2ta_core_116;
  wire popcount29_s2ta_core_117;
  wire popcount29_s2ta_core_119;
  wire popcount29_s2ta_core_122;
  wire popcount29_s2ta_core_126;
  wire popcount29_s2ta_core_128;
  wire popcount29_s2ta_core_130;
  wire popcount29_s2ta_core_134;
  wire popcount29_s2ta_core_135;
  wire popcount29_s2ta_core_136;
  wire popcount29_s2ta_core_137;
  wire popcount29_s2ta_core_139_not;
  wire popcount29_s2ta_core_140;
  wire popcount29_s2ta_core_141;
  wire popcount29_s2ta_core_142;
  wire popcount29_s2ta_core_144;
  wire popcount29_s2ta_core_145;
  wire popcount29_s2ta_core_147;
  wire popcount29_s2ta_core_150;
  wire popcount29_s2ta_core_151_not;
  wire popcount29_s2ta_core_152;
  wire popcount29_s2ta_core_155;
  wire popcount29_s2ta_core_156;
  wire popcount29_s2ta_core_158;
  wire popcount29_s2ta_core_159_not;
  wire popcount29_s2ta_core_160;
  wire popcount29_s2ta_core_161;
  wire popcount29_s2ta_core_163;
  wire popcount29_s2ta_core_165;
  wire popcount29_s2ta_core_168;
  wire popcount29_s2ta_core_169;
  wire popcount29_s2ta_core_170;
  wire popcount29_s2ta_core_171;
  wire popcount29_s2ta_core_172;
  wire popcount29_s2ta_core_178;
  wire popcount29_s2ta_core_179_not;
  wire popcount29_s2ta_core_182;
  wire popcount29_s2ta_core_183;
  wire popcount29_s2ta_core_184;
  wire popcount29_s2ta_core_185_not;
  wire popcount29_s2ta_core_186;
  wire popcount29_s2ta_core_187;
  wire popcount29_s2ta_core_188;
  wire popcount29_s2ta_core_189;
  wire popcount29_s2ta_core_191;
  wire popcount29_s2ta_core_192;
  wire popcount29_s2ta_core_193_not;
  wire popcount29_s2ta_core_194_not;
  wire popcount29_s2ta_core_195;
  wire popcount29_s2ta_core_196;
  wire popcount29_s2ta_core_197;
  wire popcount29_s2ta_core_199_not;
  wire popcount29_s2ta_core_200;
  wire popcount29_s2ta_core_203;
  wire popcount29_s2ta_core_204;
  wire popcount29_s2ta_core_206;
  wire popcount29_s2ta_core_207;

  assign popcount29_s2ta_core_031 = ~input_a[13];
  assign popcount29_s2ta_core_032 = ~input_a[18];
  assign popcount29_s2ta_core_035 = ~(input_a[5] | input_a[24]);
  assign popcount29_s2ta_core_036 = ~(input_a[12] ^ input_a[18]);
  assign popcount29_s2ta_core_038 = ~input_a[14];
  assign popcount29_s2ta_core_039 = ~input_a[0];
  assign popcount29_s2ta_core_040 = input_a[19] & input_a[20];
  assign popcount29_s2ta_core_042_not = ~input_a[21];
  assign popcount29_s2ta_core_044 = ~(input_a[22] | input_a[12]);
  assign popcount29_s2ta_core_045 = ~(input_a[24] ^ input_a[20]);
  assign popcount29_s2ta_core_047 = input_a[27] | input_a[13];
  assign popcount29_s2ta_core_051 = ~(input_a[1] ^ input_a[0]);
  assign popcount29_s2ta_core_052 = input_a[28] & input_a[15];
  assign popcount29_s2ta_core_053 = input_a[3] ^ input_a[0];
  assign popcount29_s2ta_core_055 = ~(input_a[5] ^ input_a[5]);
  assign popcount29_s2ta_core_056 = input_a[23] ^ input_a[19];
  assign popcount29_s2ta_core_057 = input_a[0] | input_a[6];
  assign popcount29_s2ta_core_058 = ~input_a[6];
  assign popcount29_s2ta_core_059 = ~input_a[5];
  assign popcount29_s2ta_core_060 = input_a[23] & input_a[4];
  assign popcount29_s2ta_core_061 = input_a[5] | input_a[15];
  assign popcount29_s2ta_core_062 = ~(input_a[27] & input_a[18]);
  assign popcount29_s2ta_core_063 = input_a[16] ^ input_a[24];
  assign popcount29_s2ta_core_064 = ~(input_a[20] | input_a[14]);
  assign popcount29_s2ta_core_065 = input_a[0] | input_a[10];
  assign popcount29_s2ta_core_066 = ~(input_a[1] ^ input_a[9]);
  assign popcount29_s2ta_core_067 = ~input_a[22];
  assign popcount29_s2ta_core_068 = ~(input_a[21] ^ input_a[14]);
  assign popcount29_s2ta_core_069 = input_a[18] ^ input_a[20];
  assign popcount29_s2ta_core_070 = ~(input_a[12] ^ input_a[27]);
  assign popcount29_s2ta_core_074 = ~(input_a[23] | input_a[6]);
  assign popcount29_s2ta_core_075 = input_a[28] & input_a[7];
  assign popcount29_s2ta_core_076 = input_a[6] | input_a[1];
  assign popcount29_s2ta_core_077 = ~(input_a[5] & input_a[19]);
  assign popcount29_s2ta_core_078 = input_a[16] ^ input_a[25];
  assign popcount29_s2ta_core_079 = ~(input_a[1] | input_a[26]);
  assign popcount29_s2ta_core_080 = ~(input_a[13] | input_a[15]);
  assign popcount29_s2ta_core_081 = input_a[26] ^ input_a[7];
  assign popcount29_s2ta_core_083 = ~(input_a[14] | input_a[20]);
  assign popcount29_s2ta_core_084 = ~(input_a[19] | input_a[3]);
  assign popcount29_s2ta_core_085 = input_a[20] & input_a[26];
  assign popcount29_s2ta_core_086 = ~(input_a[15] ^ input_a[1]);
  assign popcount29_s2ta_core_089 = ~(input_a[3] & input_a[3]);
  assign popcount29_s2ta_core_092 = ~input_a[22];
  assign popcount29_s2ta_core_094 = input_a[12] ^ input_a[9];
  assign popcount29_s2ta_core_095 = ~(input_a[28] ^ input_a[18]);
  assign popcount29_s2ta_core_099 = ~(input_a[7] ^ input_a[21]);
  assign popcount29_s2ta_core_100 = input_a[0] & input_a[20];
  assign popcount29_s2ta_core_101 = input_a[2] & input_a[1];
  assign popcount29_s2ta_core_104 = ~input_a[24];
  assign popcount29_s2ta_core_106 = input_a[6] & input_a[20];
  assign popcount29_s2ta_core_107 = input_a[3] & input_a[5];
  assign popcount29_s2ta_core_109 = input_a[1] ^ input_a[8];
  assign popcount29_s2ta_core_110 = input_a[23] | input_a[3];
  assign popcount29_s2ta_core_111 = input_a[18] ^ input_a[17];
  assign popcount29_s2ta_core_112 = input_a[4] | input_a[14];
  assign popcount29_s2ta_core_113 = input_a[13] ^ input_a[28];
  assign popcount29_s2ta_core_114 = ~input_a[15];
  assign popcount29_s2ta_core_115 = input_a[24] ^ input_a[27];
  assign popcount29_s2ta_core_116 = input_a[20] | input_a[21];
  assign popcount29_s2ta_core_117 = input_a[25] ^ input_a[3];
  assign popcount29_s2ta_core_119 = ~(input_a[8] & input_a[16]);
  assign popcount29_s2ta_core_122 = ~(input_a[23] & input_a[9]);
  assign popcount29_s2ta_core_126 = ~(input_a[15] & input_a[10]);
  assign popcount29_s2ta_core_128 = ~input_a[3];
  assign popcount29_s2ta_core_130 = input_a[27] & input_a[22];
  assign popcount29_s2ta_core_134 = ~(input_a[23] ^ input_a[16]);
  assign popcount29_s2ta_core_135 = input_a[0] & input_a[26];
  assign popcount29_s2ta_core_136 = ~(input_a[16] ^ input_a[0]);
  assign popcount29_s2ta_core_137 = ~input_a[27];
  assign popcount29_s2ta_core_139_not = ~input_a[20];
  assign popcount29_s2ta_core_140 = ~(input_a[4] & input_a[19]);
  assign popcount29_s2ta_core_141 = ~(input_a[4] & input_a[17]);
  assign popcount29_s2ta_core_142 = ~(input_a[1] ^ input_a[10]);
  assign popcount29_s2ta_core_144 = input_a[16] ^ input_a[15];
  assign popcount29_s2ta_core_145 = ~input_a[15];
  assign popcount29_s2ta_core_147 = input_a[2] & input_a[3];
  assign popcount29_s2ta_core_150 = input_a[28] & input_a[23];
  assign popcount29_s2ta_core_151_not = ~input_a[15];
  assign popcount29_s2ta_core_152 = input_a[14] | input_a[11];
  assign popcount29_s2ta_core_155 = ~(input_a[8] & input_a[23]);
  assign popcount29_s2ta_core_156 = ~(input_a[9] | input_a[0]);
  assign popcount29_s2ta_core_158 = input_a[21] & input_a[10];
  assign popcount29_s2ta_core_159_not = ~input_a[19];
  assign popcount29_s2ta_core_160 = ~(input_a[4] & input_a[1]);
  assign popcount29_s2ta_core_161 = ~(input_a[23] ^ input_a[14]);
  assign popcount29_s2ta_core_163 = ~(input_a[9] & input_a[24]);
  assign popcount29_s2ta_core_165 = ~(input_a[21] & input_a[4]);
  assign popcount29_s2ta_core_168 = ~(input_a[24] ^ input_a[10]);
  assign popcount29_s2ta_core_169 = input_a[28] ^ input_a[21];
  assign popcount29_s2ta_core_170 = ~input_a[15];
  assign popcount29_s2ta_core_171 = ~(input_a[14] | input_a[2]);
  assign popcount29_s2ta_core_172 = ~(input_a[14] | input_a[8]);
  assign popcount29_s2ta_core_178 = input_a[1] | input_a[18];
  assign popcount29_s2ta_core_179_not = ~input_a[5];
  assign popcount29_s2ta_core_182 = input_a[19] ^ input_a[16];
  assign popcount29_s2ta_core_183 = input_a[3] & input_a[26];
  assign popcount29_s2ta_core_184 = ~(input_a[12] & input_a[1]);
  assign popcount29_s2ta_core_185_not = ~input_a[13];
  assign popcount29_s2ta_core_186 = input_a[13] | input_a[3];
  assign popcount29_s2ta_core_187 = input_a[9] | input_a[5];
  assign popcount29_s2ta_core_188 = ~(input_a[6] ^ input_a[8]);
  assign popcount29_s2ta_core_189 = input_a[27] & input_a[15];
  assign popcount29_s2ta_core_191 = input_a[3] | input_a[18];
  assign popcount29_s2ta_core_192 = ~(input_a[23] | input_a[27]);
  assign popcount29_s2ta_core_193_not = ~input_a[24];
  assign popcount29_s2ta_core_194_not = ~input_a[6];
  assign popcount29_s2ta_core_195 = ~(input_a[16] | input_a[3]);
  assign popcount29_s2ta_core_196 = ~input_a[24];
  assign popcount29_s2ta_core_197 = ~(input_a[26] ^ input_a[13]);
  assign popcount29_s2ta_core_199_not = ~input_a[26];
  assign popcount29_s2ta_core_200 = ~(input_a[27] ^ input_a[18]);
  assign popcount29_s2ta_core_203 = input_a[2] & input_a[14];
  assign popcount29_s2ta_core_204 = ~(input_a[5] & input_a[12]);
  assign popcount29_s2ta_core_206 = ~(input_a[13] & input_a[18]);
  assign popcount29_s2ta_core_207 = ~input_a[0];

  assign popcount29_s2ta_out[0] = 1'b1;
  assign popcount29_s2ta_out[1] = 1'b0;
  assign popcount29_s2ta_out[2] = 1'b0;
  assign popcount29_s2ta_out[3] = 1'b0;
  assign popcount29_s2ta_out[4] = 1'b1;
endmodule