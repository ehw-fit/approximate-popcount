// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.16697
// WCE=15.0
// EP=0.855536%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount30_rptt(input [29:0] input_a, output [4:0] popcount30_rptt_out);
  wire popcount30_rptt_core_032;
  wire popcount30_rptt_core_034;
  wire popcount30_rptt_core_035;
  wire popcount30_rptt_core_036;
  wire popcount30_rptt_core_037;
  wire popcount30_rptt_core_038;
  wire popcount30_rptt_core_039;
  wire popcount30_rptt_core_041;
  wire popcount30_rptt_core_043_not;
  wire popcount30_rptt_core_044;
  wire popcount30_rptt_core_046;
  wire popcount30_rptt_core_047;
  wire popcount30_rptt_core_052;
  wire popcount30_rptt_core_053;
  wire popcount30_rptt_core_054;
  wire popcount30_rptt_core_055;
  wire popcount30_rptt_core_057_not;
  wire popcount30_rptt_core_060;
  wire popcount30_rptt_core_062;
  wire popcount30_rptt_core_064;
  wire popcount30_rptt_core_065;
  wire popcount30_rptt_core_068;
  wire popcount30_rptt_core_069;
  wire popcount30_rptt_core_071;
  wire popcount30_rptt_core_072;
  wire popcount30_rptt_core_073;
  wire popcount30_rptt_core_074;
  wire popcount30_rptt_core_076;
  wire popcount30_rptt_core_078;
  wire popcount30_rptt_core_079;
  wire popcount30_rptt_core_080;
  wire popcount30_rptt_core_081;
  wire popcount30_rptt_core_083;
  wire popcount30_rptt_core_084;
  wire popcount30_rptt_core_085_not;
  wire popcount30_rptt_core_087;
  wire popcount30_rptt_core_088;
  wire popcount30_rptt_core_090;
  wire popcount30_rptt_core_092;
  wire popcount30_rptt_core_093;
  wire popcount30_rptt_core_096;
  wire popcount30_rptt_core_098;
  wire popcount30_rptt_core_099;
  wire popcount30_rptt_core_101;
  wire popcount30_rptt_core_103;
  wire popcount30_rptt_core_105;
  wire popcount30_rptt_core_109;
  wire popcount30_rptt_core_110;
  wire popcount30_rptt_core_111;
  wire popcount30_rptt_core_113;
  wire popcount30_rptt_core_114;
  wire popcount30_rptt_core_115;
  wire popcount30_rptt_core_116;
  wire popcount30_rptt_core_117;
  wire popcount30_rptt_core_118;
  wire popcount30_rptt_core_120;
  wire popcount30_rptt_core_121;
  wire popcount30_rptt_core_123;
  wire popcount30_rptt_core_124;
  wire popcount30_rptt_core_127;
  wire popcount30_rptt_core_129;
  wire popcount30_rptt_core_130;
  wire popcount30_rptt_core_132;
  wire popcount30_rptt_core_133;
  wire popcount30_rptt_core_134;
  wire popcount30_rptt_core_135;
  wire popcount30_rptt_core_136;
  wire popcount30_rptt_core_138_not;
  wire popcount30_rptt_core_139;
  wire popcount30_rptt_core_140;
  wire popcount30_rptt_core_141;
  wire popcount30_rptt_core_143;
  wire popcount30_rptt_core_147;
  wire popcount30_rptt_core_148;
  wire popcount30_rptt_core_149;
  wire popcount30_rptt_core_150;
  wire popcount30_rptt_core_151;
  wire popcount30_rptt_core_152;
  wire popcount30_rptt_core_153;
  wire popcount30_rptt_core_154;
  wire popcount30_rptt_core_155;
  wire popcount30_rptt_core_157;
  wire popcount30_rptt_core_159;
  wire popcount30_rptt_core_160;
  wire popcount30_rptt_core_161;
  wire popcount30_rptt_core_162;
  wire popcount30_rptt_core_163;
  wire popcount30_rptt_core_167;
  wire popcount30_rptt_core_168;
  wire popcount30_rptt_core_169;
  wire popcount30_rptt_core_170;
  wire popcount30_rptt_core_173;
  wire popcount30_rptt_core_176;
  wire popcount30_rptt_core_179;
  wire popcount30_rptt_core_180;
  wire popcount30_rptt_core_181;
  wire popcount30_rptt_core_182;
  wire popcount30_rptt_core_183_not;
  wire popcount30_rptt_core_186;
  wire popcount30_rptt_core_187;
  wire popcount30_rptt_core_188;
  wire popcount30_rptt_core_189;
  wire popcount30_rptt_core_190;
  wire popcount30_rptt_core_191;
  wire popcount30_rptt_core_193;
  wire popcount30_rptt_core_197;
  wire popcount30_rptt_core_199;
  wire popcount30_rptt_core_201_not;
  wire popcount30_rptt_core_204;
  wire popcount30_rptt_core_206;
  wire popcount30_rptt_core_209;
  wire popcount30_rptt_core_211;
  wire popcount30_rptt_core_212;

  assign popcount30_rptt_core_032 = input_a[27] & input_a[24];
  assign popcount30_rptt_core_034 = ~(input_a[4] ^ input_a[16]);
  assign popcount30_rptt_core_035 = input_a[7] & input_a[5];
  assign popcount30_rptt_core_036 = ~(input_a[24] ^ input_a[9]);
  assign popcount30_rptt_core_037 = ~(input_a[15] | input_a[26]);
  assign popcount30_rptt_core_038 = input_a[24] ^ input_a[13];
  assign popcount30_rptt_core_039 = input_a[27] ^ input_a[10];
  assign popcount30_rptt_core_041 = input_a[27] | input_a[8];
  assign popcount30_rptt_core_043_not = ~input_a[5];
  assign popcount30_rptt_core_044 = input_a[25] & input_a[14];
  assign popcount30_rptt_core_046 = ~(input_a[24] | input_a[29]);
  assign popcount30_rptt_core_047 = ~(input_a[18] | input_a[23]);
  assign popcount30_rptt_core_052 = input_a[15] | input_a[10];
  assign popcount30_rptt_core_053 = input_a[8] | input_a[3];
  assign popcount30_rptt_core_054 = ~input_a[16];
  assign popcount30_rptt_core_055 = input_a[3] ^ input_a[16];
  assign popcount30_rptt_core_057_not = ~input_a[1];
  assign popcount30_rptt_core_060 = ~(input_a[18] & input_a[2]);
  assign popcount30_rptt_core_062 = input_a[24] ^ input_a[7];
  assign popcount30_rptt_core_064 = input_a[18] ^ input_a[2];
  assign popcount30_rptt_core_065 = input_a[21] & input_a[26];
  assign popcount30_rptt_core_068 = ~input_a[11];
  assign popcount30_rptt_core_069 = ~(input_a[14] ^ input_a[17]);
  assign popcount30_rptt_core_071 = ~(input_a[6] & input_a[15]);
  assign popcount30_rptt_core_072 = ~input_a[17];
  assign popcount30_rptt_core_073 = input_a[7] ^ input_a[11];
  assign popcount30_rptt_core_074 = input_a[18] | input_a[22];
  assign popcount30_rptt_core_076 = input_a[14] ^ input_a[21];
  assign popcount30_rptt_core_078 = ~input_a[12];
  assign popcount30_rptt_core_079 = ~(input_a[7] ^ input_a[0]);
  assign popcount30_rptt_core_080 = ~(input_a[4] ^ input_a[1]);
  assign popcount30_rptt_core_081 = ~(input_a[12] & input_a[1]);
  assign popcount30_rptt_core_083 = ~(input_a[28] ^ input_a[25]);
  assign popcount30_rptt_core_084 = ~(input_a[18] & input_a[19]);
  assign popcount30_rptt_core_085_not = ~input_a[17];
  assign popcount30_rptt_core_087 = input_a[27] | input_a[0];
  assign popcount30_rptt_core_088 = ~input_a[6];
  assign popcount30_rptt_core_090 = input_a[21] & input_a[2];
  assign popcount30_rptt_core_092 = input_a[5] ^ input_a[27];
  assign popcount30_rptt_core_093 = ~(input_a[1] ^ input_a[12]);
  assign popcount30_rptt_core_096 = ~(input_a[14] | input_a[26]);
  assign popcount30_rptt_core_098 = input_a[26] ^ input_a[18];
  assign popcount30_rptt_core_099 = ~input_a[23];
  assign popcount30_rptt_core_101 = ~input_a[19];
  assign popcount30_rptt_core_103 = ~input_a[26];
  assign popcount30_rptt_core_105 = input_a[20] & input_a[20];
  assign popcount30_rptt_core_109 = ~(input_a[18] & input_a[6]);
  assign popcount30_rptt_core_110 = ~(input_a[9] | input_a[17]);
  assign popcount30_rptt_core_111 = ~(input_a[7] ^ input_a[3]);
  assign popcount30_rptt_core_113 = ~input_a[18];
  assign popcount30_rptt_core_114 = input_a[17] & input_a[5];
  assign popcount30_rptt_core_115 = ~(input_a[14] & input_a[21]);
  assign popcount30_rptt_core_116 = ~(input_a[13] | input_a[27]);
  assign popcount30_rptt_core_117 = ~(input_a[19] & input_a[9]);
  assign popcount30_rptt_core_118 = input_a[11] & input_a[16];
  assign popcount30_rptt_core_120 = ~(input_a[3] ^ input_a[2]);
  assign popcount30_rptt_core_121 = input_a[6] ^ input_a[12];
  assign popcount30_rptt_core_123 = input_a[5] ^ input_a[23];
  assign popcount30_rptt_core_124 = input_a[15] ^ input_a[8];
  assign popcount30_rptt_core_127 = ~input_a[8];
  assign popcount30_rptt_core_129 = ~(input_a[18] ^ input_a[7]);
  assign popcount30_rptt_core_130 = input_a[1] | input_a[15];
  assign popcount30_rptt_core_132 = input_a[9] | input_a[1];
  assign popcount30_rptt_core_133 = input_a[25] | input_a[14];
  assign popcount30_rptt_core_134 = input_a[22] & input_a[3];
  assign popcount30_rptt_core_135 = ~input_a[3];
  assign popcount30_rptt_core_136 = ~input_a[11];
  assign popcount30_rptt_core_138_not = ~input_a[9];
  assign popcount30_rptt_core_139 = input_a[5] | input_a[17];
  assign popcount30_rptt_core_140 = ~input_a[25];
  assign popcount30_rptt_core_141 = input_a[4] | input_a[3];
  assign popcount30_rptt_core_143 = ~(input_a[2] | input_a[5]);
  assign popcount30_rptt_core_147 = ~input_a[1];
  assign popcount30_rptt_core_148 = ~(input_a[16] | input_a[25]);
  assign popcount30_rptt_core_149 = input_a[11] ^ input_a[16];
  assign popcount30_rptt_core_150 = ~(input_a[0] & input_a[26]);
  assign popcount30_rptt_core_151 = ~(input_a[2] & input_a[1]);
  assign popcount30_rptt_core_152 = input_a[24] & input_a[25];
  assign popcount30_rptt_core_153 = ~(input_a[7] | input_a[4]);
  assign popcount30_rptt_core_154 = input_a[13] | input_a[16];
  assign popcount30_rptt_core_155 = ~(input_a[21] | input_a[2]);
  assign popcount30_rptt_core_157 = ~(input_a[25] ^ input_a[19]);
  assign popcount30_rptt_core_159 = input_a[20] | input_a[16];
  assign popcount30_rptt_core_160 = input_a[10] & input_a[22];
  assign popcount30_rptt_core_161 = ~(input_a[9] & input_a[27]);
  assign popcount30_rptt_core_162 = input_a[18] & input_a[25];
  assign popcount30_rptt_core_163 = input_a[1] & input_a[9];
  assign popcount30_rptt_core_167 = ~(input_a[11] & input_a[11]);
  assign popcount30_rptt_core_168 = ~input_a[17];
  assign popcount30_rptt_core_169 = ~(input_a[17] & input_a[0]);
  assign popcount30_rptt_core_170 = ~(input_a[9] | input_a[22]);
  assign popcount30_rptt_core_173 = ~(input_a[26] ^ input_a[28]);
  assign popcount30_rptt_core_176 = input_a[29] ^ input_a[20];
  assign popcount30_rptt_core_179 = input_a[14] ^ input_a[17];
  assign popcount30_rptt_core_180 = ~(input_a[22] | input_a[24]);
  assign popcount30_rptt_core_181 = input_a[9] & input_a[22];
  assign popcount30_rptt_core_182 = ~input_a[26];
  assign popcount30_rptt_core_183_not = ~input_a[6];
  assign popcount30_rptt_core_186 = ~(input_a[19] ^ input_a[8]);
  assign popcount30_rptt_core_187 = input_a[25] & input_a[17];
  assign popcount30_rptt_core_188 = ~input_a[8];
  assign popcount30_rptt_core_189 = ~(input_a[27] | input_a[1]);
  assign popcount30_rptt_core_190 = ~input_a[1];
  assign popcount30_rptt_core_191 = ~(input_a[13] | input_a[4]);
  assign popcount30_rptt_core_193 = input_a[29] & input_a[3];
  assign popcount30_rptt_core_197 = ~(input_a[13] & input_a[7]);
  assign popcount30_rptt_core_199 = input_a[16] ^ input_a[8];
  assign popcount30_rptt_core_201_not = ~input_a[29];
  assign popcount30_rptt_core_204 = input_a[21] ^ input_a[26];
  assign popcount30_rptt_core_206 = popcount30_rptt_core_204 ^ popcount30_rptt_core_182;
  assign popcount30_rptt_core_209 = ~input_a[3];
  assign popcount30_rptt_core_211 = input_a[17] & input_a[11];
  assign popcount30_rptt_core_212 = ~(input_a[8] ^ input_a[22]);

  assign popcount30_rptt_out[0] = 1'b0;
  assign popcount30_rptt_out[1] = popcount30_rptt_core_206;
  assign popcount30_rptt_out[2] = popcount30_rptt_core_206;
  assign popcount30_rptt_out[3] = popcount30_rptt_core_206;
  assign popcount30_rptt_out[4] = input_a[21];
endmodule