// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.899
// WCE=28.0
// EP=0.961536%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount29_di19(input [28:0] input_a, output [4:0] popcount29_di19_out);
  wire popcount29_di19_core_031;
  wire popcount29_di19_core_032;
  wire popcount29_di19_core_034;
  wire popcount29_di19_core_035;
  wire popcount29_di19_core_036;
  wire popcount29_di19_core_037;
  wire popcount29_di19_core_038;
  wire popcount29_di19_core_040;
  wire popcount29_di19_core_044_not;
  wire popcount29_di19_core_045;
  wire popcount29_di19_core_047;
  wire popcount29_di19_core_048;
  wire popcount29_di19_core_049_not;
  wire popcount29_di19_core_052;
  wire popcount29_di19_core_053;
  wire popcount29_di19_core_055;
  wire popcount29_di19_core_056;
  wire popcount29_di19_core_059;
  wire popcount29_di19_core_061;
  wire popcount29_di19_core_062;
  wire popcount29_di19_core_063;
  wire popcount29_di19_core_064;
  wire popcount29_di19_core_065;
  wire popcount29_di19_core_067;
  wire popcount29_di19_core_068;
  wire popcount29_di19_core_071;
  wire popcount29_di19_core_072;
  wire popcount29_di19_core_073;
  wire popcount29_di19_core_075;
  wire popcount29_di19_core_079;
  wire popcount29_di19_core_080;
  wire popcount29_di19_core_081;
  wire popcount29_di19_core_083;
  wire popcount29_di19_core_084;
  wire popcount29_di19_core_085;
  wire popcount29_di19_core_086;
  wire popcount29_di19_core_087;
  wire popcount29_di19_core_090;
  wire popcount29_di19_core_092;
  wire popcount29_di19_core_095;
  wire popcount29_di19_core_096;
  wire popcount29_di19_core_097;
  wire popcount29_di19_core_098;
  wire popcount29_di19_core_103;
  wire popcount29_di19_core_107;
  wire popcount29_di19_core_108;
  wire popcount29_di19_core_109;
  wire popcount29_di19_core_110;
  wire popcount29_di19_core_114;
  wire popcount29_di19_core_116;
  wire popcount29_di19_core_118;
  wire popcount29_di19_core_119;
  wire popcount29_di19_core_120;
  wire popcount29_di19_core_121;
  wire popcount29_di19_core_122;
  wire popcount29_di19_core_124;
  wire popcount29_di19_core_125;
  wire popcount29_di19_core_127;
  wire popcount29_di19_core_128;
  wire popcount29_di19_core_129;
  wire popcount29_di19_core_130;
  wire popcount29_di19_core_132;
  wire popcount29_di19_core_133;
  wire popcount29_di19_core_134;
  wire popcount29_di19_core_136;
  wire popcount29_di19_core_137;
  wire popcount29_di19_core_138;
  wire popcount29_di19_core_139;
  wire popcount29_di19_core_140;
  wire popcount29_di19_core_141;
  wire popcount29_di19_core_142;
  wire popcount29_di19_core_143;
  wire popcount29_di19_core_146;
  wire popcount29_di19_core_147;
  wire popcount29_di19_core_148;
  wire popcount29_di19_core_149;
  wire popcount29_di19_core_150;
  wire popcount29_di19_core_151;
  wire popcount29_di19_core_152;
  wire popcount29_di19_core_153;
  wire popcount29_di19_core_154;
  wire popcount29_di19_core_155;
  wire popcount29_di19_core_156;
  wire popcount29_di19_core_157;
  wire popcount29_di19_core_159;
  wire popcount29_di19_core_160;
  wire popcount29_di19_core_161;
  wire popcount29_di19_core_162;
  wire popcount29_di19_core_163;
  wire popcount29_di19_core_164;
  wire popcount29_di19_core_165;
  wire popcount29_di19_core_166;
  wire popcount29_di19_core_167;
  wire popcount29_di19_core_168;
  wire popcount29_di19_core_170;
  wire popcount29_di19_core_171;
  wire popcount29_di19_core_176;
  wire popcount29_di19_core_177;
  wire popcount29_di19_core_178;
  wire popcount29_di19_core_179;
  wire popcount29_di19_core_180;
  wire popcount29_di19_core_181;
  wire popcount29_di19_core_182_not;
  wire popcount29_di19_core_183;
  wire popcount29_di19_core_184;
  wire popcount29_di19_core_185;
  wire popcount29_di19_core_186;
  wire popcount29_di19_core_187;
  wire popcount29_di19_core_188;
  wire popcount29_di19_core_189;
  wire popcount29_di19_core_191;
  wire popcount29_di19_core_192;
  wire popcount29_di19_core_193;
  wire popcount29_di19_core_194;
  wire popcount29_di19_core_195;
  wire popcount29_di19_core_196;
  wire popcount29_di19_core_197;
  wire popcount29_di19_core_198;
  wire popcount29_di19_core_199;
  wire popcount29_di19_core_200;
  wire popcount29_di19_core_201;
  wire popcount29_di19_core_203;
  wire popcount29_di19_core_205;
  wire popcount29_di19_core_206;
  wire popcount29_di19_core_207;

  assign popcount29_di19_core_031 = input_a[28] ^ input_a[23];
  assign popcount29_di19_core_032 = ~(input_a[1] ^ input_a[23]);
  assign popcount29_di19_core_034 = ~(input_a[14] ^ input_a[19]);
  assign popcount29_di19_core_035 = ~(input_a[22] ^ input_a[17]);
  assign popcount29_di19_core_036 = ~(input_a[0] ^ input_a[18]);
  assign popcount29_di19_core_037 = ~input_a[23];
  assign popcount29_di19_core_038 = ~(input_a[27] | input_a[28]);
  assign popcount29_di19_core_040 = ~(input_a[18] | input_a[20]);
  assign popcount29_di19_core_044_not = ~input_a[17];
  assign popcount29_di19_core_045 = input_a[16] | input_a[27];
  assign popcount29_di19_core_047 = ~(input_a[24] & input_a[6]);
  assign popcount29_di19_core_048 = ~(input_a[23] | input_a[2]);
  assign popcount29_di19_core_049_not = ~input_a[14];
  assign popcount29_di19_core_052 = ~input_a[7];
  assign popcount29_di19_core_053 = input_a[7] & input_a[27];
  assign popcount29_di19_core_055 = ~input_a[2];
  assign popcount29_di19_core_056 = ~input_a[9];
  assign popcount29_di19_core_059 = ~(input_a[24] & input_a[15]);
  assign popcount29_di19_core_061 = ~(input_a[26] ^ input_a[13]);
  assign popcount29_di19_core_062 = input_a[0] | input_a[0];
  assign popcount29_di19_core_063 = ~input_a[7];
  assign popcount29_di19_core_064 = ~input_a[5];
  assign popcount29_di19_core_065 = ~input_a[15];
  assign popcount29_di19_core_067 = input_a[16] & input_a[22];
  assign popcount29_di19_core_068 = ~(input_a[5] ^ input_a[1]);
  assign popcount29_di19_core_071 = ~(input_a[22] | input_a[8]);
  assign popcount29_di19_core_072 = ~input_a[14];
  assign popcount29_di19_core_073 = ~(input_a[10] & input_a[6]);
  assign popcount29_di19_core_075 = input_a[12] ^ input_a[8];
  assign popcount29_di19_core_079 = ~(input_a[18] ^ input_a[13]);
  assign popcount29_di19_core_080 = ~input_a[23];
  assign popcount29_di19_core_081 = ~(input_a[28] | input_a[16]);
  assign popcount29_di19_core_083 = ~(input_a[20] ^ input_a[20]);
  assign popcount29_di19_core_084 = ~(input_a[14] & input_a[22]);
  assign popcount29_di19_core_085 = ~(input_a[20] & input_a[1]);
  assign popcount29_di19_core_086 = input_a[11] ^ input_a[27];
  assign popcount29_di19_core_087 = input_a[16] ^ input_a[16];
  assign popcount29_di19_core_090 = ~(input_a[13] ^ input_a[25]);
  assign popcount29_di19_core_092 = ~(input_a[14] ^ input_a[8]);
  assign popcount29_di19_core_095 = input_a[28] ^ input_a[14];
  assign popcount29_di19_core_096 = ~(input_a[13] ^ input_a[16]);
  assign popcount29_di19_core_097 = ~(input_a[17] & input_a[6]);
  assign popcount29_di19_core_098 = input_a[20] ^ input_a[2];
  assign popcount29_di19_core_103 = ~(input_a[24] ^ input_a[1]);
  assign popcount29_di19_core_107 = ~(input_a[0] & input_a[5]);
  assign popcount29_di19_core_108 = ~(input_a[5] & input_a[0]);
  assign popcount29_di19_core_109 = ~input_a[2];
  assign popcount29_di19_core_110 = input_a[23] | input_a[26];
  assign popcount29_di19_core_114 = input_a[1] ^ input_a[16];
  assign popcount29_di19_core_116 = ~(input_a[16] & input_a[28]);
  assign popcount29_di19_core_118 = ~(input_a[24] | input_a[3]);
  assign popcount29_di19_core_119 = ~input_a[11];
  assign popcount29_di19_core_120 = ~(input_a[15] | input_a[10]);
  assign popcount29_di19_core_121 = ~(input_a[26] ^ input_a[5]);
  assign popcount29_di19_core_122 = input_a[11] | input_a[11];
  assign popcount29_di19_core_124 = ~(input_a[7] & input_a[9]);
  assign popcount29_di19_core_125 = ~(input_a[12] & input_a[19]);
  assign popcount29_di19_core_127 = ~(input_a[7] & input_a[6]);
  assign popcount29_di19_core_128 = ~(input_a[6] & input_a[14]);
  assign popcount29_di19_core_129 = ~(input_a[6] & input_a[7]);
  assign popcount29_di19_core_130 = ~(input_a[26] ^ input_a[25]);
  assign popcount29_di19_core_132 = input_a[24] ^ input_a[9];
  assign popcount29_di19_core_133 = input_a[7] ^ input_a[21];
  assign popcount29_di19_core_134 = ~(input_a[9] & input_a[22]);
  assign popcount29_di19_core_136 = input_a[1] & input_a[2];
  assign popcount29_di19_core_137 = ~(input_a[6] | input_a[21]);
  assign popcount29_di19_core_138 = ~(input_a[24] ^ input_a[26]);
  assign popcount29_di19_core_139 = input_a[18] ^ input_a[1];
  assign popcount29_di19_core_140 = ~(input_a[16] | input_a[25]);
  assign popcount29_di19_core_141 = ~(input_a[12] & input_a[11]);
  assign popcount29_di19_core_142 = ~(input_a[0] ^ input_a[1]);
  assign popcount29_di19_core_143 = ~(input_a[21] | input_a[3]);
  assign popcount29_di19_core_146 = input_a[2] ^ input_a[0];
  assign popcount29_di19_core_147 = ~(input_a[5] & input_a[17]);
  assign popcount29_di19_core_148 = ~(input_a[14] ^ input_a[10]);
  assign popcount29_di19_core_149 = ~(input_a[1] | input_a[23]);
  assign popcount29_di19_core_150 = ~(input_a[3] ^ input_a[8]);
  assign popcount29_di19_core_151 = ~input_a[6];
  assign popcount29_di19_core_152 = ~input_a[21];
  assign popcount29_di19_core_153 = ~(input_a[10] | input_a[17]);
  assign popcount29_di19_core_154 = ~input_a[18];
  assign popcount29_di19_core_155 = input_a[20] & input_a[21];
  assign popcount29_di19_core_156 = ~(input_a[27] | input_a[8]);
  assign popcount29_di19_core_157 = input_a[8] & input_a[20];
  assign popcount29_di19_core_159 = ~input_a[6];
  assign popcount29_di19_core_160 = ~(input_a[2] & input_a[7]);
  assign popcount29_di19_core_161 = input_a[7] & input_a[8];
  assign popcount29_di19_core_162 = input_a[5] & input_a[0];
  assign popcount29_di19_core_163 = input_a[22] & input_a[0];
  assign popcount29_di19_core_164 = ~(input_a[5] | input_a[24]);
  assign popcount29_di19_core_165 = input_a[19] | input_a[0];
  assign popcount29_di19_core_166 = input_a[24] ^ input_a[14];
  assign popcount29_di19_core_167 = ~(input_a[17] | input_a[16]);
  assign popcount29_di19_core_168 = ~input_a[5];
  assign popcount29_di19_core_170 = input_a[14] ^ input_a[15];
  assign popcount29_di19_core_171 = ~(input_a[24] & input_a[12]);
  assign popcount29_di19_core_176 = input_a[23] & input_a[24];
  assign popcount29_di19_core_177 = ~input_a[19];
  assign popcount29_di19_core_178 = ~(input_a[15] ^ input_a[0]);
  assign popcount29_di19_core_179 = ~(input_a[5] ^ input_a[27]);
  assign popcount29_di19_core_180 = ~(input_a[23] ^ input_a[1]);
  assign popcount29_di19_core_181 = ~input_a[27];
  assign popcount29_di19_core_182_not = ~input_a[23];
  assign popcount29_di19_core_183 = ~(input_a[13] & input_a[21]);
  assign popcount29_di19_core_184 = ~input_a[10];
  assign popcount29_di19_core_185 = input_a[0] | input_a[22];
  assign popcount29_di19_core_186 = input_a[11] & input_a[26];
  assign popcount29_di19_core_187 = ~input_a[17];
  assign popcount29_di19_core_188 = ~(input_a[26] & input_a[21]);
  assign popcount29_di19_core_189 = ~(input_a[10] ^ input_a[18]);
  assign popcount29_di19_core_191 = ~input_a[24];
  assign popcount29_di19_core_192 = ~(input_a[20] & input_a[0]);
  assign popcount29_di19_core_193 = ~(input_a[10] ^ input_a[3]);
  assign popcount29_di19_core_194 = input_a[21] ^ input_a[27];
  assign popcount29_di19_core_195 = ~(input_a[11] & input_a[11]);
  assign popcount29_di19_core_196 = input_a[18] ^ input_a[12];
  assign popcount29_di19_core_197 = ~(input_a[28] ^ input_a[22]);
  assign popcount29_di19_core_198 = ~(input_a[10] | input_a[7]);
  assign popcount29_di19_core_199 = input_a[3] & input_a[18];
  assign popcount29_di19_core_200 = ~input_a[28];
  assign popcount29_di19_core_201 = ~(input_a[25] | input_a[1]);
  assign popcount29_di19_core_203 = input_a[24] ^ input_a[7];
  assign popcount29_di19_core_205 = input_a[21] ^ input_a[2];
  assign popcount29_di19_core_206 = ~(input_a[18] ^ input_a[12]);
  assign popcount29_di19_core_207 = input_a[20] & input_a[0];

  assign popcount29_di19_out[0] = 1'b0;
  assign popcount29_di19_out[1] = 1'b1;
  assign popcount29_di19_out[2] = 1'b1;
  assign popcount29_di19_out[3] = input_a[26];
  assign popcount29_di19_out[4] = input_a[28];
endmodule