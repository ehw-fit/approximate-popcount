// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.66295
// WCE=18.0
// EP=0.924139%
// Printed PDK parameters:
//  Area=16470774.0
//  Delay=40807444.0
//  Power=551060.0

module popcount36_kbjb(input [35:0] input_a, output [5:0] popcount36_kbjb_out);
  wire popcount36_kbjb_core_038;
  wire popcount36_kbjb_core_039;
  wire popcount36_kbjb_core_040;
  wire popcount36_kbjb_core_041;
  wire popcount36_kbjb_core_042;
  wire popcount36_kbjb_core_044;
  wire popcount36_kbjb_core_045;
  wire popcount36_kbjb_core_046;
  wire popcount36_kbjb_core_049;
  wire popcount36_kbjb_core_050;
  wire popcount36_kbjb_core_051;
  wire popcount36_kbjb_core_053;
  wire popcount36_kbjb_core_054;
  wire popcount36_kbjb_core_055;
  wire popcount36_kbjb_core_056;
  wire popcount36_kbjb_core_057;
  wire popcount36_kbjb_core_059;
  wire popcount36_kbjb_core_062;
  wire popcount36_kbjb_core_067;
  wire popcount36_kbjb_core_069;
  wire popcount36_kbjb_core_070;
  wire popcount36_kbjb_core_071;
  wire popcount36_kbjb_core_073;
  wire popcount36_kbjb_core_080;
  wire popcount36_kbjb_core_081;
  wire popcount36_kbjb_core_083;
  wire popcount36_kbjb_core_084;
  wire popcount36_kbjb_core_085;
  wire popcount36_kbjb_core_086;
  wire popcount36_kbjb_core_087;
  wire popcount36_kbjb_core_089;
  wire popcount36_kbjb_core_091;
  wire popcount36_kbjb_core_092;
  wire popcount36_kbjb_core_094;
  wire popcount36_kbjb_core_096;
  wire popcount36_kbjb_core_097;
  wire popcount36_kbjb_core_099;
  wire popcount36_kbjb_core_100;
  wire popcount36_kbjb_core_101;
  wire popcount36_kbjb_core_102;
  wire popcount36_kbjb_core_103;
  wire popcount36_kbjb_core_104;
  wire popcount36_kbjb_core_105_not;
  wire popcount36_kbjb_core_107;
  wire popcount36_kbjb_core_108;
  wire popcount36_kbjb_core_110;
  wire popcount36_kbjb_core_113;
  wire popcount36_kbjb_core_114;
  wire popcount36_kbjb_core_116;
  wire popcount36_kbjb_core_117;
  wire popcount36_kbjb_core_118;
  wire popcount36_kbjb_core_120;
  wire popcount36_kbjb_core_121;
  wire popcount36_kbjb_core_123;
  wire popcount36_kbjb_core_124_not;
  wire popcount36_kbjb_core_125;
  wire popcount36_kbjb_core_129;
  wire popcount36_kbjb_core_131;
  wire popcount36_kbjb_core_132;
  wire popcount36_kbjb_core_135;
  wire popcount36_kbjb_core_136;
  wire popcount36_kbjb_core_137;
  wire popcount36_kbjb_core_138;
  wire popcount36_kbjb_core_139;
  wire popcount36_kbjb_core_140;
  wire popcount36_kbjb_core_145;
  wire popcount36_kbjb_core_146;
  wire popcount36_kbjb_core_147;
  wire popcount36_kbjb_core_148;
  wire popcount36_kbjb_core_150;
  wire popcount36_kbjb_core_151;
  wire popcount36_kbjb_core_155;
  wire popcount36_kbjb_core_156;
  wire popcount36_kbjb_core_158;
  wire popcount36_kbjb_core_159;
  wire popcount36_kbjb_core_160;
  wire popcount36_kbjb_core_162;
  wire popcount36_kbjb_core_163;
  wire popcount36_kbjb_core_165;
  wire popcount36_kbjb_core_167;
  wire popcount36_kbjb_core_168;
  wire popcount36_kbjb_core_170;
  wire popcount36_kbjb_core_171;
  wire popcount36_kbjb_core_175;
  wire popcount36_kbjb_core_176;
  wire popcount36_kbjb_core_177;
  wire popcount36_kbjb_core_179;
  wire popcount36_kbjb_core_180;
  wire popcount36_kbjb_core_181;
  wire popcount36_kbjb_core_182;
  wire popcount36_kbjb_core_183;
  wire popcount36_kbjb_core_184;
  wire popcount36_kbjb_core_185;
  wire popcount36_kbjb_core_186;
  wire popcount36_kbjb_core_187;
  wire popcount36_kbjb_core_188;
  wire popcount36_kbjb_core_191;
  wire popcount36_kbjb_core_192;
  wire popcount36_kbjb_core_193;
  wire popcount36_kbjb_core_194;
  wire popcount36_kbjb_core_197;
  wire popcount36_kbjb_core_200;
  wire popcount36_kbjb_core_201;
  wire popcount36_kbjb_core_205;
  wire popcount36_kbjb_core_208;
  wire popcount36_kbjb_core_209;
  wire popcount36_kbjb_core_210;
  wire popcount36_kbjb_core_214;
  wire popcount36_kbjb_core_216;
  wire popcount36_kbjb_core_217;
  wire popcount36_kbjb_core_218;
  wire popcount36_kbjb_core_219;
  wire popcount36_kbjb_core_222;
  wire popcount36_kbjb_core_223;
  wire popcount36_kbjb_core_225;
  wire popcount36_kbjb_core_228;
  wire popcount36_kbjb_core_231;
  wire popcount36_kbjb_core_232;
  wire popcount36_kbjb_core_234;
  wire popcount36_kbjb_core_236;
  wire popcount36_kbjb_core_242;
  wire popcount36_kbjb_core_243;
  wire popcount36_kbjb_core_249;
  wire popcount36_kbjb_core_254;
  wire popcount36_kbjb_core_255;
  wire popcount36_kbjb_core_256;
  wire popcount36_kbjb_core_257;
  wire popcount36_kbjb_core_258;
  wire popcount36_kbjb_core_259_not;
  wire popcount36_kbjb_core_260;
  wire popcount36_kbjb_core_261;
  wire popcount36_kbjb_core_262;
  wire popcount36_kbjb_core_263;
  wire popcount36_kbjb_core_264;
  wire popcount36_kbjb_core_265;
  wire popcount36_kbjb_core_268;
  wire popcount36_kbjb_core_269;
  wire popcount36_kbjb_core_270;
  wire popcount36_kbjb_core_271;
  wire popcount36_kbjb_core_273;
  wire popcount36_kbjb_core_276;

  assign popcount36_kbjb_core_038 = ~(input_a[29] ^ input_a[10]);
  assign popcount36_kbjb_core_039 = ~input_a[26];
  assign popcount36_kbjb_core_040 = ~(input_a[1] | input_a[23]);
  assign popcount36_kbjb_core_041 = ~(input_a[4] | input_a[5]);
  assign popcount36_kbjb_core_042 = ~(input_a[16] & input_a[22]);
  assign popcount36_kbjb_core_044 = input_a[3] ^ input_a[32];
  assign popcount36_kbjb_core_045 = input_a[29] & input_a[8];
  assign popcount36_kbjb_core_046 = input_a[29] ^ input_a[14];
  assign popcount36_kbjb_core_049 = ~(input_a[2] ^ input_a[4]);
  assign popcount36_kbjb_core_050 = ~(input_a[12] | input_a[31]);
  assign popcount36_kbjb_core_051 = ~(input_a[25] ^ input_a[20]);
  assign popcount36_kbjb_core_053 = ~(input_a[32] ^ input_a[9]);
  assign popcount36_kbjb_core_054 = input_a[6] & input_a[25];
  assign popcount36_kbjb_core_055 = input_a[4] & input_a[28];
  assign popcount36_kbjb_core_056 = ~(input_a[25] ^ input_a[6]);
  assign popcount36_kbjb_core_057 = ~(input_a[20] ^ input_a[9]);
  assign popcount36_kbjb_core_059 = ~(input_a[25] | input_a[34]);
  assign popcount36_kbjb_core_062 = ~(input_a[34] & input_a[17]);
  assign popcount36_kbjb_core_067 = input_a[26] ^ input_a[7];
  assign popcount36_kbjb_core_069 = ~(input_a[28] & input_a[22]);
  assign popcount36_kbjb_core_070 = ~input_a[3];
  assign popcount36_kbjb_core_071 = ~input_a[4];
  assign popcount36_kbjb_core_073 = ~input_a[32];
  assign popcount36_kbjb_core_080 = ~input_a[23];
  assign popcount36_kbjb_core_081 = ~(input_a[29] & input_a[4]);
  assign popcount36_kbjb_core_083 = input_a[17] ^ input_a[31];
  assign popcount36_kbjb_core_084 = input_a[3] ^ input_a[9];
  assign popcount36_kbjb_core_085 = input_a[32] | input_a[30];
  assign popcount36_kbjb_core_086 = input_a[8] | input_a[34];
  assign popcount36_kbjb_core_087 = input_a[15] & input_a[33];
  assign popcount36_kbjb_core_089 = ~(input_a[29] ^ input_a[7]);
  assign popcount36_kbjb_core_091 = ~(input_a[32] | input_a[30]);
  assign popcount36_kbjb_core_092 = input_a[34] & input_a[17];
  assign popcount36_kbjb_core_094 = input_a[5] & input_a[16];
  assign popcount36_kbjb_core_096 = input_a[1] & input_a[35];
  assign popcount36_kbjb_core_097 = popcount36_kbjb_core_094 | popcount36_kbjb_core_096;
  assign popcount36_kbjb_core_099 = ~input_a[28];
  assign popcount36_kbjb_core_100 = input_a[13] & input_a[19];
  assign popcount36_kbjb_core_101 = popcount36_kbjb_core_092 | popcount36_kbjb_core_097;
  assign popcount36_kbjb_core_102 = ~(input_a[28] & input_a[15]);
  assign popcount36_kbjb_core_103 = popcount36_kbjb_core_101 | popcount36_kbjb_core_100;
  assign popcount36_kbjb_core_104 = input_a[28] & input_a[3];
  assign popcount36_kbjb_core_105_not = ~input_a[23];
  assign popcount36_kbjb_core_107 = input_a[33] & input_a[16];
  assign popcount36_kbjb_core_108 = ~(input_a[23] ^ input_a[22]);
  assign popcount36_kbjb_core_110 = input_a[32] | input_a[0];
  assign popcount36_kbjb_core_113 = input_a[10] & input_a[3];
  assign popcount36_kbjb_core_114 = popcount36_kbjb_core_103 | popcount36_kbjb_core_113;
  assign popcount36_kbjb_core_116 = input_a[5] & input_a[28];
  assign popcount36_kbjb_core_117 = popcount36_kbjb_core_087 | popcount36_kbjb_core_114;
  assign popcount36_kbjb_core_118 = input_a[2] | input_a[0];
  assign popcount36_kbjb_core_120 = ~(input_a[6] & input_a[20]);
  assign popcount36_kbjb_core_121 = ~(input_a[28] | input_a[12]);
  assign popcount36_kbjb_core_123 = ~(input_a[25] ^ input_a[11]);
  assign popcount36_kbjb_core_124_not = ~input_a[11];
  assign popcount36_kbjb_core_125 = ~(input_a[11] & input_a[24]);
  assign popcount36_kbjb_core_129 = ~(input_a[21] & input_a[8]);
  assign popcount36_kbjb_core_131 = input_a[34] ^ input_a[10];
  assign popcount36_kbjb_core_132 = ~(input_a[16] & input_a[28]);
  assign popcount36_kbjb_core_135 = ~input_a[21];
  assign popcount36_kbjb_core_136 = popcount36_kbjb_core_045 | popcount36_kbjb_core_117;
  assign popcount36_kbjb_core_137 = input_a[5] ^ input_a[34];
  assign popcount36_kbjb_core_138 = input_a[15] & input_a[18];
  assign popcount36_kbjb_core_139 = ~(input_a[20] ^ input_a[11]);
  assign popcount36_kbjb_core_140 = input_a[17] & input_a[10];
  assign popcount36_kbjb_core_145 = input_a[28] & input_a[4];
  assign popcount36_kbjb_core_146 = ~(input_a[21] | input_a[8]);
  assign popcount36_kbjb_core_147 = input_a[31] & input_a[0];
  assign popcount36_kbjb_core_148 = ~(input_a[1] & input_a[12]);
  assign popcount36_kbjb_core_150 = ~(input_a[33] ^ input_a[32]);
  assign popcount36_kbjb_core_151 = popcount36_kbjb_core_145 & popcount36_kbjb_core_147;
  assign popcount36_kbjb_core_155 = ~(input_a[23] & input_a[30]);
  assign popcount36_kbjb_core_156 = input_a[22] | input_a[3];
  assign popcount36_kbjb_core_158 = input_a[20] | input_a[0];
  assign popcount36_kbjb_core_159 = ~(input_a[32] & input_a[34]);
  assign popcount36_kbjb_core_160 = input_a[16] ^ input_a[30];
  assign popcount36_kbjb_core_162 = input_a[22] & input_a[11];
  assign popcount36_kbjb_core_163 = ~input_a[9];
  assign popcount36_kbjb_core_165 = input_a[27] & input_a[33];
  assign popcount36_kbjb_core_167 = input_a[12] ^ input_a[20];
  assign popcount36_kbjb_core_168 = input_a[12] & input_a[20];
  assign popcount36_kbjb_core_170 = popcount36_kbjb_core_162 ^ popcount36_kbjb_core_168;
  assign popcount36_kbjb_core_171 = popcount36_kbjb_core_162 & popcount36_kbjb_core_168;
  assign popcount36_kbjb_core_175 = input_a[7] & popcount36_kbjb_core_167;
  assign popcount36_kbjb_core_176 = ~(input_a[32] | input_a[21]);
  assign popcount36_kbjb_core_177 = ~(input_a[1] ^ input_a[31]);
  assign popcount36_kbjb_core_179 = popcount36_kbjb_core_151 ^ popcount36_kbjb_core_170;
  assign popcount36_kbjb_core_180 = popcount36_kbjb_core_151 & popcount36_kbjb_core_170;
  assign popcount36_kbjb_core_181 = popcount36_kbjb_core_179 ^ popcount36_kbjb_core_175;
  assign popcount36_kbjb_core_182 = popcount36_kbjb_core_179 & popcount36_kbjb_core_175;
  assign popcount36_kbjb_core_183 = popcount36_kbjb_core_180 | popcount36_kbjb_core_182;
  assign popcount36_kbjb_core_184 = popcount36_kbjb_core_171 | popcount36_kbjb_core_183;
  assign popcount36_kbjb_core_185 = ~(input_a[33] | input_a[32]);
  assign popcount36_kbjb_core_186 = ~input_a[31];
  assign popcount36_kbjb_core_187 = ~(input_a[29] | input_a[13]);
  assign popcount36_kbjb_core_188 = ~(input_a[19] | input_a[0]);
  assign popcount36_kbjb_core_191 = ~(input_a[2] & input_a[21]);
  assign popcount36_kbjb_core_192 = ~(input_a[12] & input_a[21]);
  assign popcount36_kbjb_core_193 = ~(input_a[4] | input_a[1]);
  assign popcount36_kbjb_core_194 = ~(input_a[7] & input_a[33]);
  assign popcount36_kbjb_core_197 = ~(input_a[12] & input_a[7]);
  assign popcount36_kbjb_core_200 = input_a[34] & input_a[25];
  assign popcount36_kbjb_core_201 = input_a[12] | input_a[8];
  assign popcount36_kbjb_core_205 = input_a[4] & input_a[1];
  assign popcount36_kbjb_core_208 = input_a[18] & input_a[27];
  assign popcount36_kbjb_core_209 = input_a[18] | input_a[9];
  assign popcount36_kbjb_core_210 = input_a[5] ^ input_a[5];
  assign popcount36_kbjb_core_214 = ~(input_a[34] ^ input_a[2]);
  assign popcount36_kbjb_core_216 = input_a[5] | input_a[16];
  assign popcount36_kbjb_core_217 = input_a[21] & input_a[25];
  assign popcount36_kbjb_core_218 = input_a[26] ^ input_a[31];
  assign popcount36_kbjb_core_219 = input_a[12] & input_a[34];
  assign popcount36_kbjb_core_222 = input_a[28] & input_a[16];
  assign popcount36_kbjb_core_223 = popcount36_kbjb_core_208 | popcount36_kbjb_core_217;
  assign popcount36_kbjb_core_225 = input_a[12] | input_a[11];
  assign popcount36_kbjb_core_228 = input_a[34] | input_a[9];
  assign popcount36_kbjb_core_231 = ~(input_a[1] ^ input_a[18]);
  assign popcount36_kbjb_core_232 = input_a[2] & input_a[14];
  assign popcount36_kbjb_core_234 = ~input_a[26];
  assign popcount36_kbjb_core_236 = popcount36_kbjb_core_181 & popcount36_kbjb_core_223;
  assign popcount36_kbjb_core_242 = popcount36_kbjb_core_184 ^ popcount36_kbjb_core_236;
  assign popcount36_kbjb_core_243 = popcount36_kbjb_core_184 & popcount36_kbjb_core_236;
  assign popcount36_kbjb_core_249 = ~input_a[1];
  assign popcount36_kbjb_core_254 = ~input_a[25];
  assign popcount36_kbjb_core_255 = input_a[14] & input_a[25];
  assign popcount36_kbjb_core_256 = ~input_a[13];
  assign popcount36_kbjb_core_257 = input_a[11] & input_a[4];
  assign popcount36_kbjb_core_258 = ~(input_a[10] | input_a[16]);
  assign popcount36_kbjb_core_259_not = ~input_a[17];
  assign popcount36_kbjb_core_260 = input_a[9] | input_a[34];
  assign popcount36_kbjb_core_261 = input_a[5] & input_a[16];
  assign popcount36_kbjb_core_262 = popcount36_kbjb_core_136 ^ popcount36_kbjb_core_242;
  assign popcount36_kbjb_core_263 = popcount36_kbjb_core_136 & popcount36_kbjb_core_242;
  assign popcount36_kbjb_core_264 = ~input_a[28];
  assign popcount36_kbjb_core_265 = ~(input_a[1] | input_a[32]);
  assign popcount36_kbjb_core_268 = input_a[10] & input_a[17];
  assign popcount36_kbjb_core_269 = popcount36_kbjb_core_243 | popcount36_kbjb_core_263;
  assign popcount36_kbjb_core_270 = input_a[25] ^ input_a[34];
  assign popcount36_kbjb_core_271 = ~input_a[7];
  assign popcount36_kbjb_core_273 = ~input_a[13];
  assign popcount36_kbjb_core_276 = ~(input_a[6] ^ input_a[4]);

  assign popcount36_kbjb_out[0] = input_a[6];
  assign popcount36_kbjb_out[1] = 1'b1;
  assign popcount36_kbjb_out[2] = 1'b1;
  assign popcount36_kbjb_out[3] = popcount36_kbjb_core_262;
  assign popcount36_kbjb_out[4] = popcount36_kbjb_core_269;
  assign popcount36_kbjb_out[5] = 1'b0;
endmodule