// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.58235
// WCE=26.0
// EP=0.974549%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_gyrw(input [31:0] input_a, output [5:0] popcount32_gyrw_out);
  wire popcount32_gyrw_core_035;
  wire popcount32_gyrw_core_036;
  wire popcount32_gyrw_core_037;
  wire popcount32_gyrw_core_039;
  wire popcount32_gyrw_core_041;
  wire popcount32_gyrw_core_042;
  wire popcount32_gyrw_core_043;
  wire popcount32_gyrw_core_044;
  wire popcount32_gyrw_core_045;
  wire popcount32_gyrw_core_047;
  wire popcount32_gyrw_core_048;
  wire popcount32_gyrw_core_049;
  wire popcount32_gyrw_core_050;
  wire popcount32_gyrw_core_051;
  wire popcount32_gyrw_core_055;
  wire popcount32_gyrw_core_056;
  wire popcount32_gyrw_core_057;
  wire popcount32_gyrw_core_058;
  wire popcount32_gyrw_core_059;
  wire popcount32_gyrw_core_060;
  wire popcount32_gyrw_core_064;
  wire popcount32_gyrw_core_065;
  wire popcount32_gyrw_core_069;
  wire popcount32_gyrw_core_070;
  wire popcount32_gyrw_core_072;
  wire popcount32_gyrw_core_074;
  wire popcount32_gyrw_core_075;
  wire popcount32_gyrw_core_077;
  wire popcount32_gyrw_core_079;
  wire popcount32_gyrw_core_081;
  wire popcount32_gyrw_core_082;
  wire popcount32_gyrw_core_084;
  wire popcount32_gyrw_core_085;
  wire popcount32_gyrw_core_086;
  wire popcount32_gyrw_core_087;
  wire popcount32_gyrw_core_088;
  wire popcount32_gyrw_core_089;
  wire popcount32_gyrw_core_090;
  wire popcount32_gyrw_core_092;
  wire popcount32_gyrw_core_093;
  wire popcount32_gyrw_core_097;
  wire popcount32_gyrw_core_098;
  wire popcount32_gyrw_core_099;
  wire popcount32_gyrw_core_100_not;
  wire popcount32_gyrw_core_103;
  wire popcount32_gyrw_core_104;
  wire popcount32_gyrw_core_105;
  wire popcount32_gyrw_core_106;
  wire popcount32_gyrw_core_107;
  wire popcount32_gyrw_core_112;
  wire popcount32_gyrw_core_114;
  wire popcount32_gyrw_core_116;
  wire popcount32_gyrw_core_117;
  wire popcount32_gyrw_core_118;
  wire popcount32_gyrw_core_120;
  wire popcount32_gyrw_core_121;
  wire popcount32_gyrw_core_124;
  wire popcount32_gyrw_core_125;
  wire popcount32_gyrw_core_126_not;
  wire popcount32_gyrw_core_127;
  wire popcount32_gyrw_core_128;
  wire popcount32_gyrw_core_130;
  wire popcount32_gyrw_core_134;
  wire popcount32_gyrw_core_136;
  wire popcount32_gyrw_core_137;
  wire popcount32_gyrw_core_138;
  wire popcount32_gyrw_core_141;
  wire popcount32_gyrw_core_142;
  wire popcount32_gyrw_core_146;
  wire popcount32_gyrw_core_147;
  wire popcount32_gyrw_core_148;
  wire popcount32_gyrw_core_149;
  wire popcount32_gyrw_core_150;
  wire popcount32_gyrw_core_151;
  wire popcount32_gyrw_core_152;
  wire popcount32_gyrw_core_153;
  wire popcount32_gyrw_core_154;
  wire popcount32_gyrw_core_158;
  wire popcount32_gyrw_core_159;
  wire popcount32_gyrw_core_161;
  wire popcount32_gyrw_core_162;
  wire popcount32_gyrw_core_163;
  wire popcount32_gyrw_core_164;
  wire popcount32_gyrw_core_165;
  wire popcount32_gyrw_core_167;
  wire popcount32_gyrw_core_171;
  wire popcount32_gyrw_core_172;
  wire popcount32_gyrw_core_175;
  wire popcount32_gyrw_core_176;
  wire popcount32_gyrw_core_177;
  wire popcount32_gyrw_core_178;
  wire popcount32_gyrw_core_179;
  wire popcount32_gyrw_core_180;
  wire popcount32_gyrw_core_181;
  wire popcount32_gyrw_core_184;
  wire popcount32_gyrw_core_185;
  wire popcount32_gyrw_core_187;
  wire popcount32_gyrw_core_189;
  wire popcount32_gyrw_core_190;
  wire popcount32_gyrw_core_192;
  wire popcount32_gyrw_core_193;
  wire popcount32_gyrw_core_195;
  wire popcount32_gyrw_core_196;
  wire popcount32_gyrw_core_197;
  wire popcount32_gyrw_core_198;
  wire popcount32_gyrw_core_203;
  wire popcount32_gyrw_core_204;
  wire popcount32_gyrw_core_205;
  wire popcount32_gyrw_core_209;
  wire popcount32_gyrw_core_210;
  wire popcount32_gyrw_core_214;
  wire popcount32_gyrw_core_215;
  wire popcount32_gyrw_core_217;
  wire popcount32_gyrw_core_218;
  wire popcount32_gyrw_core_220;
  wire popcount32_gyrw_core_221;
  wire popcount32_gyrw_core_222;
  wire popcount32_gyrw_core_223;
  wire popcount32_gyrw_core_224;
  wire popcount32_gyrw_core_225;

  assign popcount32_gyrw_core_035 = ~input_a[20];
  assign popcount32_gyrw_core_036 = input_a[19] ^ input_a[14];
  assign popcount32_gyrw_core_037 = input_a[29] | input_a[7];
  assign popcount32_gyrw_core_039 = ~(input_a[26] ^ input_a[10]);
  assign popcount32_gyrw_core_041 = ~input_a[11];
  assign popcount32_gyrw_core_042 = input_a[2] | input_a[18];
  assign popcount32_gyrw_core_043 = ~(input_a[29] & input_a[1]);
  assign popcount32_gyrw_core_044 = ~(input_a[20] | input_a[4]);
  assign popcount32_gyrw_core_045 = ~(input_a[9] ^ input_a[7]);
  assign popcount32_gyrw_core_047 = ~(input_a[14] & input_a[28]);
  assign popcount32_gyrw_core_048 = ~(input_a[9] & input_a[8]);
  assign popcount32_gyrw_core_049 = ~(input_a[30] | input_a[7]);
  assign popcount32_gyrw_core_050 = input_a[5] ^ input_a[29];
  assign popcount32_gyrw_core_051 = input_a[4] | input_a[28];
  assign popcount32_gyrw_core_055 = input_a[2] & input_a[18];
  assign popcount32_gyrw_core_056 = input_a[12] ^ input_a[23];
  assign popcount32_gyrw_core_057 = input_a[14] ^ input_a[13];
  assign popcount32_gyrw_core_058 = input_a[23] ^ input_a[15];
  assign popcount32_gyrw_core_059 = ~(input_a[4] & input_a[21]);
  assign popcount32_gyrw_core_060 = ~(input_a[13] ^ input_a[6]);
  assign popcount32_gyrw_core_064 = ~(input_a[6] & input_a[7]);
  assign popcount32_gyrw_core_065 = ~(input_a[10] | input_a[19]);
  assign popcount32_gyrw_core_069 = input_a[9] & input_a[8];
  assign popcount32_gyrw_core_070 = ~(input_a[16] & input_a[14]);
  assign popcount32_gyrw_core_072 = ~(input_a[3] ^ input_a[13]);
  assign popcount32_gyrw_core_074 = input_a[12] ^ input_a[4];
  assign popcount32_gyrw_core_075 = ~(input_a[22] | input_a[21]);
  assign popcount32_gyrw_core_077 = ~(input_a[12] | input_a[20]);
  assign popcount32_gyrw_core_079 = input_a[26] | input_a[22];
  assign popcount32_gyrw_core_081 = input_a[9] & input_a[16];
  assign popcount32_gyrw_core_082 = ~(input_a[9] | input_a[14]);
  assign popcount32_gyrw_core_084 = ~(input_a[30] & input_a[24]);
  assign popcount32_gyrw_core_085 = ~(input_a[20] | input_a[29]);
  assign popcount32_gyrw_core_086 = input_a[30] | input_a[5];
  assign popcount32_gyrw_core_087 = ~input_a[12];
  assign popcount32_gyrw_core_088 = input_a[6] ^ input_a[22];
  assign popcount32_gyrw_core_089 = input_a[12] & input_a[12];
  assign popcount32_gyrw_core_090 = input_a[24] | input_a[2];
  assign popcount32_gyrw_core_092 = input_a[24] ^ input_a[13];
  assign popcount32_gyrw_core_093 = ~input_a[3];
  assign popcount32_gyrw_core_097 = ~(input_a[19] | input_a[30]);
  assign popcount32_gyrw_core_098 = input_a[13] ^ input_a[1];
  assign popcount32_gyrw_core_099 = ~(input_a[17] ^ input_a[24]);
  assign popcount32_gyrw_core_100_not = ~input_a[8];
  assign popcount32_gyrw_core_103 = ~(input_a[2] ^ input_a[27]);
  assign popcount32_gyrw_core_104 = input_a[29] | input_a[28];
  assign popcount32_gyrw_core_105 = ~(input_a[16] | input_a[27]);
  assign popcount32_gyrw_core_106 = ~(input_a[27] & input_a[11]);
  assign popcount32_gyrw_core_107 = ~(input_a[25] & input_a[1]);
  assign popcount32_gyrw_core_112 = input_a[0] | input_a[18];
  assign popcount32_gyrw_core_114 = ~(input_a[4] & input_a[24]);
  assign popcount32_gyrw_core_116 = input_a[28] & input_a[25];
  assign popcount32_gyrw_core_117 = input_a[29] | input_a[19];
  assign popcount32_gyrw_core_118 = ~(input_a[23] | input_a[22]);
  assign popcount32_gyrw_core_120 = ~(input_a[0] | input_a[11]);
  assign popcount32_gyrw_core_121 = ~input_a[2];
  assign popcount32_gyrw_core_124 = input_a[6] & input_a[24];
  assign popcount32_gyrw_core_125 = ~(input_a[23] | input_a[23]);
  assign popcount32_gyrw_core_126_not = ~input_a[17];
  assign popcount32_gyrw_core_127 = ~(input_a[19] ^ input_a[12]);
  assign popcount32_gyrw_core_128 = ~(input_a[14] | input_a[14]);
  assign popcount32_gyrw_core_130 = input_a[13] ^ input_a[12];
  assign popcount32_gyrw_core_134 = input_a[27] & input_a[22];
  assign popcount32_gyrw_core_136 = input_a[26] | input_a[23];
  assign popcount32_gyrw_core_137 = ~(input_a[24] | input_a[4]);
  assign popcount32_gyrw_core_138 = ~(input_a[19] | input_a[18]);
  assign popcount32_gyrw_core_141 = input_a[10] ^ input_a[3];
  assign popcount32_gyrw_core_142 = input_a[15] | input_a[4];
  assign popcount32_gyrw_core_146 = input_a[23] | input_a[15];
  assign popcount32_gyrw_core_147 = input_a[3] | input_a[9];
  assign popcount32_gyrw_core_148 = ~(input_a[7] ^ input_a[1]);
  assign popcount32_gyrw_core_149 = ~(input_a[28] | input_a[25]);
  assign popcount32_gyrw_core_150 = ~input_a[21];
  assign popcount32_gyrw_core_151 = ~input_a[16];
  assign popcount32_gyrw_core_152 = ~(input_a[27] ^ input_a[30]);
  assign popcount32_gyrw_core_153 = ~(input_a[3] ^ input_a[8]);
  assign popcount32_gyrw_core_154 = input_a[28] ^ input_a[22];
  assign popcount32_gyrw_core_158 = ~(input_a[6] ^ input_a[26]);
  assign popcount32_gyrw_core_159 = input_a[16] & input_a[16];
  assign popcount32_gyrw_core_161 = input_a[0] ^ input_a[12];
  assign popcount32_gyrw_core_162 = ~input_a[8];
  assign popcount32_gyrw_core_163 = ~(input_a[0] & input_a[19]);
  assign popcount32_gyrw_core_164 = ~(input_a[10] & input_a[7]);
  assign popcount32_gyrw_core_165 = input_a[9] | input_a[19];
  assign popcount32_gyrw_core_167 = ~input_a[19];
  assign popcount32_gyrw_core_171 = ~(input_a[25] | input_a[28]);
  assign popcount32_gyrw_core_172 = ~(input_a[11] & input_a[26]);
  assign popcount32_gyrw_core_175 = input_a[8] | input_a[16];
  assign popcount32_gyrw_core_176 = input_a[25] | input_a[31];
  assign popcount32_gyrw_core_177 = input_a[28] | input_a[8];
  assign popcount32_gyrw_core_178 = ~(input_a[27] & input_a[29]);
  assign popcount32_gyrw_core_179 = ~(input_a[13] | input_a[27]);
  assign popcount32_gyrw_core_180 = ~(input_a[18] ^ input_a[29]);
  assign popcount32_gyrw_core_181 = input_a[3] & input_a[20];
  assign popcount32_gyrw_core_184 = input_a[16] | input_a[28];
  assign popcount32_gyrw_core_185 = input_a[25] ^ input_a[16];
  assign popcount32_gyrw_core_187 = ~(input_a[13] ^ input_a[26]);
  assign popcount32_gyrw_core_189 = ~(input_a[19] & input_a[29]);
  assign popcount32_gyrw_core_190 = ~(input_a[6] ^ input_a[0]);
  assign popcount32_gyrw_core_192 = input_a[19] & input_a[21];
  assign popcount32_gyrw_core_193 = ~input_a[1];
  assign popcount32_gyrw_core_195 = input_a[26] | input_a[22];
  assign popcount32_gyrw_core_196 = ~(input_a[14] ^ input_a[29]);
  assign popcount32_gyrw_core_197 = ~(input_a[30] ^ input_a[17]);
  assign popcount32_gyrw_core_198 = ~(input_a[14] | input_a[10]);
  assign popcount32_gyrw_core_203 = input_a[31] & input_a[10];
  assign popcount32_gyrw_core_204 = ~(input_a[9] | input_a[29]);
  assign popcount32_gyrw_core_205 = ~(input_a[18] & input_a[22]);
  assign popcount32_gyrw_core_209 = ~(input_a[11] | input_a[0]);
  assign popcount32_gyrw_core_210 = input_a[6] & input_a[13];
  assign popcount32_gyrw_core_214 = ~(input_a[14] ^ input_a[14]);
  assign popcount32_gyrw_core_215 = input_a[18] ^ input_a[1];
  assign popcount32_gyrw_core_217 = input_a[11] & input_a[16];
  assign popcount32_gyrw_core_218 = ~input_a[27];
  assign popcount32_gyrw_core_220 = ~input_a[8];
  assign popcount32_gyrw_core_221 = ~(input_a[15] & input_a[12]);
  assign popcount32_gyrw_core_222 = input_a[9] | input_a[20];
  assign popcount32_gyrw_core_223 = input_a[3] ^ input_a[5];
  assign popcount32_gyrw_core_224 = ~(input_a[2] | input_a[22]);
  assign popcount32_gyrw_core_225 = ~(input_a[13] ^ input_a[9]);

  assign popcount32_gyrw_out[0] = input_a[0];
  assign popcount32_gyrw_out[1] = 1'b0;
  assign popcount32_gyrw_out[2] = 1'b1;
  assign popcount32_gyrw_out[3] = input_a[18];
  assign popcount32_gyrw_out[4] = 1'b0;
  assign popcount32_gyrw_out[5] = 1'b0;
endmodule