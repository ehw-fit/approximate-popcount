// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=17.3797
// WCE=51.0
// EP=0.943353%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount38_1bs7(input [37:0] input_a, output [5:0] popcount38_1bs7_out);
  wire popcount38_1bs7_core_041;
  wire popcount38_1bs7_core_042;
  wire popcount38_1bs7_core_043;
  wire popcount38_1bs7_core_045;
  wire popcount38_1bs7_core_046;
  wire popcount38_1bs7_core_048;
  wire popcount38_1bs7_core_050;
  wire popcount38_1bs7_core_051;
  wire popcount38_1bs7_core_052;
  wire popcount38_1bs7_core_053;
  wire popcount38_1bs7_core_055;
  wire popcount38_1bs7_core_056;
  wire popcount38_1bs7_core_058;
  wire popcount38_1bs7_core_062;
  wire popcount38_1bs7_core_063;
  wire popcount38_1bs7_core_064;
  wire popcount38_1bs7_core_065;
  wire popcount38_1bs7_core_068;
  wire popcount38_1bs7_core_072;
  wire popcount38_1bs7_core_073_not;
  wire popcount38_1bs7_core_074;
  wire popcount38_1bs7_core_078;
  wire popcount38_1bs7_core_079;
  wire popcount38_1bs7_core_080;
  wire popcount38_1bs7_core_081;
  wire popcount38_1bs7_core_082;
  wire popcount38_1bs7_core_084;
  wire popcount38_1bs7_core_085;
  wire popcount38_1bs7_core_087;
  wire popcount38_1bs7_core_088;
  wire popcount38_1bs7_core_089;
  wire popcount38_1bs7_core_090;
  wire popcount38_1bs7_core_093;
  wire popcount38_1bs7_core_094;
  wire popcount38_1bs7_core_095;
  wire popcount38_1bs7_core_096;
  wire popcount38_1bs7_core_097;
  wire popcount38_1bs7_core_098;
  wire popcount38_1bs7_core_100;
  wire popcount38_1bs7_core_103;
  wire popcount38_1bs7_core_104;
  wire popcount38_1bs7_core_105;
  wire popcount38_1bs7_core_106;
  wire popcount38_1bs7_core_109;
  wire popcount38_1bs7_core_111;
  wire popcount38_1bs7_core_112;
  wire popcount38_1bs7_core_114_not;
  wire popcount38_1bs7_core_115;
  wire popcount38_1bs7_core_116;
  wire popcount38_1bs7_core_120;
  wire popcount38_1bs7_core_121;
  wire popcount38_1bs7_core_122;
  wire popcount38_1bs7_core_123;
  wire popcount38_1bs7_core_124;
  wire popcount38_1bs7_core_127;
  wire popcount38_1bs7_core_128;
  wire popcount38_1bs7_core_129;
  wire popcount38_1bs7_core_130;
  wire popcount38_1bs7_core_131;
  wire popcount38_1bs7_core_135;
  wire popcount38_1bs7_core_137;
  wire popcount38_1bs7_core_139;
  wire popcount38_1bs7_core_140;
  wire popcount38_1bs7_core_141;
  wire popcount38_1bs7_core_142;
  wire popcount38_1bs7_core_144;
  wire popcount38_1bs7_core_146;
  wire popcount38_1bs7_core_147;
  wire popcount38_1bs7_core_148;
  wire popcount38_1bs7_core_150;
  wire popcount38_1bs7_core_151;
  wire popcount38_1bs7_core_152;
  wire popcount38_1bs7_core_155;
  wire popcount38_1bs7_core_156;
  wire popcount38_1bs7_core_157;
  wire popcount38_1bs7_core_159;
  wire popcount38_1bs7_core_160;
  wire popcount38_1bs7_core_162;
  wire popcount38_1bs7_core_163;
  wire popcount38_1bs7_core_164;
  wire popcount38_1bs7_core_165;
  wire popcount38_1bs7_core_166;
  wire popcount38_1bs7_core_167;
  wire popcount38_1bs7_core_168;
  wire popcount38_1bs7_core_171;
  wire popcount38_1bs7_core_172;
  wire popcount38_1bs7_core_173;
  wire popcount38_1bs7_core_174;
  wire popcount38_1bs7_core_176;
  wire popcount38_1bs7_core_178;
  wire popcount38_1bs7_core_179;
  wire popcount38_1bs7_core_181;
  wire popcount38_1bs7_core_182;
  wire popcount38_1bs7_core_183;
  wire popcount38_1bs7_core_184;
  wire popcount38_1bs7_core_185;
  wire popcount38_1bs7_core_187_not;
  wire popcount38_1bs7_core_189;
  wire popcount38_1bs7_core_191;
  wire popcount38_1bs7_core_194;
  wire popcount38_1bs7_core_195;
  wire popcount38_1bs7_core_196;
  wire popcount38_1bs7_core_197;
  wire popcount38_1bs7_core_199;
  wire popcount38_1bs7_core_201;
  wire popcount38_1bs7_core_202;
  wire popcount38_1bs7_core_203;
  wire popcount38_1bs7_core_204;
  wire popcount38_1bs7_core_205;
  wire popcount38_1bs7_core_208;
  wire popcount38_1bs7_core_211;
  wire popcount38_1bs7_core_214;
  wire popcount38_1bs7_core_215;
  wire popcount38_1bs7_core_216;
  wire popcount38_1bs7_core_218;
  wire popcount38_1bs7_core_219;
  wire popcount38_1bs7_core_220;
  wire popcount38_1bs7_core_221;
  wire popcount38_1bs7_core_223;
  wire popcount38_1bs7_core_224;
  wire popcount38_1bs7_core_225;
  wire popcount38_1bs7_core_226;
  wire popcount38_1bs7_core_227;
  wire popcount38_1bs7_core_229;
  wire popcount38_1bs7_core_231;
  wire popcount38_1bs7_core_232;
  wire popcount38_1bs7_core_234;
  wire popcount38_1bs7_core_235;
  wire popcount38_1bs7_core_236;
  wire popcount38_1bs7_core_237;
  wire popcount38_1bs7_core_239;
  wire popcount38_1bs7_core_242;
  wire popcount38_1bs7_core_243;
  wire popcount38_1bs7_core_244;
  wire popcount38_1bs7_core_247;
  wire popcount38_1bs7_core_248;
  wire popcount38_1bs7_core_249;
  wire popcount38_1bs7_core_251;
  wire popcount38_1bs7_core_254;
  wire popcount38_1bs7_core_257;
  wire popcount38_1bs7_core_258;
  wire popcount38_1bs7_core_260;
  wire popcount38_1bs7_core_261_not;
  wire popcount38_1bs7_core_262;
  wire popcount38_1bs7_core_264;
  wire popcount38_1bs7_core_265;
  wire popcount38_1bs7_core_267;
  wire popcount38_1bs7_core_268;
  wire popcount38_1bs7_core_269;
  wire popcount38_1bs7_core_270;
  wire popcount38_1bs7_core_272;
  wire popcount38_1bs7_core_273;
  wire popcount38_1bs7_core_274;
  wire popcount38_1bs7_core_275;
  wire popcount38_1bs7_core_276;
  wire popcount38_1bs7_core_277;
  wire popcount38_1bs7_core_280;
  wire popcount38_1bs7_core_282;
  wire popcount38_1bs7_core_285;
  wire popcount38_1bs7_core_286;
  wire popcount38_1bs7_core_287;
  wire popcount38_1bs7_core_289;
  wire popcount38_1bs7_core_290;
  wire popcount38_1bs7_core_292;
  wire popcount38_1bs7_core_293;
  wire popcount38_1bs7_core_295;

  assign popcount38_1bs7_core_041 = input_a[4] & input_a[1];
  assign popcount38_1bs7_core_042 = input_a[11] & input_a[8];
  assign popcount38_1bs7_core_043 = ~(input_a[29] & input_a[17]);
  assign popcount38_1bs7_core_045 = ~(input_a[11] ^ input_a[9]);
  assign popcount38_1bs7_core_046 = ~(input_a[0] & input_a[28]);
  assign popcount38_1bs7_core_048 = ~(input_a[2] ^ input_a[23]);
  assign popcount38_1bs7_core_050 = ~input_a[9];
  assign popcount38_1bs7_core_051 = ~(input_a[4] & input_a[37]);
  assign popcount38_1bs7_core_052 = input_a[17] ^ input_a[1];
  assign popcount38_1bs7_core_053 = input_a[20] & input_a[26];
  assign popcount38_1bs7_core_055 = ~(input_a[4] | input_a[24]);
  assign popcount38_1bs7_core_056 = ~(input_a[13] | input_a[16]);
  assign popcount38_1bs7_core_058 = ~(input_a[30] | input_a[37]);
  assign popcount38_1bs7_core_062 = input_a[2] & input_a[5];
  assign popcount38_1bs7_core_063 = ~(input_a[7] & input_a[23]);
  assign popcount38_1bs7_core_064 = ~(input_a[19] | input_a[36]);
  assign popcount38_1bs7_core_065 = ~(input_a[8] & input_a[30]);
  assign popcount38_1bs7_core_068 = input_a[3] ^ input_a[31];
  assign popcount38_1bs7_core_072 = ~(input_a[24] ^ input_a[27]);
  assign popcount38_1bs7_core_073_not = ~input_a[27];
  assign popcount38_1bs7_core_074 = ~(input_a[7] | input_a[1]);
  assign popcount38_1bs7_core_078 = ~input_a[32];
  assign popcount38_1bs7_core_079 = input_a[27] & input_a[33];
  assign popcount38_1bs7_core_080 = ~(input_a[15] ^ input_a[11]);
  assign popcount38_1bs7_core_081 = ~(input_a[2] | input_a[8]);
  assign popcount38_1bs7_core_082 = input_a[14] & input_a[28];
  assign popcount38_1bs7_core_084 = ~input_a[2];
  assign popcount38_1bs7_core_085 = input_a[28] & input_a[11];
  assign popcount38_1bs7_core_087 = ~(input_a[28] & input_a[22]);
  assign popcount38_1bs7_core_088 = input_a[13] & input_a[37];
  assign popcount38_1bs7_core_089 = input_a[35] & input_a[14];
  assign popcount38_1bs7_core_090 = ~input_a[30];
  assign popcount38_1bs7_core_093 = input_a[26] ^ input_a[33];
  assign popcount38_1bs7_core_094 = input_a[17] & input_a[17];
  assign popcount38_1bs7_core_095 = input_a[22] | input_a[1];
  assign popcount38_1bs7_core_096 = ~(input_a[10] & input_a[28]);
  assign popcount38_1bs7_core_097 = input_a[34] & input_a[18];
  assign popcount38_1bs7_core_098 = input_a[16] ^ input_a[3];
  assign popcount38_1bs7_core_100 = ~(input_a[35] & input_a[33]);
  assign popcount38_1bs7_core_103 = input_a[2] | input_a[30];
  assign popcount38_1bs7_core_104 = ~(input_a[1] & input_a[31]);
  assign popcount38_1bs7_core_105 = ~input_a[21];
  assign popcount38_1bs7_core_106 = ~(input_a[13] | input_a[12]);
  assign popcount38_1bs7_core_109 = input_a[24] | input_a[3];
  assign popcount38_1bs7_core_111 = ~(input_a[23] & input_a[8]);
  assign popcount38_1bs7_core_112 = input_a[9] & input_a[1];
  assign popcount38_1bs7_core_114_not = ~input_a[0];
  assign popcount38_1bs7_core_115 = ~(input_a[1] & input_a[18]);
  assign popcount38_1bs7_core_116 = input_a[25] | input_a[21];
  assign popcount38_1bs7_core_120 = ~(input_a[24] | input_a[26]);
  assign popcount38_1bs7_core_121 = input_a[30] | input_a[33];
  assign popcount38_1bs7_core_122 = ~(input_a[6] & input_a[4]);
  assign popcount38_1bs7_core_123 = ~(input_a[12] & input_a[23]);
  assign popcount38_1bs7_core_124 = input_a[10] ^ input_a[3];
  assign popcount38_1bs7_core_127 = input_a[23] & input_a[7];
  assign popcount38_1bs7_core_128 = input_a[9] | input_a[17];
  assign popcount38_1bs7_core_129 = input_a[31] & input_a[29];
  assign popcount38_1bs7_core_130 = ~(input_a[0] & input_a[9]);
  assign popcount38_1bs7_core_131 = ~(input_a[23] ^ input_a[28]);
  assign popcount38_1bs7_core_135 = ~(input_a[11] & input_a[10]);
  assign popcount38_1bs7_core_137 = ~(input_a[18] | input_a[34]);
  assign popcount38_1bs7_core_139 = input_a[4] | input_a[1];
  assign popcount38_1bs7_core_140 = input_a[25] ^ input_a[25];
  assign popcount38_1bs7_core_141 = ~(input_a[30] & input_a[7]);
  assign popcount38_1bs7_core_142 = ~(input_a[27] & input_a[27]);
  assign popcount38_1bs7_core_144 = ~(input_a[32] | input_a[13]);
  assign popcount38_1bs7_core_146 = ~(input_a[7] | input_a[22]);
  assign popcount38_1bs7_core_147 = ~(input_a[8] | input_a[10]);
  assign popcount38_1bs7_core_148 = input_a[5] ^ input_a[19];
  assign popcount38_1bs7_core_150 = ~(input_a[3] | input_a[16]);
  assign popcount38_1bs7_core_151 = ~(input_a[15] | input_a[13]);
  assign popcount38_1bs7_core_152 = input_a[14] & input_a[11];
  assign popcount38_1bs7_core_155 = ~(input_a[23] | input_a[24]);
  assign popcount38_1bs7_core_156 = input_a[16] ^ input_a[12];
  assign popcount38_1bs7_core_157 = input_a[10] | input_a[10];
  assign popcount38_1bs7_core_159 = ~(input_a[33] ^ input_a[27]);
  assign popcount38_1bs7_core_160 = input_a[16] & input_a[1];
  assign popcount38_1bs7_core_162 = input_a[5] | input_a[15];
  assign popcount38_1bs7_core_163 = ~input_a[22];
  assign popcount38_1bs7_core_164 = input_a[11] ^ input_a[34];
  assign popcount38_1bs7_core_165 = input_a[31] | input_a[17];
  assign popcount38_1bs7_core_166 = input_a[21] ^ input_a[7];
  assign popcount38_1bs7_core_167 = input_a[23] ^ input_a[22];
  assign popcount38_1bs7_core_168 = input_a[14] | input_a[26];
  assign popcount38_1bs7_core_171 = input_a[10] | input_a[32];
  assign popcount38_1bs7_core_172 = input_a[0] | input_a[16];
  assign popcount38_1bs7_core_173 = ~(input_a[5] | input_a[35]);
  assign popcount38_1bs7_core_174 = ~input_a[15];
  assign popcount38_1bs7_core_176 = input_a[9] & input_a[24];
  assign popcount38_1bs7_core_178 = input_a[36] ^ input_a[18];
  assign popcount38_1bs7_core_179 = input_a[22] | input_a[23];
  assign popcount38_1bs7_core_181 = input_a[9] ^ input_a[11];
  assign popcount38_1bs7_core_182 = input_a[5] | input_a[29];
  assign popcount38_1bs7_core_183 = ~input_a[33];
  assign popcount38_1bs7_core_184 = input_a[37] & input_a[12];
  assign popcount38_1bs7_core_185 = input_a[35] ^ input_a[25];
  assign popcount38_1bs7_core_187_not = ~input_a[16];
  assign popcount38_1bs7_core_189 = ~input_a[4];
  assign popcount38_1bs7_core_191 = ~input_a[4];
  assign popcount38_1bs7_core_194 = ~(input_a[29] & input_a[3]);
  assign popcount38_1bs7_core_195 = ~(input_a[27] | input_a[9]);
  assign popcount38_1bs7_core_196 = input_a[2] | input_a[9];
  assign popcount38_1bs7_core_197 = input_a[0] & input_a[25];
  assign popcount38_1bs7_core_199 = input_a[6] & input_a[11];
  assign popcount38_1bs7_core_201 = ~(input_a[19] & input_a[31]);
  assign popcount38_1bs7_core_202 = input_a[34] ^ input_a[26];
  assign popcount38_1bs7_core_203 = ~(input_a[25] ^ input_a[34]);
  assign popcount38_1bs7_core_204 = ~input_a[29];
  assign popcount38_1bs7_core_205 = input_a[26] & input_a[11];
  assign popcount38_1bs7_core_208 = input_a[32] | input_a[31];
  assign popcount38_1bs7_core_211 = input_a[36] ^ input_a[28];
  assign popcount38_1bs7_core_214 = input_a[33] & input_a[33];
  assign popcount38_1bs7_core_215 = input_a[35] | input_a[7];
  assign popcount38_1bs7_core_216 = input_a[11] ^ input_a[17];
  assign popcount38_1bs7_core_218 = input_a[10] & input_a[12];
  assign popcount38_1bs7_core_219 = ~(input_a[30] | input_a[8]);
  assign popcount38_1bs7_core_220 = input_a[32] ^ input_a[36];
  assign popcount38_1bs7_core_221 = ~(input_a[7] & input_a[8]);
  assign popcount38_1bs7_core_223 = ~(input_a[2] | input_a[12]);
  assign popcount38_1bs7_core_224 = input_a[21] ^ input_a[28];
  assign popcount38_1bs7_core_225 = input_a[22] & input_a[19];
  assign popcount38_1bs7_core_226 = input_a[36] & input_a[22];
  assign popcount38_1bs7_core_227 = input_a[33] & input_a[21];
  assign popcount38_1bs7_core_229 = ~(input_a[21] | input_a[16]);
  assign popcount38_1bs7_core_231 = input_a[23] & input_a[36];
  assign popcount38_1bs7_core_232 = input_a[34] ^ input_a[28];
  assign popcount38_1bs7_core_234 = ~input_a[7];
  assign popcount38_1bs7_core_235 = input_a[10] & input_a[26];
  assign popcount38_1bs7_core_236 = input_a[7] & input_a[17];
  assign popcount38_1bs7_core_237 = ~(input_a[30] & input_a[35]);
  assign popcount38_1bs7_core_239 = input_a[37] | input_a[17];
  assign popcount38_1bs7_core_242 = input_a[0] | input_a[20];
  assign popcount38_1bs7_core_243 = ~(input_a[2] & input_a[20]);
  assign popcount38_1bs7_core_244 = ~input_a[24];
  assign popcount38_1bs7_core_247 = ~input_a[36];
  assign popcount38_1bs7_core_248 = ~(input_a[11] & input_a[35]);
  assign popcount38_1bs7_core_249 = ~input_a[5];
  assign popcount38_1bs7_core_251 = ~(input_a[33] & input_a[36]);
  assign popcount38_1bs7_core_254 = input_a[37] | input_a[7];
  assign popcount38_1bs7_core_257 = input_a[37] & input_a[11];
  assign popcount38_1bs7_core_258 = input_a[30] ^ input_a[32];
  assign popcount38_1bs7_core_260 = ~input_a[27];
  assign popcount38_1bs7_core_261_not = ~input_a[31];
  assign popcount38_1bs7_core_262 = input_a[9] & input_a[11];
  assign popcount38_1bs7_core_264 = ~(input_a[8] & input_a[32]);
  assign popcount38_1bs7_core_265 = input_a[4] | input_a[1];
  assign popcount38_1bs7_core_267 = input_a[5] & input_a[23];
  assign popcount38_1bs7_core_268 = ~(input_a[28] ^ input_a[5]);
  assign popcount38_1bs7_core_269 = ~input_a[6];
  assign popcount38_1bs7_core_270 = input_a[11] ^ input_a[1];
  assign popcount38_1bs7_core_272 = ~input_a[7];
  assign popcount38_1bs7_core_273 = ~(input_a[33] | input_a[28]);
  assign popcount38_1bs7_core_274 = input_a[17] & input_a[4];
  assign popcount38_1bs7_core_275 = ~(input_a[35] ^ input_a[5]);
  assign popcount38_1bs7_core_276 = ~(input_a[27] & input_a[18]);
  assign popcount38_1bs7_core_277 = ~(input_a[15] & input_a[2]);
  assign popcount38_1bs7_core_280 = ~input_a[9];
  assign popcount38_1bs7_core_282 = input_a[22] ^ input_a[0];
  assign popcount38_1bs7_core_285 = input_a[30] & input_a[14];
  assign popcount38_1bs7_core_286 = input_a[12] & input_a[3];
  assign popcount38_1bs7_core_287 = input_a[21] ^ input_a[28];
  assign popcount38_1bs7_core_289 = input_a[21] ^ input_a[33];
  assign popcount38_1bs7_core_290 = ~(input_a[6] & input_a[3]);
  assign popcount38_1bs7_core_292 = input_a[33] & input_a[0];
  assign popcount38_1bs7_core_293 = ~(input_a[7] & input_a[22]);
  assign popcount38_1bs7_core_295 = input_a[33] | input_a[29];

  assign popcount38_1bs7_out[0] = input_a[17];
  assign popcount38_1bs7_out[1] = input_a[27];
  assign popcount38_1bs7_out[2] = input_a[20];
  assign popcount38_1bs7_out[3] = 1'b0;
  assign popcount38_1bs7_out[4] = 1'b1;
  assign popcount38_1bs7_out[5] = input_a[0];
endmodule