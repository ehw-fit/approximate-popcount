// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.05348
// WCE=20.0
// EP=0.89872%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount35_19t3(input [34:0] input_a, output [5:0] popcount35_19t3_out);
  wire popcount35_19t3_core_037;
  wire popcount35_19t3_core_038;
  wire popcount35_19t3_core_039;
  wire popcount35_19t3_core_040;
  wire popcount35_19t3_core_041;
  wire popcount35_19t3_core_042;
  wire popcount35_19t3_core_043_not;
  wire popcount35_19t3_core_044;
  wire popcount35_19t3_core_047;
  wire popcount35_19t3_core_049;
  wire popcount35_19t3_core_050;
  wire popcount35_19t3_core_051;
  wire popcount35_19t3_core_052;
  wire popcount35_19t3_core_055;
  wire popcount35_19t3_core_057;
  wire popcount35_19t3_core_060;
  wire popcount35_19t3_core_061;
  wire popcount35_19t3_core_065;
  wire popcount35_19t3_core_066;
  wire popcount35_19t3_core_067;
  wire popcount35_19t3_core_069;
  wire popcount35_19t3_core_070;
  wire popcount35_19t3_core_071;
  wire popcount35_19t3_core_073;
  wire popcount35_19t3_core_074_not;
  wire popcount35_19t3_core_075;
  wire popcount35_19t3_core_076;
  wire popcount35_19t3_core_077;
  wire popcount35_19t3_core_079;
  wire popcount35_19t3_core_082;
  wire popcount35_19t3_core_083;
  wire popcount35_19t3_core_085;
  wire popcount35_19t3_core_089;
  wire popcount35_19t3_core_090;
  wire popcount35_19t3_core_091;
  wire popcount35_19t3_core_093;
  wire popcount35_19t3_core_094;
  wire popcount35_19t3_core_095;
  wire popcount35_19t3_core_096;
  wire popcount35_19t3_core_097;
  wire popcount35_19t3_core_103;
  wire popcount35_19t3_core_104;
  wire popcount35_19t3_core_105;
  wire popcount35_19t3_core_106;
  wire popcount35_19t3_core_107;
  wire popcount35_19t3_core_108;
  wire popcount35_19t3_core_109_not;
  wire popcount35_19t3_core_110;
  wire popcount35_19t3_core_111;
  wire popcount35_19t3_core_112;
  wire popcount35_19t3_core_113;
  wire popcount35_19t3_core_114;
  wire popcount35_19t3_core_117;
  wire popcount35_19t3_core_118;
  wire popcount35_19t3_core_119;
  wire popcount35_19t3_core_120;
  wire popcount35_19t3_core_121;
  wire popcount35_19t3_core_122;
  wire popcount35_19t3_core_123;
  wire popcount35_19t3_core_124;
  wire popcount35_19t3_core_125;
  wire popcount35_19t3_core_126;
  wire popcount35_19t3_core_127;
  wire popcount35_19t3_core_129;
  wire popcount35_19t3_core_130;
  wire popcount35_19t3_core_131;
  wire popcount35_19t3_core_132;
  wire popcount35_19t3_core_133;
  wire popcount35_19t3_core_134;
  wire popcount35_19t3_core_135;
  wire popcount35_19t3_core_136;
  wire popcount35_19t3_core_137;
  wire popcount35_19t3_core_139;
  wire popcount35_19t3_core_140;
  wire popcount35_19t3_core_141;
  wire popcount35_19t3_core_143;
  wire popcount35_19t3_core_145;
  wire popcount35_19t3_core_148;
  wire popcount35_19t3_core_152;
  wire popcount35_19t3_core_153;
  wire popcount35_19t3_core_156;
  wire popcount35_19t3_core_157;
  wire popcount35_19t3_core_158;
  wire popcount35_19t3_core_161;
  wire popcount35_19t3_core_162;
  wire popcount35_19t3_core_163;
  wire popcount35_19t3_core_165;
  wire popcount35_19t3_core_167;
  wire popcount35_19t3_core_168;
  wire popcount35_19t3_core_171;
  wire popcount35_19t3_core_174;
  wire popcount35_19t3_core_175;
  wire popcount35_19t3_core_177;
  wire popcount35_19t3_core_178;
  wire popcount35_19t3_core_179;
  wire popcount35_19t3_core_180;
  wire popcount35_19t3_core_181;
  wire popcount35_19t3_core_182;
  wire popcount35_19t3_core_183;
  wire popcount35_19t3_core_184;
  wire popcount35_19t3_core_185;
  wire popcount35_19t3_core_187;
  wire popcount35_19t3_core_191;
  wire popcount35_19t3_core_192;
  wire popcount35_19t3_core_193;
  wire popcount35_19t3_core_195;
  wire popcount35_19t3_core_196;
  wire popcount35_19t3_core_197;
  wire popcount35_19t3_core_199;
  wire popcount35_19t3_core_200;
  wire popcount35_19t3_core_201;
  wire popcount35_19t3_core_203;
  wire popcount35_19t3_core_204;
  wire popcount35_19t3_core_205;
  wire popcount35_19t3_core_208;
  wire popcount35_19t3_core_209_not;
  wire popcount35_19t3_core_210;
  wire popcount35_19t3_core_211;
  wire popcount35_19t3_core_213;
  wire popcount35_19t3_core_214;
  wire popcount35_19t3_core_215;
  wire popcount35_19t3_core_216;
  wire popcount35_19t3_core_218;
  wire popcount35_19t3_core_223;
  wire popcount35_19t3_core_224;
  wire popcount35_19t3_core_225;
  wire popcount35_19t3_core_226;
  wire popcount35_19t3_core_227;
  wire popcount35_19t3_core_228;
  wire popcount35_19t3_core_233;
  wire popcount35_19t3_core_236;
  wire popcount35_19t3_core_237;
  wire popcount35_19t3_core_239;
  wire popcount35_19t3_core_240;
  wire popcount35_19t3_core_243;
  wire popcount35_19t3_core_244;
  wire popcount35_19t3_core_245;
  wire popcount35_19t3_core_249;
  wire popcount35_19t3_core_250;
  wire popcount35_19t3_core_252;
  wire popcount35_19t3_core_253;
  wire popcount35_19t3_core_254;
  wire popcount35_19t3_core_256;
  wire popcount35_19t3_core_257;
  wire popcount35_19t3_core_258;
  wire popcount35_19t3_core_262;
  wire popcount35_19t3_core_263;
  wire popcount35_19t3_core_264;

  assign popcount35_19t3_core_037 = ~(input_a[27] | input_a[2]);
  assign popcount35_19t3_core_038 = input_a[0] | input_a[8];
  assign popcount35_19t3_core_039 = ~(input_a[21] | input_a[3]);
  assign popcount35_19t3_core_040 = input_a[31] & input_a[18];
  assign popcount35_19t3_core_041 = ~(input_a[13] | input_a[18]);
  assign popcount35_19t3_core_042 = input_a[2] | input_a[5];
  assign popcount35_19t3_core_043_not = ~input_a[11];
  assign popcount35_19t3_core_044 = input_a[15] ^ input_a[29];
  assign popcount35_19t3_core_047 = input_a[20] | input_a[8];
  assign popcount35_19t3_core_049 = ~input_a[33];
  assign popcount35_19t3_core_050 = ~input_a[8];
  assign popcount35_19t3_core_051 = ~input_a[7];
  assign popcount35_19t3_core_052 = input_a[27] ^ input_a[23];
  assign popcount35_19t3_core_055 = ~(input_a[6] & input_a[18]);
  assign popcount35_19t3_core_057 = ~(input_a[9] | input_a[24]);
  assign popcount35_19t3_core_060 = ~(input_a[32] ^ input_a[12]);
  assign popcount35_19t3_core_061 = ~input_a[9];
  assign popcount35_19t3_core_065 = ~input_a[6];
  assign popcount35_19t3_core_066 = input_a[5] & input_a[15];
  assign popcount35_19t3_core_067 = ~(input_a[10] | input_a[4]);
  assign popcount35_19t3_core_069 = input_a[9] & input_a[15];
  assign popcount35_19t3_core_070 = ~input_a[16];
  assign popcount35_19t3_core_071 = ~(input_a[23] | input_a[32]);
  assign popcount35_19t3_core_073 = ~input_a[32];
  assign popcount35_19t3_core_074_not = ~input_a[2];
  assign popcount35_19t3_core_075 = ~(input_a[29] ^ input_a[14]);
  assign popcount35_19t3_core_076 = input_a[31] & input_a[11];
  assign popcount35_19t3_core_077 = input_a[10] | input_a[22];
  assign popcount35_19t3_core_079 = ~input_a[19];
  assign popcount35_19t3_core_082 = ~(input_a[1] | input_a[6]);
  assign popcount35_19t3_core_083 = ~(input_a[19] ^ input_a[16]);
  assign popcount35_19t3_core_085 = ~(input_a[3] & input_a[19]);
  assign popcount35_19t3_core_089 = ~(input_a[33] & input_a[8]);
  assign popcount35_19t3_core_090 = ~input_a[32];
  assign popcount35_19t3_core_091 = ~(input_a[30] | input_a[30]);
  assign popcount35_19t3_core_093 = ~(input_a[0] | input_a[24]);
  assign popcount35_19t3_core_094 = input_a[1] & input_a[25];
  assign popcount35_19t3_core_095 = input_a[23] & input_a[17];
  assign popcount35_19t3_core_096 = input_a[28] | input_a[32];
  assign popcount35_19t3_core_097 = input_a[2] ^ input_a[30];
  assign popcount35_19t3_core_103 = ~(input_a[34] | input_a[14]);
  assign popcount35_19t3_core_104 = ~(input_a[9] ^ input_a[28]);
  assign popcount35_19t3_core_105 = ~(input_a[1] | input_a[33]);
  assign popcount35_19t3_core_106 = ~(input_a[31] & input_a[20]);
  assign popcount35_19t3_core_107 = ~(input_a[29] & input_a[18]);
  assign popcount35_19t3_core_108 = input_a[1] ^ input_a[15];
  assign popcount35_19t3_core_109_not = ~input_a[23];
  assign popcount35_19t3_core_110 = ~input_a[23];
  assign popcount35_19t3_core_111 = ~(input_a[27] ^ input_a[21]);
  assign popcount35_19t3_core_112 = ~input_a[21];
  assign popcount35_19t3_core_113 = input_a[27] & input_a[31];
  assign popcount35_19t3_core_114 = input_a[20] | input_a[3];
  assign popcount35_19t3_core_117 = input_a[16] | input_a[20];
  assign popcount35_19t3_core_118 = input_a[31] ^ input_a[25];
  assign popcount35_19t3_core_119 = ~(input_a[34] | input_a[32]);
  assign popcount35_19t3_core_120 = ~(input_a[10] ^ input_a[11]);
  assign popcount35_19t3_core_121 = ~(input_a[10] & input_a[8]);
  assign popcount35_19t3_core_122 = ~input_a[30];
  assign popcount35_19t3_core_123 = input_a[14] | input_a[9];
  assign popcount35_19t3_core_124 = ~input_a[10];
  assign popcount35_19t3_core_125 = input_a[19] | input_a[12];
  assign popcount35_19t3_core_126 = ~(input_a[6] ^ input_a[30]);
  assign popcount35_19t3_core_127 = input_a[30] & input_a[14];
  assign popcount35_19t3_core_129 = ~(input_a[11] | input_a[33]);
  assign popcount35_19t3_core_130 = ~input_a[13];
  assign popcount35_19t3_core_131 = input_a[20] | input_a[21];
  assign popcount35_19t3_core_132 = input_a[4] & input_a[5];
  assign popcount35_19t3_core_133 = input_a[9] ^ input_a[15];
  assign popcount35_19t3_core_134 = ~(input_a[16] & input_a[19]);
  assign popcount35_19t3_core_135 = ~input_a[4];
  assign popcount35_19t3_core_136 = ~(input_a[6] | input_a[17]);
  assign popcount35_19t3_core_137 = ~(input_a[20] & input_a[5]);
  assign popcount35_19t3_core_139 = ~(input_a[23] & input_a[24]);
  assign popcount35_19t3_core_140 = ~(input_a[25] | input_a[2]);
  assign popcount35_19t3_core_141 = input_a[11] & input_a[33];
  assign popcount35_19t3_core_143 = input_a[6] ^ input_a[17];
  assign popcount35_19t3_core_145 = input_a[31] & input_a[22];
  assign popcount35_19t3_core_148 = ~(input_a[25] | input_a[4]);
  assign popcount35_19t3_core_152 = input_a[10] | input_a[31];
  assign popcount35_19t3_core_153 = ~(input_a[4] ^ input_a[17]);
  assign popcount35_19t3_core_156 = ~input_a[7];
  assign popcount35_19t3_core_157 = input_a[25] | input_a[31];
  assign popcount35_19t3_core_158 = ~(input_a[13] ^ input_a[7]);
  assign popcount35_19t3_core_161 = ~(input_a[34] ^ input_a[26]);
  assign popcount35_19t3_core_162 = ~(input_a[18] & input_a[24]);
  assign popcount35_19t3_core_163 = ~(input_a[22] ^ input_a[24]);
  assign popcount35_19t3_core_165 = ~(input_a[7] & input_a[33]);
  assign popcount35_19t3_core_167 = ~(input_a[29] & input_a[3]);
  assign popcount35_19t3_core_168 = ~(input_a[22] ^ input_a[26]);
  assign popcount35_19t3_core_171 = ~(input_a[34] ^ input_a[29]);
  assign popcount35_19t3_core_174 = ~(input_a[6] & input_a[24]);
  assign popcount35_19t3_core_175 = ~(input_a[1] | input_a[21]);
  assign popcount35_19t3_core_177 = input_a[33] & input_a[9];
  assign popcount35_19t3_core_178 = ~input_a[14];
  assign popcount35_19t3_core_179 = input_a[15] ^ input_a[25];
  assign popcount35_19t3_core_180 = ~input_a[7];
  assign popcount35_19t3_core_181 = ~input_a[14];
  assign popcount35_19t3_core_182 = ~(input_a[6] | input_a[11]);
  assign popcount35_19t3_core_183 = ~(input_a[19] & input_a[5]);
  assign popcount35_19t3_core_184 = ~(input_a[14] & input_a[18]);
  assign popcount35_19t3_core_185 = ~(input_a[10] | input_a[21]);
  assign popcount35_19t3_core_187 = input_a[0] & input_a[5];
  assign popcount35_19t3_core_191 = input_a[16] ^ input_a[28];
  assign popcount35_19t3_core_192 = ~(input_a[28] & input_a[8]);
  assign popcount35_19t3_core_193 = ~(input_a[29] & input_a[7]);
  assign popcount35_19t3_core_195 = input_a[27] & input_a[17];
  assign popcount35_19t3_core_196 = input_a[7] | input_a[21];
  assign popcount35_19t3_core_197 = ~(input_a[13] & input_a[24]);
  assign popcount35_19t3_core_199 = input_a[6] & input_a[24];
  assign popcount35_19t3_core_200 = ~(input_a[14] | input_a[0]);
  assign popcount35_19t3_core_201 = input_a[1] | input_a[6];
  assign popcount35_19t3_core_203 = input_a[34] & input_a[20];
  assign popcount35_19t3_core_204 = input_a[27] | input_a[25];
  assign popcount35_19t3_core_205 = ~input_a[34];
  assign popcount35_19t3_core_208 = ~(input_a[6] & input_a[25]);
  assign popcount35_19t3_core_209_not = ~input_a[10];
  assign popcount35_19t3_core_210 = input_a[11] | input_a[28];
  assign popcount35_19t3_core_211 = ~(input_a[4] | input_a[23]);
  assign popcount35_19t3_core_213 = input_a[6] & input_a[13];
  assign popcount35_19t3_core_214 = ~input_a[34];
  assign popcount35_19t3_core_215 = input_a[3] & input_a[9];
  assign popcount35_19t3_core_216 = ~(input_a[4] & input_a[9]);
  assign popcount35_19t3_core_218 = input_a[15] & input_a[20];
  assign popcount35_19t3_core_223 = ~(input_a[1] | input_a[8]);
  assign popcount35_19t3_core_224 = input_a[10] ^ input_a[1];
  assign popcount35_19t3_core_225 = input_a[23] | input_a[27];
  assign popcount35_19t3_core_226 = ~(input_a[13] ^ input_a[28]);
  assign popcount35_19t3_core_227 = ~(input_a[30] ^ input_a[25]);
  assign popcount35_19t3_core_228 = input_a[5] & input_a[15];
  assign popcount35_19t3_core_233 = ~(input_a[10] | input_a[22]);
  assign popcount35_19t3_core_236 = ~(input_a[33] | input_a[28]);
  assign popcount35_19t3_core_237 = ~input_a[8];
  assign popcount35_19t3_core_239 = ~(input_a[7] & input_a[23]);
  assign popcount35_19t3_core_240 = ~(input_a[8] | input_a[34]);
  assign popcount35_19t3_core_243 = ~(input_a[20] | input_a[6]);
  assign popcount35_19t3_core_244 = ~input_a[3];
  assign popcount35_19t3_core_245 = input_a[31] ^ input_a[17];
  assign popcount35_19t3_core_249 = ~(input_a[2] | input_a[15]);
  assign popcount35_19t3_core_250 = input_a[0] ^ input_a[11];
  assign popcount35_19t3_core_252 = input_a[24] | input_a[16];
  assign popcount35_19t3_core_253 = ~(input_a[34] | input_a[31]);
  assign popcount35_19t3_core_254 = input_a[13] | input_a[30];
  assign popcount35_19t3_core_256 = ~input_a[22];
  assign popcount35_19t3_core_257 = ~(input_a[13] | input_a[13]);
  assign popcount35_19t3_core_258 = input_a[1] | input_a[14];
  assign popcount35_19t3_core_262 = ~(input_a[18] | input_a[21]);
  assign popcount35_19t3_core_263 = ~input_a[25];
  assign popcount35_19t3_core_264 = input_a[3] & input_a[17];

  assign popcount35_19t3_out[0] = input_a[19];
  assign popcount35_19t3_out[1] = input_a[3];
  assign popcount35_19t3_out[2] = input_a[5];
  assign popcount35_19t3_out[3] = 1'b0;
  assign popcount35_19t3_out[4] = 1'b1;
  assign popcount35_19t3_out[5] = 1'b0;
endmodule