// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.30917
// WCE=17.0
// EP=0.864166%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_vhmp(input [33:0] input_a, output [5:0] popcount34_vhmp_out);
  wire popcount34_vhmp_core_037;
  wire popcount34_vhmp_core_041;
  wire popcount34_vhmp_core_043;
  wire popcount34_vhmp_core_047;
  wire popcount34_vhmp_core_049;
  wire popcount34_vhmp_core_051;
  wire popcount34_vhmp_core_052;
  wire popcount34_vhmp_core_053;
  wire popcount34_vhmp_core_054;
  wire popcount34_vhmp_core_055_not;
  wire popcount34_vhmp_core_056;
  wire popcount34_vhmp_core_057;
  wire popcount34_vhmp_core_058;
  wire popcount34_vhmp_core_063;
  wire popcount34_vhmp_core_065;
  wire popcount34_vhmp_core_070;
  wire popcount34_vhmp_core_071;
  wire popcount34_vhmp_core_072;
  wire popcount34_vhmp_core_073;
  wire popcount34_vhmp_core_074;
  wire popcount34_vhmp_core_075;
  wire popcount34_vhmp_core_077_not;
  wire popcount34_vhmp_core_079;
  wire popcount34_vhmp_core_081;
  wire popcount34_vhmp_core_084;
  wire popcount34_vhmp_core_085;
  wire popcount34_vhmp_core_086;
  wire popcount34_vhmp_core_087;
  wire popcount34_vhmp_core_089;
  wire popcount34_vhmp_core_090;
  wire popcount34_vhmp_core_092;
  wire popcount34_vhmp_core_093;
  wire popcount34_vhmp_core_094;
  wire popcount34_vhmp_core_095;
  wire popcount34_vhmp_core_096;
  wire popcount34_vhmp_core_098;
  wire popcount34_vhmp_core_099;
  wire popcount34_vhmp_core_100;
  wire popcount34_vhmp_core_101;
  wire popcount34_vhmp_core_102;
  wire popcount34_vhmp_core_103;
  wire popcount34_vhmp_core_104;
  wire popcount34_vhmp_core_105;
  wire popcount34_vhmp_core_106;
  wire popcount34_vhmp_core_110;
  wire popcount34_vhmp_core_111;
  wire popcount34_vhmp_core_112;
  wire popcount34_vhmp_core_113;
  wire popcount34_vhmp_core_115;
  wire popcount34_vhmp_core_117;
  wire popcount34_vhmp_core_118;
  wire popcount34_vhmp_core_119;
  wire popcount34_vhmp_core_120;
  wire popcount34_vhmp_core_124;
  wire popcount34_vhmp_core_125;
  wire popcount34_vhmp_core_126;
  wire popcount34_vhmp_core_127;
  wire popcount34_vhmp_core_128;
  wire popcount34_vhmp_core_129;
  wire popcount34_vhmp_core_130;
  wire popcount34_vhmp_core_131;
  wire popcount34_vhmp_core_133;
  wire popcount34_vhmp_core_134_not;
  wire popcount34_vhmp_core_135;
  wire popcount34_vhmp_core_140;
  wire popcount34_vhmp_core_141;
  wire popcount34_vhmp_core_144;
  wire popcount34_vhmp_core_145_not;
  wire popcount34_vhmp_core_150;
  wire popcount34_vhmp_core_151;
  wire popcount34_vhmp_core_152;
  wire popcount34_vhmp_core_153;
  wire popcount34_vhmp_core_154;
  wire popcount34_vhmp_core_155;
  wire popcount34_vhmp_core_160;
  wire popcount34_vhmp_core_161;
  wire popcount34_vhmp_core_162_not;
  wire popcount34_vhmp_core_163;
  wire popcount34_vhmp_core_164;
  wire popcount34_vhmp_core_165;
  wire popcount34_vhmp_core_166;
  wire popcount34_vhmp_core_168;
  wire popcount34_vhmp_core_169;
  wire popcount34_vhmp_core_170;
  wire popcount34_vhmp_core_172;
  wire popcount34_vhmp_core_173;
  wire popcount34_vhmp_core_174;
  wire popcount34_vhmp_core_175;
  wire popcount34_vhmp_core_178;
  wire popcount34_vhmp_core_179;
  wire popcount34_vhmp_core_180;
  wire popcount34_vhmp_core_181;
  wire popcount34_vhmp_core_182;
  wire popcount34_vhmp_core_184;
  wire popcount34_vhmp_core_186;
  wire popcount34_vhmp_core_187_not;
  wire popcount34_vhmp_core_188;
  wire popcount34_vhmp_core_189;
  wire popcount34_vhmp_core_191;
  wire popcount34_vhmp_core_192;
  wire popcount34_vhmp_core_193;
  wire popcount34_vhmp_core_194;
  wire popcount34_vhmp_core_196;
  wire popcount34_vhmp_core_197;
  wire popcount34_vhmp_core_198;
  wire popcount34_vhmp_core_199;
  wire popcount34_vhmp_core_201;
  wire popcount34_vhmp_core_202;
  wire popcount34_vhmp_core_203_not;
  wire popcount34_vhmp_core_205;
  wire popcount34_vhmp_core_207;
  wire popcount34_vhmp_core_210;
  wire popcount34_vhmp_core_213;
  wire popcount34_vhmp_core_214;
  wire popcount34_vhmp_core_215_not;
  wire popcount34_vhmp_core_216;
  wire popcount34_vhmp_core_217;
  wire popcount34_vhmp_core_220;
  wire popcount34_vhmp_core_221;
  wire popcount34_vhmp_core_223;
  wire popcount34_vhmp_core_224;
  wire popcount34_vhmp_core_225;
  wire popcount34_vhmp_core_226;
  wire popcount34_vhmp_core_228;
  wire popcount34_vhmp_core_230;
  wire popcount34_vhmp_core_232;
  wire popcount34_vhmp_core_234;
  wire popcount34_vhmp_core_235;
  wire popcount34_vhmp_core_236_not;
  wire popcount34_vhmp_core_237;
  wire popcount34_vhmp_core_238;
  wire popcount34_vhmp_core_239;
  wire popcount34_vhmp_core_240;
  wire popcount34_vhmp_core_243;
  wire popcount34_vhmp_core_244;
  wire popcount34_vhmp_core_246;
  wire popcount34_vhmp_core_247;
  wire popcount34_vhmp_core_251;

  assign popcount34_vhmp_core_037 = ~(input_a[29] & input_a[18]);
  assign popcount34_vhmp_core_041 = input_a[3] & input_a[9];
  assign popcount34_vhmp_core_043 = input_a[22] & input_a[13];
  assign popcount34_vhmp_core_047 = input_a[27] ^ input_a[24];
  assign popcount34_vhmp_core_049 = input_a[6] | input_a[22];
  assign popcount34_vhmp_core_051 = input_a[2] ^ input_a[33];
  assign popcount34_vhmp_core_052 = ~(input_a[3] ^ input_a[14]);
  assign popcount34_vhmp_core_053 = input_a[20] | input_a[32];
  assign popcount34_vhmp_core_054 = ~(input_a[25] ^ input_a[28]);
  assign popcount34_vhmp_core_055_not = ~input_a[3];
  assign popcount34_vhmp_core_056 = input_a[26] & input_a[7];
  assign popcount34_vhmp_core_057 = input_a[12] ^ input_a[25];
  assign popcount34_vhmp_core_058 = input_a[7] | input_a[18];
  assign popcount34_vhmp_core_063 = ~(input_a[13] & input_a[12]);
  assign popcount34_vhmp_core_065 = ~(input_a[9] ^ input_a[30]);
  assign popcount34_vhmp_core_070 = ~input_a[29];
  assign popcount34_vhmp_core_071 = ~input_a[16];
  assign popcount34_vhmp_core_072 = ~(input_a[20] | input_a[19]);
  assign popcount34_vhmp_core_073 = ~(input_a[21] & input_a[4]);
  assign popcount34_vhmp_core_074 = ~(input_a[22] & input_a[11]);
  assign popcount34_vhmp_core_075 = input_a[6] ^ input_a[8];
  assign popcount34_vhmp_core_077_not = ~input_a[31];
  assign popcount34_vhmp_core_079 = input_a[13] & input_a[17];
  assign popcount34_vhmp_core_081 = ~(input_a[11] | input_a[32]);
  assign popcount34_vhmp_core_084 = ~(input_a[26] ^ input_a[5]);
  assign popcount34_vhmp_core_085 = ~(input_a[22] & input_a[23]);
  assign popcount34_vhmp_core_086 = ~(input_a[16] & input_a[23]);
  assign popcount34_vhmp_core_087 = ~(input_a[8] | input_a[13]);
  assign popcount34_vhmp_core_089 = ~(input_a[12] | input_a[22]);
  assign popcount34_vhmp_core_090 = ~(input_a[7] | input_a[32]);
  assign popcount34_vhmp_core_092 = ~(input_a[25] ^ input_a[24]);
  assign popcount34_vhmp_core_093 = input_a[31] | input_a[9];
  assign popcount34_vhmp_core_094 = ~(input_a[9] ^ input_a[19]);
  assign popcount34_vhmp_core_095 = ~(input_a[4] ^ input_a[9]);
  assign popcount34_vhmp_core_096 = input_a[9] | input_a[2];
  assign popcount34_vhmp_core_098 = ~input_a[4];
  assign popcount34_vhmp_core_099 = ~(input_a[30] & input_a[7]);
  assign popcount34_vhmp_core_100 = ~(input_a[32] & input_a[5]);
  assign popcount34_vhmp_core_101 = input_a[26] & input_a[9];
  assign popcount34_vhmp_core_102 = ~(input_a[32] ^ input_a[32]);
  assign popcount34_vhmp_core_103 = ~input_a[24];
  assign popcount34_vhmp_core_104 = input_a[6] ^ input_a[18];
  assign popcount34_vhmp_core_105 = input_a[13] ^ input_a[15];
  assign popcount34_vhmp_core_106 = input_a[21] & input_a[21];
  assign popcount34_vhmp_core_110 = ~input_a[3];
  assign popcount34_vhmp_core_111 = ~(input_a[13] ^ input_a[13]);
  assign popcount34_vhmp_core_112 = ~(input_a[11] & input_a[14]);
  assign popcount34_vhmp_core_113 = input_a[19] ^ input_a[19];
  assign popcount34_vhmp_core_115 = ~(input_a[11] | input_a[31]);
  assign popcount34_vhmp_core_117 = ~(input_a[0] ^ input_a[9]);
  assign popcount34_vhmp_core_118 = input_a[18] | input_a[14];
  assign popcount34_vhmp_core_119 = ~(input_a[30] & input_a[29]);
  assign popcount34_vhmp_core_120 = ~input_a[31];
  assign popcount34_vhmp_core_124 = input_a[33] & input_a[1];
  assign popcount34_vhmp_core_125 = ~(input_a[21] | input_a[20]);
  assign popcount34_vhmp_core_126 = ~(input_a[29] & input_a[3]);
  assign popcount34_vhmp_core_127 = ~(input_a[12] | input_a[21]);
  assign popcount34_vhmp_core_128 = ~(input_a[21] & input_a[16]);
  assign popcount34_vhmp_core_129 = input_a[9] | input_a[19];
  assign popcount34_vhmp_core_130 = input_a[24] ^ input_a[23];
  assign popcount34_vhmp_core_131 = ~(input_a[1] ^ input_a[29]);
  assign popcount34_vhmp_core_133 = ~input_a[22];
  assign popcount34_vhmp_core_134_not = ~input_a[31];
  assign popcount34_vhmp_core_135 = ~(input_a[30] ^ input_a[8]);
  assign popcount34_vhmp_core_140 = input_a[0] | input_a[15];
  assign popcount34_vhmp_core_141 = ~input_a[33];
  assign popcount34_vhmp_core_144 = ~(input_a[15] & input_a[30]);
  assign popcount34_vhmp_core_145_not = ~input_a[2];
  assign popcount34_vhmp_core_150 = ~(input_a[23] & input_a[3]);
  assign popcount34_vhmp_core_151 = input_a[9] & input_a[12];
  assign popcount34_vhmp_core_152 = ~(input_a[30] ^ input_a[21]);
  assign popcount34_vhmp_core_153 = input_a[2] & input_a[22];
  assign popcount34_vhmp_core_154 = ~(input_a[5] & input_a[30]);
  assign popcount34_vhmp_core_155 = ~(input_a[10] | input_a[21]);
  assign popcount34_vhmp_core_160 = ~(input_a[4] & input_a[32]);
  assign popcount34_vhmp_core_161 = input_a[33] | input_a[29];
  assign popcount34_vhmp_core_162_not = ~input_a[11];
  assign popcount34_vhmp_core_163 = ~input_a[22];
  assign popcount34_vhmp_core_164 = input_a[16] & input_a[13];
  assign popcount34_vhmp_core_165 = ~(input_a[20] | input_a[26]);
  assign popcount34_vhmp_core_166 = input_a[25] & input_a[13];
  assign popcount34_vhmp_core_168 = ~input_a[17];
  assign popcount34_vhmp_core_169 = ~(input_a[5] ^ input_a[29]);
  assign popcount34_vhmp_core_170 = ~(input_a[23] | input_a[19]);
  assign popcount34_vhmp_core_172 = input_a[24] ^ input_a[13];
  assign popcount34_vhmp_core_173 = input_a[27] | input_a[3];
  assign popcount34_vhmp_core_174 = ~(input_a[29] ^ input_a[24]);
  assign popcount34_vhmp_core_175 = ~(input_a[20] ^ input_a[9]);
  assign popcount34_vhmp_core_178 = ~input_a[16];
  assign popcount34_vhmp_core_179 = input_a[27] & input_a[4];
  assign popcount34_vhmp_core_180 = input_a[8] & input_a[11];
  assign popcount34_vhmp_core_181 = input_a[22] & input_a[26];
  assign popcount34_vhmp_core_182 = ~(input_a[30] | input_a[5]);
  assign popcount34_vhmp_core_184 = input_a[19] ^ input_a[8];
  assign popcount34_vhmp_core_186 = input_a[3] & input_a[2];
  assign popcount34_vhmp_core_187_not = ~input_a[0];
  assign popcount34_vhmp_core_188 = ~input_a[27];
  assign popcount34_vhmp_core_189 = input_a[1] & input_a[13];
  assign popcount34_vhmp_core_191 = ~(input_a[23] & input_a[26]);
  assign popcount34_vhmp_core_192 = input_a[11] ^ input_a[6];
  assign popcount34_vhmp_core_193 = ~input_a[16];
  assign popcount34_vhmp_core_194 = input_a[15] & input_a[12];
  assign popcount34_vhmp_core_196 = ~(input_a[12] | input_a[15]);
  assign popcount34_vhmp_core_197 = ~input_a[20];
  assign popcount34_vhmp_core_198 = input_a[4] & input_a[22];
  assign popcount34_vhmp_core_199 = input_a[14] | input_a[4];
  assign popcount34_vhmp_core_201 = input_a[19] & input_a[7];
  assign popcount34_vhmp_core_202 = input_a[3] | input_a[23];
  assign popcount34_vhmp_core_203_not = ~input_a[11];
  assign popcount34_vhmp_core_205 = ~(input_a[6] & input_a[10]);
  assign popcount34_vhmp_core_207 = ~(input_a[24] & input_a[31]);
  assign popcount34_vhmp_core_210 = ~(input_a[2] | input_a[6]);
  assign popcount34_vhmp_core_213 = ~(input_a[26] & input_a[12]);
  assign popcount34_vhmp_core_214 = input_a[24] ^ input_a[19];
  assign popcount34_vhmp_core_215_not = ~input_a[20];
  assign popcount34_vhmp_core_216 = ~(input_a[24] & input_a[30]);
  assign popcount34_vhmp_core_217 = input_a[19] | input_a[15];
  assign popcount34_vhmp_core_220 = ~(input_a[19] | input_a[24]);
  assign popcount34_vhmp_core_221 = input_a[13] ^ input_a[8];
  assign popcount34_vhmp_core_223 = ~input_a[26];
  assign popcount34_vhmp_core_224 = input_a[19] ^ input_a[8];
  assign popcount34_vhmp_core_225 = ~(input_a[15] ^ input_a[31]);
  assign popcount34_vhmp_core_226 = input_a[26] ^ input_a[31];
  assign popcount34_vhmp_core_228 = input_a[31] ^ input_a[16];
  assign popcount34_vhmp_core_230 = input_a[15] | input_a[24];
  assign popcount34_vhmp_core_232 = input_a[13] & input_a[17];
  assign popcount34_vhmp_core_234 = ~input_a[14];
  assign popcount34_vhmp_core_235 = ~(input_a[14] & input_a[5]);
  assign popcount34_vhmp_core_236_not = ~input_a[18];
  assign popcount34_vhmp_core_237 = ~(input_a[24] ^ input_a[21]);
  assign popcount34_vhmp_core_238 = ~(input_a[4] | input_a[23]);
  assign popcount34_vhmp_core_239 = ~(input_a[15] & input_a[11]);
  assign popcount34_vhmp_core_240 = input_a[17] & input_a[17];
  assign popcount34_vhmp_core_243 = ~(input_a[6] ^ input_a[14]);
  assign popcount34_vhmp_core_244 = input_a[24] | input_a[6];
  assign popcount34_vhmp_core_246 = ~input_a[12];
  assign popcount34_vhmp_core_247 = ~(input_a[14] | input_a[11]);
  assign popcount34_vhmp_core_251 = ~(input_a[22] & input_a[2]);

  assign popcount34_vhmp_out[0] = 1'b0;
  assign popcount34_vhmp_out[1] = input_a[24];
  assign popcount34_vhmp_out[2] = 1'b0;
  assign popcount34_vhmp_out[3] = 1'b0;
  assign popcount34_vhmp_out[4] = 1'b1;
  assign popcount34_vhmp_out[5] = 1'b0;
endmodule