// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.75851
// WCE=16.0
// EP=0.931808%
// Printed PDK parameters:
//  Area=228420.0
//  Delay=565706.94
//  Power=878.4483

module popcount24_dyrt(input [23:0] input_a, output [4:0] popcount24_dyrt_out);
  wire popcount24_dyrt_core_026;
  wire popcount24_dyrt_core_030;
  wire popcount24_dyrt_core_031;
  wire popcount24_dyrt_core_032;
  wire popcount24_dyrt_core_034;
  wire popcount24_dyrt_core_035;
  wire popcount24_dyrt_core_037;
  wire popcount24_dyrt_core_038;
  wire popcount24_dyrt_core_039;
  wire popcount24_dyrt_core_042;
  wire popcount24_dyrt_core_044;
  wire popcount24_dyrt_core_045;
  wire popcount24_dyrt_core_046;
  wire popcount24_dyrt_core_047;
  wire popcount24_dyrt_core_049;
  wire popcount24_dyrt_core_052;
  wire popcount24_dyrt_core_053;
  wire popcount24_dyrt_core_054;
  wire popcount24_dyrt_core_055;
  wire popcount24_dyrt_core_056;
  wire popcount24_dyrt_core_057;
  wire popcount24_dyrt_core_058;
  wire popcount24_dyrt_core_060;
  wire popcount24_dyrt_core_063;
  wire popcount24_dyrt_core_064;
  wire popcount24_dyrt_core_065;
  wire popcount24_dyrt_core_066;
  wire popcount24_dyrt_core_068;
  wire popcount24_dyrt_core_069;
  wire popcount24_dyrt_core_070;
  wire popcount24_dyrt_core_071;
  wire popcount24_dyrt_core_074;
  wire popcount24_dyrt_core_075;
  wire popcount24_dyrt_core_076_not;
  wire popcount24_dyrt_core_078;
  wire popcount24_dyrt_core_079;
  wire popcount24_dyrt_core_080;
  wire popcount24_dyrt_core_081;
  wire popcount24_dyrt_core_082;
  wire popcount24_dyrt_core_083;
  wire popcount24_dyrt_core_088;
  wire popcount24_dyrt_core_089;
  wire popcount24_dyrt_core_090;
  wire popcount24_dyrt_core_092;
  wire popcount24_dyrt_core_093;
  wire popcount24_dyrt_core_094;
  wire popcount24_dyrt_core_095;
  wire popcount24_dyrt_core_096;
  wire popcount24_dyrt_core_097;
  wire popcount24_dyrt_core_099;
  wire popcount24_dyrt_core_100;
  wire popcount24_dyrt_core_102;
  wire popcount24_dyrt_core_105_not;
  wire popcount24_dyrt_core_110;
  wire popcount24_dyrt_core_111;
  wire popcount24_dyrt_core_113;
  wire popcount24_dyrt_core_115;
  wire popcount24_dyrt_core_118;
  wire popcount24_dyrt_core_120;
  wire popcount24_dyrt_core_121;
  wire popcount24_dyrt_core_122;
  wire popcount24_dyrt_core_123;
  wire popcount24_dyrt_core_124;
  wire popcount24_dyrt_core_125;
  wire popcount24_dyrt_core_126;
  wire popcount24_dyrt_core_127;
  wire popcount24_dyrt_core_128;
  wire popcount24_dyrt_core_130;
  wire popcount24_dyrt_core_131;
  wire popcount24_dyrt_core_132;
  wire popcount24_dyrt_core_134;
  wire popcount24_dyrt_core_135;
  wire popcount24_dyrt_core_137;
  wire popcount24_dyrt_core_139_not;
  wire popcount24_dyrt_core_140;
  wire popcount24_dyrt_core_141;
  wire popcount24_dyrt_core_142;
  wire popcount24_dyrt_core_143;
  wire popcount24_dyrt_core_144;
  wire popcount24_dyrt_core_145_not;
  wire popcount24_dyrt_core_146_not;
  wire popcount24_dyrt_core_148;
  wire popcount24_dyrt_core_149_not;
  wire popcount24_dyrt_core_150;
  wire popcount24_dyrt_core_151;
  wire popcount24_dyrt_core_153;
  wire popcount24_dyrt_core_154;
  wire popcount24_dyrt_core_155;
  wire popcount24_dyrt_core_156;
  wire popcount24_dyrt_core_157;
  wire popcount24_dyrt_core_160;
  wire popcount24_dyrt_core_163;
  wire popcount24_dyrt_core_166;
  wire popcount24_dyrt_core_168;
  wire popcount24_dyrt_core_169;
  wire popcount24_dyrt_core_170;
  wire popcount24_dyrt_core_172;
  wire popcount24_dyrt_core_173;
  wire popcount24_dyrt_core_174;
  wire popcount24_dyrt_core_175;

  assign popcount24_dyrt_core_026 = ~(input_a[9] | input_a[15]);
  assign popcount24_dyrt_core_030 = ~(input_a[0] | input_a[22]);
  assign popcount24_dyrt_core_031 = ~(input_a[5] ^ input_a[8]);
  assign popcount24_dyrt_core_032 = input_a[9] | input_a[12];
  assign popcount24_dyrt_core_034 = ~(input_a[5] & input_a[4]);
  assign popcount24_dyrt_core_035 = ~(input_a[20] | input_a[9]);
  assign popcount24_dyrt_core_037 = ~input_a[1];
  assign popcount24_dyrt_core_038 = ~(input_a[5] & input_a[22]);
  assign popcount24_dyrt_core_039 = input_a[12] ^ input_a[11];
  assign popcount24_dyrt_core_042 = ~(input_a[11] ^ input_a[22]);
  assign popcount24_dyrt_core_044 = input_a[5] & input_a[9];
  assign popcount24_dyrt_core_045 = ~input_a[23];
  assign popcount24_dyrt_core_046 = ~(input_a[8] ^ input_a[18]);
  assign popcount24_dyrt_core_047 = ~(input_a[3] | input_a[1]);
  assign popcount24_dyrt_core_049 = ~(input_a[22] ^ input_a[7]);
  assign popcount24_dyrt_core_052 = ~(input_a[13] | input_a[7]);
  assign popcount24_dyrt_core_053 = input_a[19] | input_a[12];
  assign popcount24_dyrt_core_054 = ~(input_a[14] | input_a[13]);
  assign popcount24_dyrt_core_055 = ~(input_a[2] & input_a[19]);
  assign popcount24_dyrt_core_056 = input_a[3] ^ input_a[4];
  assign popcount24_dyrt_core_057 = ~(input_a[18] | input_a[13]);
  assign popcount24_dyrt_core_058 = ~(input_a[14] & input_a[3]);
  assign popcount24_dyrt_core_060 = input_a[2] & input_a[6];
  assign popcount24_dyrt_core_063 = ~(input_a[12] & input_a[19]);
  assign popcount24_dyrt_core_064 = ~(input_a[9] & input_a[13]);
  assign popcount24_dyrt_core_065 = ~(input_a[18] ^ input_a[10]);
  assign popcount24_dyrt_core_066 = ~(input_a[16] ^ input_a[2]);
  assign popcount24_dyrt_core_068 = ~(input_a[0] | input_a[21]);
  assign popcount24_dyrt_core_069 = ~input_a[23];
  assign popcount24_dyrt_core_070 = input_a[13] ^ input_a[15];
  assign popcount24_dyrt_core_071 = ~(input_a[9] | input_a[19]);
  assign popcount24_dyrt_core_074 = ~(input_a[18] ^ input_a[15]);
  assign popcount24_dyrt_core_075 = input_a[20] & input_a[10];
  assign popcount24_dyrt_core_076_not = ~input_a[17];
  assign popcount24_dyrt_core_078 = ~(input_a[3] | input_a[22]);
  assign popcount24_dyrt_core_079 = input_a[21] | input_a[20];
  assign popcount24_dyrt_core_080 = ~input_a[23];
  assign popcount24_dyrt_core_081 = input_a[22] ^ input_a[22];
  assign popcount24_dyrt_core_082 = input_a[19] & input_a[21];
  assign popcount24_dyrt_core_083 = input_a[17] ^ input_a[23];
  assign popcount24_dyrt_core_088 = input_a[17] & input_a[16];
  assign popcount24_dyrt_core_089 = input_a[13] & input_a[9];
  assign popcount24_dyrt_core_090 = ~input_a[14];
  assign popcount24_dyrt_core_092 = input_a[9] ^ input_a[15];
  assign popcount24_dyrt_core_093 = ~(input_a[16] & input_a[7]);
  assign popcount24_dyrt_core_094 = ~input_a[23];
  assign popcount24_dyrt_core_095 = input_a[12] & input_a[20];
  assign popcount24_dyrt_core_096 = input_a[16] ^ input_a[22];
  assign popcount24_dyrt_core_097 = input_a[14] ^ input_a[7];
  assign popcount24_dyrt_core_099 = ~(input_a[21] ^ input_a[22]);
  assign popcount24_dyrt_core_100 = ~(input_a[14] ^ input_a[10]);
  assign popcount24_dyrt_core_102 = input_a[4] ^ input_a[16];
  assign popcount24_dyrt_core_105_not = ~input_a[5];
  assign popcount24_dyrt_core_110 = input_a[1] ^ input_a[13];
  assign popcount24_dyrt_core_111 = ~(input_a[18] & input_a[13]);
  assign popcount24_dyrt_core_113 = ~(input_a[21] | input_a[19]);
  assign popcount24_dyrt_core_115 = ~(input_a[15] ^ input_a[9]);
  assign popcount24_dyrt_core_118 = input_a[7] | input_a[16];
  assign popcount24_dyrt_core_120 = ~(input_a[19] & input_a[2]);
  assign popcount24_dyrt_core_121 = input_a[20] ^ input_a[19];
  assign popcount24_dyrt_core_122 = ~(input_a[5] | input_a[4]);
  assign popcount24_dyrt_core_123 = input_a[1] | input_a[15];
  assign popcount24_dyrt_core_124 = input_a[0] & input_a[8];
  assign popcount24_dyrt_core_125 = ~input_a[4];
  assign popcount24_dyrt_core_126 = ~input_a[12];
  assign popcount24_dyrt_core_127 = input_a[11] | input_a[11];
  assign popcount24_dyrt_core_128 = ~input_a[12];
  assign popcount24_dyrt_core_130 = input_a[20] & input_a[12];
  assign popcount24_dyrt_core_131 = input_a[9] & input_a[7];
  assign popcount24_dyrt_core_132 = ~input_a[17];
  assign popcount24_dyrt_core_134 = input_a[22] | input_a[23];
  assign popcount24_dyrt_core_135 = ~input_a[18];
  assign popcount24_dyrt_core_137 = input_a[15] | input_a[18];
  assign popcount24_dyrt_core_139_not = ~input_a[23];
  assign popcount24_dyrt_core_140 = ~(input_a[19] & input_a[20]);
  assign popcount24_dyrt_core_141 = ~(input_a[0] ^ input_a[19]);
  assign popcount24_dyrt_core_142 = ~(input_a[17] & input_a[16]);
  assign popcount24_dyrt_core_143 = ~(input_a[8] | input_a[2]);
  assign popcount24_dyrt_core_144 = input_a[4] | input_a[9];
  assign popcount24_dyrt_core_145_not = ~input_a[22];
  assign popcount24_dyrt_core_146_not = ~input_a[4];
  assign popcount24_dyrt_core_148 = input_a[16] | input_a[3];
  assign popcount24_dyrt_core_149_not = ~input_a[18];
  assign popcount24_dyrt_core_150 = input_a[5] | input_a[5];
  assign popcount24_dyrt_core_151 = ~input_a[14];
  assign popcount24_dyrt_core_153 = ~(input_a[19] ^ input_a[23]);
  assign popcount24_dyrt_core_154 = ~(input_a[22] & input_a[4]);
  assign popcount24_dyrt_core_155 = ~input_a[5];
  assign popcount24_dyrt_core_156 = ~input_a[12];
  assign popcount24_dyrt_core_157 = input_a[19] | input_a[20];
  assign popcount24_dyrt_core_160 = input_a[9] ^ input_a[4];
  assign popcount24_dyrt_core_163 = ~(input_a[21] | input_a[0]);
  assign popcount24_dyrt_core_166 = input_a[3] | input_a[21];
  assign popcount24_dyrt_core_168 = input_a[8] ^ input_a[2];
  assign popcount24_dyrt_core_169 = ~(input_a[8] ^ input_a[20]);
  assign popcount24_dyrt_core_170 = input_a[12] ^ input_a[11];
  assign popcount24_dyrt_core_172 = input_a[10] | input_a[15];
  assign popcount24_dyrt_core_173 = ~(input_a[5] | input_a[22]);
  assign popcount24_dyrt_core_174 = ~input_a[12];
  assign popcount24_dyrt_core_175 = input_a[13] & input_a[4];

  assign popcount24_dyrt_out[0] = input_a[11];
  assign popcount24_dyrt_out[1] = input_a[18];
  assign popcount24_dyrt_out[2] = 1'b0;
  assign popcount24_dyrt_out[3] = popcount24_dyrt_core_094;
  assign popcount24_dyrt_out[4] = input_a[23];
endmodule