// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=3.28464
// WCE=20.0
// EP=0.907855%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_fozj(input [32:0] input_a, output [5:0] popcount33_fozj_out);
  wire popcount33_fozj_core_035;
  wire popcount33_fozj_core_036;
  wire popcount33_fozj_core_037;
  wire popcount33_fozj_core_038;
  wire popcount33_fozj_core_040;
  wire popcount33_fozj_core_041;
  wire popcount33_fozj_core_044;
  wire popcount33_fozj_core_045;
  wire popcount33_fozj_core_048;
  wire popcount33_fozj_core_049_not;
  wire popcount33_fozj_core_050;
  wire popcount33_fozj_core_051;
  wire popcount33_fozj_core_053;
  wire popcount33_fozj_core_054;
  wire popcount33_fozj_core_055;
  wire popcount33_fozj_core_056;
  wire popcount33_fozj_core_059;
  wire popcount33_fozj_core_060;
  wire popcount33_fozj_core_062;
  wire popcount33_fozj_core_063;
  wire popcount33_fozj_core_064;
  wire popcount33_fozj_core_065_not;
  wire popcount33_fozj_core_066;
  wire popcount33_fozj_core_067;
  wire popcount33_fozj_core_068;
  wire popcount33_fozj_core_074;
  wire popcount33_fozj_core_075;
  wire popcount33_fozj_core_079;
  wire popcount33_fozj_core_080;
  wire popcount33_fozj_core_081;
  wire popcount33_fozj_core_082;
  wire popcount33_fozj_core_083;
  wire popcount33_fozj_core_084;
  wire popcount33_fozj_core_085_not;
  wire popcount33_fozj_core_087;
  wire popcount33_fozj_core_090;
  wire popcount33_fozj_core_091;
  wire popcount33_fozj_core_092;
  wire popcount33_fozj_core_093;
  wire popcount33_fozj_core_096;
  wire popcount33_fozj_core_101;
  wire popcount33_fozj_core_102;
  wire popcount33_fozj_core_104_not;
  wire popcount33_fozj_core_105;
  wire popcount33_fozj_core_107;
  wire popcount33_fozj_core_108;
  wire popcount33_fozj_core_110;
  wire popcount33_fozj_core_111;
  wire popcount33_fozj_core_112;
  wire popcount33_fozj_core_113;
  wire popcount33_fozj_core_114;
  wire popcount33_fozj_core_115;
  wire popcount33_fozj_core_116;
  wire popcount33_fozj_core_117;
  wire popcount33_fozj_core_121;
  wire popcount33_fozj_core_122;
  wire popcount33_fozj_core_123;
  wire popcount33_fozj_core_124;
  wire popcount33_fozj_core_125;
  wire popcount33_fozj_core_126;
  wire popcount33_fozj_core_130;
  wire popcount33_fozj_core_133;
  wire popcount33_fozj_core_134;
  wire popcount33_fozj_core_137;
  wire popcount33_fozj_core_139;
  wire popcount33_fozj_core_140;
  wire popcount33_fozj_core_142;
  wire popcount33_fozj_core_144;
  wire popcount33_fozj_core_145;
  wire popcount33_fozj_core_146;
  wire popcount33_fozj_core_149;
  wire popcount33_fozj_core_151;
  wire popcount33_fozj_core_152;
  wire popcount33_fozj_core_153;
  wire popcount33_fozj_core_156;
  wire popcount33_fozj_core_157;
  wire popcount33_fozj_core_158;
  wire popcount33_fozj_core_159;
  wire popcount33_fozj_core_160;
  wire popcount33_fozj_core_161;
  wire popcount33_fozj_core_162;
  wire popcount33_fozj_core_163;
  wire popcount33_fozj_core_164;
  wire popcount33_fozj_core_165;
  wire popcount33_fozj_core_167;
  wire popcount33_fozj_core_168;
  wire popcount33_fozj_core_169;
  wire popcount33_fozj_core_171;
  wire popcount33_fozj_core_172;
  wire popcount33_fozj_core_173;
  wire popcount33_fozj_core_174;
  wire popcount33_fozj_core_175;
  wire popcount33_fozj_core_179;
  wire popcount33_fozj_core_180;
  wire popcount33_fozj_core_181;
  wire popcount33_fozj_core_182;
  wire popcount33_fozj_core_184;
  wire popcount33_fozj_core_185;
  wire popcount33_fozj_core_187;
  wire popcount33_fozj_core_188;
  wire popcount33_fozj_core_190;
  wire popcount33_fozj_core_191;
  wire popcount33_fozj_core_194;
  wire popcount33_fozj_core_195;
  wire popcount33_fozj_core_196;
  wire popcount33_fozj_core_197;
  wire popcount33_fozj_core_198;
  wire popcount33_fozj_core_200;
  wire popcount33_fozj_core_202;
  wire popcount33_fozj_core_203;
  wire popcount33_fozj_core_204;
  wire popcount33_fozj_core_206;
  wire popcount33_fozj_core_207;
  wire popcount33_fozj_core_208;
  wire popcount33_fozj_core_209;
  wire popcount33_fozj_core_210;
  wire popcount33_fozj_core_211;
  wire popcount33_fozj_core_212;
  wire popcount33_fozj_core_213;
  wire popcount33_fozj_core_218;
  wire popcount33_fozj_core_219;
  wire popcount33_fozj_core_221;
  wire popcount33_fozj_core_223;
  wire popcount33_fozj_core_225;
  wire popcount33_fozj_core_226;
  wire popcount33_fozj_core_227;
  wire popcount33_fozj_core_228;
  wire popcount33_fozj_core_229;
  wire popcount33_fozj_core_234;
  wire popcount33_fozj_core_235;
  wire popcount33_fozj_core_237;
  wire popcount33_fozj_core_238;

  assign popcount33_fozj_core_035 = input_a[25] & input_a[29];
  assign popcount33_fozj_core_036 = input_a[28] | input_a[8];
  assign popcount33_fozj_core_037 = input_a[6] ^ input_a[20];
  assign popcount33_fozj_core_038 = ~(input_a[19] & input_a[30]);
  assign popcount33_fozj_core_040 = ~input_a[6];
  assign popcount33_fozj_core_041 = input_a[20] | input_a[8];
  assign popcount33_fozj_core_044 = input_a[22] ^ input_a[6];
  assign popcount33_fozj_core_045 = ~(input_a[32] & input_a[22]);
  assign popcount33_fozj_core_048 = ~input_a[8];
  assign popcount33_fozj_core_049_not = ~input_a[29];
  assign popcount33_fozj_core_050 = ~(input_a[30] ^ input_a[11]);
  assign popcount33_fozj_core_051 = ~(input_a[9] | input_a[21]);
  assign popcount33_fozj_core_053 = ~input_a[15];
  assign popcount33_fozj_core_054 = ~(input_a[3] & input_a[18]);
  assign popcount33_fozj_core_055 = input_a[21] & input_a[10];
  assign popcount33_fozj_core_056 = ~(input_a[23] | input_a[18]);
  assign popcount33_fozj_core_059 = input_a[3] ^ input_a[2];
  assign popcount33_fozj_core_060 = input_a[25] & input_a[30];
  assign popcount33_fozj_core_062 = ~(input_a[27] ^ input_a[17]);
  assign popcount33_fozj_core_063 = input_a[29] ^ input_a[14];
  assign popcount33_fozj_core_064 = ~(input_a[32] | input_a[26]);
  assign popcount33_fozj_core_065_not = ~input_a[11];
  assign popcount33_fozj_core_066 = ~(input_a[1] | input_a[16]);
  assign popcount33_fozj_core_067 = ~(input_a[7] & input_a[12]);
  assign popcount33_fozj_core_068 = input_a[3] | input_a[10];
  assign popcount33_fozj_core_074 = input_a[18] ^ input_a[25];
  assign popcount33_fozj_core_075 = input_a[14] ^ input_a[21];
  assign popcount33_fozj_core_079 = ~(input_a[3] | input_a[5]);
  assign popcount33_fozj_core_080 = ~(input_a[31] ^ input_a[19]);
  assign popcount33_fozj_core_081 = input_a[15] ^ input_a[6];
  assign popcount33_fozj_core_082 = ~(input_a[18] ^ input_a[25]);
  assign popcount33_fozj_core_083 = ~(input_a[31] ^ input_a[8]);
  assign popcount33_fozj_core_084 = ~(input_a[30] & input_a[3]);
  assign popcount33_fozj_core_085_not = ~input_a[19];
  assign popcount33_fozj_core_087 = input_a[12] & input_a[29];
  assign popcount33_fozj_core_090 = input_a[28] & input_a[14];
  assign popcount33_fozj_core_091 = input_a[27] & input_a[31];
  assign popcount33_fozj_core_092 = ~(input_a[0] & input_a[29]);
  assign popcount33_fozj_core_093 = ~input_a[13];
  assign popcount33_fozj_core_096 = input_a[27] ^ input_a[17];
  assign popcount33_fozj_core_101 = ~input_a[9];
  assign popcount33_fozj_core_102 = input_a[32] | input_a[16];
  assign popcount33_fozj_core_104_not = ~input_a[7];
  assign popcount33_fozj_core_105 = ~(input_a[26] | input_a[13]);
  assign popcount33_fozj_core_107 = input_a[4] | input_a[8];
  assign popcount33_fozj_core_108 = ~input_a[9];
  assign popcount33_fozj_core_110 = input_a[9] ^ input_a[26];
  assign popcount33_fozj_core_111 = input_a[3] ^ input_a[5];
  assign popcount33_fozj_core_112 = ~(input_a[22] | input_a[7]);
  assign popcount33_fozj_core_113 = ~(input_a[16] | input_a[21]);
  assign popcount33_fozj_core_114 = input_a[3] ^ input_a[8];
  assign popcount33_fozj_core_115 = input_a[19] | input_a[4];
  assign popcount33_fozj_core_116 = input_a[17] | input_a[24];
  assign popcount33_fozj_core_117 = input_a[19] ^ input_a[29];
  assign popcount33_fozj_core_121 = input_a[23] & input_a[24];
  assign popcount33_fozj_core_122 = ~input_a[26];
  assign popcount33_fozj_core_123 = ~(input_a[9] | input_a[3]);
  assign popcount33_fozj_core_124 = ~(input_a[29] | input_a[9]);
  assign popcount33_fozj_core_125 = input_a[32] ^ input_a[29];
  assign popcount33_fozj_core_126 = input_a[26] ^ input_a[3];
  assign popcount33_fozj_core_130 = input_a[19] | input_a[6];
  assign popcount33_fozj_core_133 = ~(input_a[3] & input_a[13]);
  assign popcount33_fozj_core_134 = input_a[5] & input_a[26];
  assign popcount33_fozj_core_137 = input_a[24] & input_a[27];
  assign popcount33_fozj_core_139 = input_a[23] ^ input_a[15];
  assign popcount33_fozj_core_140 = ~input_a[23];
  assign popcount33_fozj_core_142 = ~(input_a[9] | input_a[15]);
  assign popcount33_fozj_core_144 = input_a[4] ^ input_a[3];
  assign popcount33_fozj_core_145 = ~(input_a[19] & input_a[17]);
  assign popcount33_fozj_core_146 = ~input_a[1];
  assign popcount33_fozj_core_149 = ~(input_a[6] & input_a[29]);
  assign popcount33_fozj_core_151 = input_a[8] & input_a[21];
  assign popcount33_fozj_core_152 = input_a[20] ^ input_a[26];
  assign popcount33_fozj_core_153 = ~input_a[22];
  assign popcount33_fozj_core_156 = input_a[10] ^ input_a[32];
  assign popcount33_fozj_core_157 = input_a[25] & input_a[10];
  assign popcount33_fozj_core_158 = input_a[8] | input_a[25];
  assign popcount33_fozj_core_159 = ~input_a[2];
  assign popcount33_fozj_core_160 = input_a[15] & input_a[10];
  assign popcount33_fozj_core_161 = input_a[0] ^ input_a[16];
  assign popcount33_fozj_core_162 = input_a[19] & input_a[21];
  assign popcount33_fozj_core_163 = ~input_a[10];
  assign popcount33_fozj_core_164 = input_a[30] | input_a[25];
  assign popcount33_fozj_core_165 = ~(input_a[29] & input_a[12]);
  assign popcount33_fozj_core_167 = input_a[22] | input_a[26];
  assign popcount33_fozj_core_168 = input_a[18] ^ input_a[7];
  assign popcount33_fozj_core_169 = ~input_a[31];
  assign popcount33_fozj_core_171 = input_a[21] | input_a[0];
  assign popcount33_fozj_core_172 = input_a[4] | input_a[25];
  assign popcount33_fozj_core_173 = ~(input_a[30] ^ input_a[5]);
  assign popcount33_fozj_core_174 = input_a[18] ^ input_a[32];
  assign popcount33_fozj_core_175 = ~(input_a[2] ^ input_a[9]);
  assign popcount33_fozj_core_179 = input_a[19] ^ input_a[15];
  assign popcount33_fozj_core_180 = ~input_a[1];
  assign popcount33_fozj_core_181 = input_a[16] & input_a[0];
  assign popcount33_fozj_core_182 = ~(input_a[0] & input_a[20]);
  assign popcount33_fozj_core_184 = ~(input_a[3] ^ input_a[8]);
  assign popcount33_fozj_core_185 = input_a[20] & input_a[31];
  assign popcount33_fozj_core_187 = input_a[4] ^ input_a[1];
  assign popcount33_fozj_core_188 = ~(input_a[30] ^ input_a[2]);
  assign popcount33_fozj_core_190 = ~(input_a[20] | input_a[0]);
  assign popcount33_fozj_core_191 = ~(input_a[12] | input_a[0]);
  assign popcount33_fozj_core_194 = input_a[20] & input_a[8];
  assign popcount33_fozj_core_195 = ~(input_a[11] & input_a[18]);
  assign popcount33_fozj_core_196 = ~(input_a[3] & input_a[13]);
  assign popcount33_fozj_core_197 = ~input_a[13];
  assign popcount33_fozj_core_198 = ~input_a[29];
  assign popcount33_fozj_core_200 = ~(input_a[31] & input_a[3]);
  assign popcount33_fozj_core_202 = input_a[18] & input_a[2];
  assign popcount33_fozj_core_203 = input_a[17] ^ input_a[24];
  assign popcount33_fozj_core_204 = input_a[25] ^ input_a[29];
  assign popcount33_fozj_core_206 = ~(input_a[17] & input_a[27]);
  assign popcount33_fozj_core_207 = input_a[6] | input_a[4];
  assign popcount33_fozj_core_208 = input_a[10] & input_a[9];
  assign popcount33_fozj_core_209 = input_a[5] ^ input_a[25];
  assign popcount33_fozj_core_210 = input_a[10] & input_a[24];
  assign popcount33_fozj_core_211 = ~(input_a[25] & input_a[19]);
  assign popcount33_fozj_core_212 = input_a[0] & input_a[23];
  assign popcount33_fozj_core_213 = input_a[1] ^ input_a[17];
  assign popcount33_fozj_core_218 = ~(input_a[26] ^ input_a[25]);
  assign popcount33_fozj_core_219 = ~(input_a[19] ^ input_a[8]);
  assign popcount33_fozj_core_221 = ~(input_a[21] ^ input_a[7]);
  assign popcount33_fozj_core_223 = ~(input_a[30] ^ input_a[16]);
  assign popcount33_fozj_core_225 = ~(input_a[3] | input_a[12]);
  assign popcount33_fozj_core_226 = ~(input_a[0] | input_a[11]);
  assign popcount33_fozj_core_227 = ~(input_a[27] & input_a[8]);
  assign popcount33_fozj_core_228 = input_a[24] & input_a[10];
  assign popcount33_fozj_core_229 = ~input_a[13];
  assign popcount33_fozj_core_234 = ~(input_a[9] | input_a[15]);
  assign popcount33_fozj_core_235 = input_a[14] & input_a[12];
  assign popcount33_fozj_core_237 = input_a[26] ^ input_a[22];
  assign popcount33_fozj_core_238 = input_a[28] | input_a[32];

  assign popcount33_fozj_out[0] = 1'b0;
  assign popcount33_fozj_out[1] = input_a[21];
  assign popcount33_fozj_out[2] = input_a[32];
  assign popcount33_fozj_out[3] = 1'b0;
  assign popcount33_fozj_out[4] = 1'b1;
  assign popcount33_fozj_out[5] = 1'b0;
endmodule