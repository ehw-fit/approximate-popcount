// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.57029
// WCE=27.0
// EP=0.980915%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount34_gs0l(input [33:0] input_a, output [5:0] popcount34_gs0l_out);
  wire popcount34_gs0l_core_036;
  wire popcount34_gs0l_core_039_not;
  wire popcount34_gs0l_core_041;
  wire popcount34_gs0l_core_043;
  wire popcount34_gs0l_core_044;
  wire popcount34_gs0l_core_046;
  wire popcount34_gs0l_core_047;
  wire popcount34_gs0l_core_048;
  wire popcount34_gs0l_core_050;
  wire popcount34_gs0l_core_051;
  wire popcount34_gs0l_core_053;
  wire popcount34_gs0l_core_054;
  wire popcount34_gs0l_core_057;
  wire popcount34_gs0l_core_061;
  wire popcount34_gs0l_core_066;
  wire popcount34_gs0l_core_067;
  wire popcount34_gs0l_core_069;
  wire popcount34_gs0l_core_070;
  wire popcount34_gs0l_core_071;
  wire popcount34_gs0l_core_073;
  wire popcount34_gs0l_core_074;
  wire popcount34_gs0l_core_075;
  wire popcount34_gs0l_core_077;
  wire popcount34_gs0l_core_079;
  wire popcount34_gs0l_core_080;
  wire popcount34_gs0l_core_085;
  wire popcount34_gs0l_core_087;
  wire popcount34_gs0l_core_088;
  wire popcount34_gs0l_core_089;
  wire popcount34_gs0l_core_091;
  wire popcount34_gs0l_core_092;
  wire popcount34_gs0l_core_095;
  wire popcount34_gs0l_core_097;
  wire popcount34_gs0l_core_099;
  wire popcount34_gs0l_core_104;
  wire popcount34_gs0l_core_105;
  wire popcount34_gs0l_core_109_not;
  wire popcount34_gs0l_core_110;
  wire popcount34_gs0l_core_111;
  wire popcount34_gs0l_core_112;
  wire popcount34_gs0l_core_113;
  wire popcount34_gs0l_core_114;
  wire popcount34_gs0l_core_115;
  wire popcount34_gs0l_core_116_not;
  wire popcount34_gs0l_core_117;
  wire popcount34_gs0l_core_118;
  wire popcount34_gs0l_core_120;
  wire popcount34_gs0l_core_121;
  wire popcount34_gs0l_core_122;
  wire popcount34_gs0l_core_123;
  wire popcount34_gs0l_core_126;
  wire popcount34_gs0l_core_129_not;
  wire popcount34_gs0l_core_131;
  wire popcount34_gs0l_core_134;
  wire popcount34_gs0l_core_135;
  wire popcount34_gs0l_core_136;
  wire popcount34_gs0l_core_139;
  wire popcount34_gs0l_core_143;
  wire popcount34_gs0l_core_145;
  wire popcount34_gs0l_core_149;
  wire popcount34_gs0l_core_150;
  wire popcount34_gs0l_core_151;
  wire popcount34_gs0l_core_152;
  wire popcount34_gs0l_core_155;
  wire popcount34_gs0l_core_156;
  wire popcount34_gs0l_core_158;
  wire popcount34_gs0l_core_161;
  wire popcount34_gs0l_core_162;
  wire popcount34_gs0l_core_164;
  wire popcount34_gs0l_core_167;
  wire popcount34_gs0l_core_168;
  wire popcount34_gs0l_core_169_not;
  wire popcount34_gs0l_core_170;
  wire popcount34_gs0l_core_171;
  wire popcount34_gs0l_core_172;
  wire popcount34_gs0l_core_174;
  wire popcount34_gs0l_core_175;
  wire popcount34_gs0l_core_177;
  wire popcount34_gs0l_core_179;
  wire popcount34_gs0l_core_180;
  wire popcount34_gs0l_core_181;
  wire popcount34_gs0l_core_183;
  wire popcount34_gs0l_core_184;
  wire popcount34_gs0l_core_185;
  wire popcount34_gs0l_core_186;
  wire popcount34_gs0l_core_187;
  wire popcount34_gs0l_core_189;
  wire popcount34_gs0l_core_190;
  wire popcount34_gs0l_core_191;
  wire popcount34_gs0l_core_192;
  wire popcount34_gs0l_core_194;
  wire popcount34_gs0l_core_195;
  wire popcount34_gs0l_core_196;
  wire popcount34_gs0l_core_198;
  wire popcount34_gs0l_core_199;
  wire popcount34_gs0l_core_201;
  wire popcount34_gs0l_core_203;
  wire popcount34_gs0l_core_204;
  wire popcount34_gs0l_core_205;
  wire popcount34_gs0l_core_206;
  wire popcount34_gs0l_core_208;
  wire popcount34_gs0l_core_209;
  wire popcount34_gs0l_core_210;
  wire popcount34_gs0l_core_212;
  wire popcount34_gs0l_core_213;
  wire popcount34_gs0l_core_214;
  wire popcount34_gs0l_core_215;
  wire popcount34_gs0l_core_219_not;
  wire popcount34_gs0l_core_226;
  wire popcount34_gs0l_core_229;
  wire popcount34_gs0l_core_230;
  wire popcount34_gs0l_core_231;
  wire popcount34_gs0l_core_232;
  wire popcount34_gs0l_core_234;
  wire popcount34_gs0l_core_235;
  wire popcount34_gs0l_core_239;
  wire popcount34_gs0l_core_242;
  wire popcount34_gs0l_core_243;
  wire popcount34_gs0l_core_244;
  wire popcount34_gs0l_core_245;
  wire popcount34_gs0l_core_246;
  wire popcount34_gs0l_core_247;
  wire popcount34_gs0l_core_248;
  wire popcount34_gs0l_core_249;
  wire popcount34_gs0l_core_250;
  wire popcount34_gs0l_core_251;
  wire popcount34_gs0l_core_252;

  assign popcount34_gs0l_core_036 = input_a[12] ^ input_a[0];
  assign popcount34_gs0l_core_039_not = ~input_a[27];
  assign popcount34_gs0l_core_041 = ~(input_a[22] & input_a[1]);
  assign popcount34_gs0l_core_043 = input_a[1] & input_a[10];
  assign popcount34_gs0l_core_044 = input_a[23] & input_a[10];
  assign popcount34_gs0l_core_046 = ~(input_a[28] | input_a[20]);
  assign popcount34_gs0l_core_047 = input_a[23] & input_a[28];
  assign popcount34_gs0l_core_048 = ~(input_a[13] & input_a[21]);
  assign popcount34_gs0l_core_050 = input_a[19] | input_a[20];
  assign popcount34_gs0l_core_051 = ~input_a[3];
  assign popcount34_gs0l_core_053 = ~(input_a[0] & input_a[3]);
  assign popcount34_gs0l_core_054 = ~(input_a[24] | input_a[30]);
  assign popcount34_gs0l_core_057 = input_a[31] ^ input_a[8];
  assign popcount34_gs0l_core_061 = ~(input_a[27] & input_a[14]);
  assign popcount34_gs0l_core_066 = input_a[1] | input_a[31];
  assign popcount34_gs0l_core_067 = ~(input_a[12] & input_a[3]);
  assign popcount34_gs0l_core_069 = input_a[2] ^ input_a[20];
  assign popcount34_gs0l_core_070 = ~(input_a[4] ^ input_a[3]);
  assign popcount34_gs0l_core_071 = input_a[31] ^ input_a[3];
  assign popcount34_gs0l_core_073 = ~(input_a[2] & input_a[10]);
  assign popcount34_gs0l_core_074 = ~(input_a[22] ^ input_a[32]);
  assign popcount34_gs0l_core_075 = ~(input_a[2] | input_a[6]);
  assign popcount34_gs0l_core_077 = ~input_a[6];
  assign popcount34_gs0l_core_079 = ~(input_a[20] ^ input_a[14]);
  assign popcount34_gs0l_core_080 = ~(input_a[33] ^ input_a[13]);
  assign popcount34_gs0l_core_085 = input_a[7] | input_a[3];
  assign popcount34_gs0l_core_087 = ~(input_a[16] | input_a[11]);
  assign popcount34_gs0l_core_088 = input_a[26] ^ input_a[27];
  assign popcount34_gs0l_core_089 = input_a[18] ^ input_a[26];
  assign popcount34_gs0l_core_091 = ~(input_a[11] & input_a[5]);
  assign popcount34_gs0l_core_092 = input_a[0] & input_a[15];
  assign popcount34_gs0l_core_095 = input_a[29] ^ input_a[8];
  assign popcount34_gs0l_core_097 = input_a[19] & input_a[2];
  assign popcount34_gs0l_core_099 = ~(input_a[17] & input_a[24]);
  assign popcount34_gs0l_core_104 = ~(input_a[12] & input_a[14]);
  assign popcount34_gs0l_core_105 = ~(input_a[33] & input_a[8]);
  assign popcount34_gs0l_core_109_not = ~input_a[15];
  assign popcount34_gs0l_core_110 = ~(input_a[22] & input_a[27]);
  assign popcount34_gs0l_core_111 = ~(input_a[29] & input_a[28]);
  assign popcount34_gs0l_core_112 = ~(input_a[6] & input_a[28]);
  assign popcount34_gs0l_core_113 = ~(input_a[8] ^ input_a[31]);
  assign popcount34_gs0l_core_114 = ~input_a[24];
  assign popcount34_gs0l_core_115 = input_a[12] | input_a[14];
  assign popcount34_gs0l_core_116_not = ~input_a[11];
  assign popcount34_gs0l_core_117 = input_a[17] | input_a[31];
  assign popcount34_gs0l_core_118 = input_a[31] & input_a[16];
  assign popcount34_gs0l_core_120 = input_a[30] & input_a[22];
  assign popcount34_gs0l_core_121 = ~(input_a[21] | input_a[11]);
  assign popcount34_gs0l_core_122 = ~(input_a[10] & input_a[11]);
  assign popcount34_gs0l_core_123 = input_a[12] | input_a[10];
  assign popcount34_gs0l_core_126 = input_a[11] | input_a[2];
  assign popcount34_gs0l_core_129_not = ~input_a[11];
  assign popcount34_gs0l_core_131 = ~input_a[32];
  assign popcount34_gs0l_core_134 = input_a[29] ^ input_a[4];
  assign popcount34_gs0l_core_135 = ~input_a[25];
  assign popcount34_gs0l_core_136 = input_a[6] ^ input_a[3];
  assign popcount34_gs0l_core_139 = input_a[14] ^ input_a[11];
  assign popcount34_gs0l_core_143 = ~(input_a[15] | input_a[6]);
  assign popcount34_gs0l_core_145 = ~(input_a[7] | input_a[30]);
  assign popcount34_gs0l_core_149 = input_a[29] | input_a[4];
  assign popcount34_gs0l_core_150 = input_a[16] | input_a[2];
  assign popcount34_gs0l_core_151 = input_a[28] | input_a[31];
  assign popcount34_gs0l_core_152 = ~(input_a[29] & input_a[25]);
  assign popcount34_gs0l_core_155 = ~input_a[32];
  assign popcount34_gs0l_core_156 = ~input_a[0];
  assign popcount34_gs0l_core_158 = ~input_a[1];
  assign popcount34_gs0l_core_161 = ~(input_a[15] ^ input_a[15]);
  assign popcount34_gs0l_core_162 = ~(input_a[29] | input_a[8]);
  assign popcount34_gs0l_core_164 = input_a[18] | input_a[18];
  assign popcount34_gs0l_core_167 = input_a[21] ^ input_a[17];
  assign popcount34_gs0l_core_168 = input_a[28] ^ input_a[30];
  assign popcount34_gs0l_core_169_not = ~input_a[10];
  assign popcount34_gs0l_core_170 = input_a[1] ^ input_a[33];
  assign popcount34_gs0l_core_171 = input_a[2] ^ input_a[28];
  assign popcount34_gs0l_core_172 = input_a[27] ^ input_a[5];
  assign popcount34_gs0l_core_174 = ~(input_a[19] ^ input_a[19]);
  assign popcount34_gs0l_core_175 = ~input_a[3];
  assign popcount34_gs0l_core_177 = ~input_a[15];
  assign popcount34_gs0l_core_179 = ~input_a[25];
  assign popcount34_gs0l_core_180 = input_a[23] & input_a[22];
  assign popcount34_gs0l_core_181 = input_a[27] ^ input_a[11];
  assign popcount34_gs0l_core_183 = ~(input_a[22] ^ input_a[16]);
  assign popcount34_gs0l_core_184 = input_a[7] ^ input_a[23];
  assign popcount34_gs0l_core_185 = ~(input_a[12] ^ input_a[13]);
  assign popcount34_gs0l_core_186 = ~(input_a[12] ^ input_a[23]);
  assign popcount34_gs0l_core_187 = ~(input_a[26] ^ input_a[0]);
  assign popcount34_gs0l_core_189 = ~(input_a[16] | input_a[16]);
  assign popcount34_gs0l_core_190 = ~(input_a[22] ^ input_a[16]);
  assign popcount34_gs0l_core_191 = input_a[20] ^ input_a[22];
  assign popcount34_gs0l_core_192 = ~(input_a[18] ^ input_a[12]);
  assign popcount34_gs0l_core_194 = input_a[24] | input_a[22];
  assign popcount34_gs0l_core_195 = ~input_a[24];
  assign popcount34_gs0l_core_196 = ~(input_a[5] ^ input_a[17]);
  assign popcount34_gs0l_core_198 = ~(input_a[13] & input_a[21]);
  assign popcount34_gs0l_core_199 = ~(input_a[2] ^ input_a[11]);
  assign popcount34_gs0l_core_201 = input_a[28] & input_a[11];
  assign popcount34_gs0l_core_203 = ~(input_a[25] | input_a[5]);
  assign popcount34_gs0l_core_204 = ~(input_a[3] | input_a[27]);
  assign popcount34_gs0l_core_205 = ~(input_a[27] ^ input_a[29]);
  assign popcount34_gs0l_core_206 = ~input_a[4];
  assign popcount34_gs0l_core_208 = input_a[1] ^ input_a[11];
  assign popcount34_gs0l_core_209 = input_a[8] | input_a[1];
  assign popcount34_gs0l_core_210 = ~(input_a[3] | input_a[6]);
  assign popcount34_gs0l_core_212 = ~(input_a[27] | input_a[32]);
  assign popcount34_gs0l_core_213 = ~input_a[9];
  assign popcount34_gs0l_core_214 = input_a[31] & input_a[2];
  assign popcount34_gs0l_core_215 = input_a[23] ^ input_a[30];
  assign popcount34_gs0l_core_219_not = ~input_a[19];
  assign popcount34_gs0l_core_226 = input_a[4] & input_a[27];
  assign popcount34_gs0l_core_229 = input_a[28] | input_a[0];
  assign popcount34_gs0l_core_230 = ~(input_a[27] ^ input_a[15]);
  assign popcount34_gs0l_core_231 = ~(input_a[3] ^ input_a[8]);
  assign popcount34_gs0l_core_232 = ~(input_a[22] & input_a[20]);
  assign popcount34_gs0l_core_234 = input_a[7] & input_a[22];
  assign popcount34_gs0l_core_235 = input_a[11] | input_a[25];
  assign popcount34_gs0l_core_239 = ~(input_a[13] ^ input_a[15]);
  assign popcount34_gs0l_core_242 = ~(input_a[23] | input_a[9]);
  assign popcount34_gs0l_core_243 = input_a[2] & input_a[23];
  assign popcount34_gs0l_core_244 = input_a[11] ^ input_a[2];
  assign popcount34_gs0l_core_245 = ~(input_a[30] & input_a[16]);
  assign popcount34_gs0l_core_246 = input_a[24] ^ input_a[20];
  assign popcount34_gs0l_core_247 = ~(input_a[22] ^ input_a[17]);
  assign popcount34_gs0l_core_248 = input_a[8] ^ input_a[13];
  assign popcount34_gs0l_core_249 = ~(input_a[33] ^ input_a[0]);
  assign popcount34_gs0l_core_250 = ~(input_a[25] ^ input_a[4]);
  assign popcount34_gs0l_core_251 = ~(input_a[10] | input_a[31]);
  assign popcount34_gs0l_core_252 = ~input_a[2];

  assign popcount34_gs0l_out[0] = input_a[28];
  assign popcount34_gs0l_out[1] = input_a[26];
  assign popcount34_gs0l_out[2] = input_a[14];
  assign popcount34_gs0l_out[3] = 1'b1;
  assign popcount34_gs0l_out[4] = input_a[25];
  assign popcount34_gs0l_out[5] = 1'b0;
endmodule