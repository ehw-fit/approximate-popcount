// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.80263
// WCE=28.0
// EP=0.964362%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_lwvc(input [27:0] input_a, output [4:0] popcount28_lwvc_out);
  wire popcount28_lwvc_core_031;
  wire popcount28_lwvc_core_033;
  wire popcount28_lwvc_core_035;
  wire popcount28_lwvc_core_036;
  wire popcount28_lwvc_core_037;
  wire popcount28_lwvc_core_039;
  wire popcount28_lwvc_core_040;
  wire popcount28_lwvc_core_041;
  wire popcount28_lwvc_core_044;
  wire popcount28_lwvc_core_047;
  wire popcount28_lwvc_core_048;
  wire popcount28_lwvc_core_049;
  wire popcount28_lwvc_core_050;
  wire popcount28_lwvc_core_051;
  wire popcount28_lwvc_core_052;
  wire popcount28_lwvc_core_053_not;
  wire popcount28_lwvc_core_055;
  wire popcount28_lwvc_core_057;
  wire popcount28_lwvc_core_058;
  wire popcount28_lwvc_core_060;
  wire popcount28_lwvc_core_063;
  wire popcount28_lwvc_core_064;
  wire popcount28_lwvc_core_065;
  wire popcount28_lwvc_core_066;
  wire popcount28_lwvc_core_068;
  wire popcount28_lwvc_core_069;
  wire popcount28_lwvc_core_070;
  wire popcount28_lwvc_core_072;
  wire popcount28_lwvc_core_077;
  wire popcount28_lwvc_core_080;
  wire popcount28_lwvc_core_082;
  wire popcount28_lwvc_core_085;
  wire popcount28_lwvc_core_087;
  wire popcount28_lwvc_core_089;
  wire popcount28_lwvc_core_090;
  wire popcount28_lwvc_core_091;
  wire popcount28_lwvc_core_094;
  wire popcount28_lwvc_core_095;
  wire popcount28_lwvc_core_096;
  wire popcount28_lwvc_core_097;
  wire popcount28_lwvc_core_098;
  wire popcount28_lwvc_core_099;
  wire popcount28_lwvc_core_100;
  wire popcount28_lwvc_core_101;
  wire popcount28_lwvc_core_102;
  wire popcount28_lwvc_core_104;
  wire popcount28_lwvc_core_105;
  wire popcount28_lwvc_core_106;
  wire popcount28_lwvc_core_107;
  wire popcount28_lwvc_core_108;
  wire popcount28_lwvc_core_109;
  wire popcount28_lwvc_core_110;
  wire popcount28_lwvc_core_111;
  wire popcount28_lwvc_core_113;
  wire popcount28_lwvc_core_115;
  wire popcount28_lwvc_core_117;
  wire popcount28_lwvc_core_120;
  wire popcount28_lwvc_core_121;
  wire popcount28_lwvc_core_122;
  wire popcount28_lwvc_core_123;
  wire popcount28_lwvc_core_124;
  wire popcount28_lwvc_core_127;
  wire popcount28_lwvc_core_128;
  wire popcount28_lwvc_core_130;
  wire popcount28_lwvc_core_132;
  wire popcount28_lwvc_core_135;
  wire popcount28_lwvc_core_136;
  wire popcount28_lwvc_core_139;
  wire popcount28_lwvc_core_140;
  wire popcount28_lwvc_core_142;
  wire popcount28_lwvc_core_143;
  wire popcount28_lwvc_core_144;
  wire popcount28_lwvc_core_145;
  wire popcount28_lwvc_core_147;
  wire popcount28_lwvc_core_148_not;
  wire popcount28_lwvc_core_151;
  wire popcount28_lwvc_core_153;
  wire popcount28_lwvc_core_154;
  wire popcount28_lwvc_core_157;
  wire popcount28_lwvc_core_158;
  wire popcount28_lwvc_core_163;
  wire popcount28_lwvc_core_165;
  wire popcount28_lwvc_core_166;
  wire popcount28_lwvc_core_168;
  wire popcount28_lwvc_core_170;
  wire popcount28_lwvc_core_171;
  wire popcount28_lwvc_core_173;
  wire popcount28_lwvc_core_174;
  wire popcount28_lwvc_core_175_not;
  wire popcount28_lwvc_core_177;
  wire popcount28_lwvc_core_179;
  wire popcount28_lwvc_core_183;
  wire popcount28_lwvc_core_188_not;
  wire popcount28_lwvc_core_189;
  wire popcount28_lwvc_core_190;
  wire popcount28_lwvc_core_195;
  wire popcount28_lwvc_core_197;
  wire popcount28_lwvc_core_201;

  assign popcount28_lwvc_core_031 = input_a[2] ^ input_a[15];
  assign popcount28_lwvc_core_033 = input_a[7] ^ input_a[9];
  assign popcount28_lwvc_core_035 = ~input_a[27];
  assign popcount28_lwvc_core_036 = input_a[6] ^ input_a[2];
  assign popcount28_lwvc_core_037 = ~(input_a[8] | input_a[9]);
  assign popcount28_lwvc_core_039 = input_a[2] & input_a[16];
  assign popcount28_lwvc_core_040 = ~(input_a[20] | input_a[14]);
  assign popcount28_lwvc_core_041 = ~(input_a[7] ^ input_a[15]);
  assign popcount28_lwvc_core_044 = ~(input_a[5] & input_a[14]);
  assign popcount28_lwvc_core_047 = input_a[18] | input_a[15];
  assign popcount28_lwvc_core_048 = input_a[6] ^ input_a[12];
  assign popcount28_lwvc_core_049 = input_a[5] | input_a[9];
  assign popcount28_lwvc_core_050 = ~(input_a[16] ^ input_a[5]);
  assign popcount28_lwvc_core_051 = ~(input_a[8] & input_a[14]);
  assign popcount28_lwvc_core_052 = ~(input_a[9] | input_a[17]);
  assign popcount28_lwvc_core_053_not = ~input_a[12];
  assign popcount28_lwvc_core_055 = input_a[13] | input_a[2];
  assign popcount28_lwvc_core_057 = ~(input_a[10] ^ input_a[8]);
  assign popcount28_lwvc_core_058 = ~(input_a[16] | input_a[18]);
  assign popcount28_lwvc_core_060 = ~(input_a[21] | input_a[16]);
  assign popcount28_lwvc_core_063 = input_a[8] ^ input_a[12];
  assign popcount28_lwvc_core_064 = ~(input_a[7] ^ input_a[20]);
  assign popcount28_lwvc_core_065 = input_a[12] | input_a[10];
  assign popcount28_lwvc_core_066 = ~input_a[27];
  assign popcount28_lwvc_core_068 = ~(input_a[4] & input_a[23]);
  assign popcount28_lwvc_core_069 = ~(input_a[15] & input_a[15]);
  assign popcount28_lwvc_core_070 = ~(input_a[1] & input_a[15]);
  assign popcount28_lwvc_core_072 = ~(input_a[4] | input_a[21]);
  assign popcount28_lwvc_core_077 = ~(input_a[25] & input_a[10]);
  assign popcount28_lwvc_core_080 = input_a[3] ^ input_a[21];
  assign popcount28_lwvc_core_082 = input_a[27] ^ input_a[13];
  assign popcount28_lwvc_core_085 = input_a[12] & input_a[19];
  assign popcount28_lwvc_core_087 = input_a[23] | input_a[25];
  assign popcount28_lwvc_core_089 = ~(input_a[18] & input_a[20]);
  assign popcount28_lwvc_core_090 = input_a[24] & input_a[10];
  assign popcount28_lwvc_core_091 = ~(input_a[13] & input_a[5]);
  assign popcount28_lwvc_core_094 = ~(input_a[19] ^ input_a[27]);
  assign popcount28_lwvc_core_095 = ~(input_a[11] ^ input_a[23]);
  assign popcount28_lwvc_core_096 = input_a[0] | input_a[18];
  assign popcount28_lwvc_core_097 = ~(input_a[16] | input_a[3]);
  assign popcount28_lwvc_core_098 = input_a[10] | input_a[14];
  assign popcount28_lwvc_core_099 = ~input_a[23];
  assign popcount28_lwvc_core_100 = ~(input_a[8] ^ input_a[6]);
  assign popcount28_lwvc_core_101 = input_a[19] ^ input_a[5];
  assign popcount28_lwvc_core_102 = ~input_a[25];
  assign popcount28_lwvc_core_104 = ~input_a[0];
  assign popcount28_lwvc_core_105 = ~input_a[7];
  assign popcount28_lwvc_core_106 = ~(input_a[21] ^ input_a[23]);
  assign popcount28_lwvc_core_107 = input_a[27] ^ input_a[8];
  assign popcount28_lwvc_core_108 = input_a[19] & input_a[12];
  assign popcount28_lwvc_core_109 = input_a[9] & input_a[15];
  assign popcount28_lwvc_core_110 = input_a[12] & input_a[5];
  assign popcount28_lwvc_core_111 = ~(input_a[14] & input_a[4]);
  assign popcount28_lwvc_core_113 = ~input_a[27];
  assign popcount28_lwvc_core_115 = input_a[23] & input_a[14];
  assign popcount28_lwvc_core_117 = input_a[15] | input_a[7];
  assign popcount28_lwvc_core_120 = input_a[1] | input_a[18];
  assign popcount28_lwvc_core_121 = ~(input_a[9] ^ input_a[20]);
  assign popcount28_lwvc_core_122 = ~(input_a[14] & input_a[16]);
  assign popcount28_lwvc_core_123 = input_a[10] | input_a[20];
  assign popcount28_lwvc_core_124 = input_a[10] ^ input_a[1];
  assign popcount28_lwvc_core_127 = input_a[2] & input_a[17];
  assign popcount28_lwvc_core_128 = ~(input_a[22] & input_a[15]);
  assign popcount28_lwvc_core_130 = ~input_a[1];
  assign popcount28_lwvc_core_132 = ~input_a[16];
  assign popcount28_lwvc_core_135 = ~input_a[14];
  assign popcount28_lwvc_core_136 = ~(input_a[7] ^ input_a[19]);
  assign popcount28_lwvc_core_139 = input_a[17] ^ input_a[3];
  assign popcount28_lwvc_core_140 = ~(input_a[20] ^ input_a[0]);
  assign popcount28_lwvc_core_142 = ~(input_a[12] ^ input_a[8]);
  assign popcount28_lwvc_core_143 = ~(input_a[1] & input_a[23]);
  assign popcount28_lwvc_core_144 = ~(input_a[25] & input_a[20]);
  assign popcount28_lwvc_core_145 = ~input_a[2];
  assign popcount28_lwvc_core_147 = input_a[2] & input_a[24];
  assign popcount28_lwvc_core_148_not = ~input_a[0];
  assign popcount28_lwvc_core_151 = ~input_a[6];
  assign popcount28_lwvc_core_153 = input_a[16] & input_a[3];
  assign popcount28_lwvc_core_154 = ~(input_a[21] & input_a[26]);
  assign popcount28_lwvc_core_157 = ~(input_a[27] ^ input_a[0]);
  assign popcount28_lwvc_core_158 = input_a[20] & input_a[2];
  assign popcount28_lwvc_core_163 = ~(input_a[11] | input_a[16]);
  assign popcount28_lwvc_core_165 = input_a[10] ^ input_a[13];
  assign popcount28_lwvc_core_166 = ~input_a[26];
  assign popcount28_lwvc_core_168 = input_a[20] ^ input_a[20];
  assign popcount28_lwvc_core_170 = ~(input_a[21] & input_a[27]);
  assign popcount28_lwvc_core_171 = ~input_a[5];
  assign popcount28_lwvc_core_173 = ~(input_a[7] | input_a[22]);
  assign popcount28_lwvc_core_174 = input_a[27] | input_a[22];
  assign popcount28_lwvc_core_175_not = ~input_a[9];
  assign popcount28_lwvc_core_177 = ~(input_a[20] ^ input_a[10]);
  assign popcount28_lwvc_core_179 = ~(input_a[4] ^ input_a[3]);
  assign popcount28_lwvc_core_183 = ~(input_a[8] | input_a[6]);
  assign popcount28_lwvc_core_188_not = ~input_a[10];
  assign popcount28_lwvc_core_189 = ~(input_a[9] & input_a[25]);
  assign popcount28_lwvc_core_190 = ~(input_a[24] ^ input_a[11]);
  assign popcount28_lwvc_core_195 = ~(input_a[23] | input_a[0]);
  assign popcount28_lwvc_core_197 = input_a[18] ^ input_a[18];
  assign popcount28_lwvc_core_201 = ~(input_a[4] & input_a[1]);

  assign popcount28_lwvc_out[0] = 1'b1;
  assign popcount28_lwvc_out[1] = input_a[14];
  assign popcount28_lwvc_out[2] = input_a[2];
  assign popcount28_lwvc_out[3] = 1'b1;
  assign popcount28_lwvc_out[4] = input_a[17];
endmodule