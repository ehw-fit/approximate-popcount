// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.49501
// WCE=11.0
// EP=0.790214%
// Printed PDK parameters:
//  Area=47984588.0
//  Delay=67266408.0
//  Power=2249400.0

module popcount30_u8tp(input [29:0] input_a, output [4:0] popcount30_u8tp_out);
  wire popcount30_u8tp_core_032;
  wire popcount30_u8tp_core_033;
  wire popcount30_u8tp_core_034;
  wire popcount30_u8tp_core_035;
  wire popcount30_u8tp_core_036;
  wire popcount30_u8tp_core_039;
  wire popcount30_u8tp_core_040;
  wire popcount30_u8tp_core_041;
  wire popcount30_u8tp_core_042;
  wire popcount30_u8tp_core_044;
  wire popcount30_u8tp_core_045;
  wire popcount30_u8tp_core_046;
  wire popcount30_u8tp_core_051;
  wire popcount30_u8tp_core_052;
  wire popcount30_u8tp_core_054;
  wire popcount30_u8tp_core_058;
  wire popcount30_u8tp_core_059;
  wire popcount30_u8tp_core_060;
  wire popcount30_u8tp_core_061;
  wire popcount30_u8tp_core_062;
  wire popcount30_u8tp_core_064;
  wire popcount30_u8tp_core_065;
  wire popcount30_u8tp_core_066;
  wire popcount30_u8tp_core_067;
  wire popcount30_u8tp_core_068;
  wire popcount30_u8tp_core_069;
  wire popcount30_u8tp_core_070;
  wire popcount30_u8tp_core_071;
  wire popcount30_u8tp_core_072;
  wire popcount30_u8tp_core_073;
  wire popcount30_u8tp_core_074;
  wire popcount30_u8tp_core_075;
  wire popcount30_u8tp_core_076;
  wire popcount30_u8tp_core_078;
  wire popcount30_u8tp_core_079;
  wire popcount30_u8tp_core_080;
  wire popcount30_u8tp_core_083;
  wire popcount30_u8tp_core_084;
  wire popcount30_u8tp_core_085;
  wire popcount30_u8tp_core_086;
  wire popcount30_u8tp_core_087;
  wire popcount30_u8tp_core_088;
  wire popcount30_u8tp_core_089;
  wire popcount30_u8tp_core_091;
  wire popcount30_u8tp_core_094;
  wire popcount30_u8tp_core_095_not;
  wire popcount30_u8tp_core_096;
  wire popcount30_u8tp_core_097;
  wire popcount30_u8tp_core_098;
  wire popcount30_u8tp_core_100;
  wire popcount30_u8tp_core_102;
  wire popcount30_u8tp_core_103;
  wire popcount30_u8tp_core_104;
  wire popcount30_u8tp_core_105;
  wire popcount30_u8tp_core_106;
  wire popcount30_u8tp_core_108;
  wire popcount30_u8tp_core_110;
  wire popcount30_u8tp_core_111;
  wire popcount30_u8tp_core_112;
  wire popcount30_u8tp_core_113;
  wire popcount30_u8tp_core_114;
  wire popcount30_u8tp_core_115;
  wire popcount30_u8tp_core_116;
  wire popcount30_u8tp_core_119;
  wire popcount30_u8tp_core_121;
  wire popcount30_u8tp_core_123;
  wire popcount30_u8tp_core_125;
  wire popcount30_u8tp_core_127_not;
  wire popcount30_u8tp_core_128;
  wire popcount30_u8tp_core_129;
  wire popcount30_u8tp_core_131;
  wire popcount30_u8tp_core_132;
  wire popcount30_u8tp_core_133;
  wire popcount30_u8tp_core_134;
  wire popcount30_u8tp_core_135;
  wire popcount30_u8tp_core_137;
  wire popcount30_u8tp_core_139;
  wire popcount30_u8tp_core_142;
  wire popcount30_u8tp_core_143;
  wire popcount30_u8tp_core_144;
  wire popcount30_u8tp_core_147;
  wire popcount30_u8tp_core_149;
  wire popcount30_u8tp_core_152;
  wire popcount30_u8tp_core_153;
  wire popcount30_u8tp_core_157;
  wire popcount30_u8tp_core_161;
  wire popcount30_u8tp_core_163;
  wire popcount30_u8tp_core_165;
  wire popcount30_u8tp_core_166;
  wire popcount30_u8tp_core_168;
  wire popcount30_u8tp_core_170;
  wire popcount30_u8tp_core_171;
  wire popcount30_u8tp_core_172;
  wire popcount30_u8tp_core_173;
  wire popcount30_u8tp_core_175;
  wire popcount30_u8tp_core_176;
  wire popcount30_u8tp_core_177;
  wire popcount30_u8tp_core_178;
  wire popcount30_u8tp_core_179;
  wire popcount30_u8tp_core_180;
  wire popcount30_u8tp_core_181;
  wire popcount30_u8tp_core_182;
  wire popcount30_u8tp_core_183;
  wire popcount30_u8tp_core_184;
  wire popcount30_u8tp_core_185;
  wire popcount30_u8tp_core_186;
  wire popcount30_u8tp_core_189;
  wire popcount30_u8tp_core_190;
  wire popcount30_u8tp_core_191;
  wire popcount30_u8tp_core_193;
  wire popcount30_u8tp_core_194;
  wire popcount30_u8tp_core_195;
  wire popcount30_u8tp_core_196;
  wire popcount30_u8tp_core_197;
  wire popcount30_u8tp_core_198;
  wire popcount30_u8tp_core_199;
  wire popcount30_u8tp_core_200;
  wire popcount30_u8tp_core_201;
  wire popcount30_u8tp_core_202;
  wire popcount30_u8tp_core_203;
  wire popcount30_u8tp_core_204;
  wire popcount30_u8tp_core_205;
  wire popcount30_u8tp_core_206;
  wire popcount30_u8tp_core_207;
  wire popcount30_u8tp_core_208;
  wire popcount30_u8tp_core_210;
  wire popcount30_u8tp_core_213_not;

  assign popcount30_u8tp_core_032 = input_a[1] | input_a[2];
  assign popcount30_u8tp_core_033 = input_a[1] & input_a[2];
  assign popcount30_u8tp_core_034 = ~input_a[29];
  assign popcount30_u8tp_core_035 = input_a[4] & popcount30_u8tp_core_032;
  assign popcount30_u8tp_core_036 = popcount30_u8tp_core_033 | popcount30_u8tp_core_035;
  assign popcount30_u8tp_core_039 = ~(input_a[29] ^ input_a[16]);
  assign popcount30_u8tp_core_040 = input_a[6] ^ input_a[3];
  assign popcount30_u8tp_core_041 = input_a[5] & input_a[6];
  assign popcount30_u8tp_core_042 = ~(input_a[28] | input_a[18]);
  assign popcount30_u8tp_core_044 = input_a[5] ^ input_a[3];
  assign popcount30_u8tp_core_045 = input_a[3] & popcount30_u8tp_core_041;
  assign popcount30_u8tp_core_046 = popcount30_u8tp_core_044 | popcount30_u8tp_core_040;
  assign popcount30_u8tp_core_051 = popcount30_u8tp_core_036 ^ popcount30_u8tp_core_046;
  assign popcount30_u8tp_core_052 = popcount30_u8tp_core_036 & popcount30_u8tp_core_046;
  assign popcount30_u8tp_core_054 = input_a[3] & input_a[26];
  assign popcount30_u8tp_core_058 = popcount30_u8tp_core_045 | popcount30_u8tp_core_052;
  assign popcount30_u8tp_core_059 = input_a[17] & input_a[10];
  assign popcount30_u8tp_core_060 = input_a[6] & input_a[28];
  assign popcount30_u8tp_core_061 = input_a[27] | input_a[4];
  assign popcount30_u8tp_core_062 = input_a[20] & input_a[9];
  assign popcount30_u8tp_core_064 = input_a[8] & input_a[10];
  assign popcount30_u8tp_core_065 = ~input_a[12];
  assign popcount30_u8tp_core_066 = input_a[11] & input_a[18];
  assign popcount30_u8tp_core_067 = popcount30_u8tp_core_062 | popcount30_u8tp_core_064;
  assign popcount30_u8tp_core_068 = ~(input_a[9] ^ input_a[23]);
  assign popcount30_u8tp_core_069 = popcount30_u8tp_core_067 | popcount30_u8tp_core_066;
  assign popcount30_u8tp_core_070 = ~(input_a[8] | input_a[20]);
  assign popcount30_u8tp_core_071 = ~input_a[5];
  assign popcount30_u8tp_core_072 = input_a[18] | input_a[12];
  assign popcount30_u8tp_core_073 = ~input_a[7];
  assign popcount30_u8tp_core_074 = ~(input_a[15] | input_a[1]);
  assign popcount30_u8tp_core_075 = ~(input_a[23] ^ input_a[4]);
  assign popcount30_u8tp_core_076 = input_a[15] | input_a[22];
  assign popcount30_u8tp_core_078 = ~(input_a[18] & input_a[0]);
  assign popcount30_u8tp_core_079 = input_a[21] | input_a[9];
  assign popcount30_u8tp_core_080 = input_a[11] | popcount30_u8tp_core_072;
  assign popcount30_u8tp_core_083 = input_a[17] | input_a[17];
  assign popcount30_u8tp_core_084 = input_a[14] & input_a[13];
  assign popcount30_u8tp_core_085 = popcount30_u8tp_core_069 ^ popcount30_u8tp_core_080;
  assign popcount30_u8tp_core_086 = popcount30_u8tp_core_069 & popcount30_u8tp_core_080;
  assign popcount30_u8tp_core_087 = popcount30_u8tp_core_085 ^ popcount30_u8tp_core_084;
  assign popcount30_u8tp_core_088 = popcount30_u8tp_core_085 & popcount30_u8tp_core_084;
  assign popcount30_u8tp_core_089 = popcount30_u8tp_core_086 | popcount30_u8tp_core_088;
  assign popcount30_u8tp_core_091 = ~input_a[12];
  assign popcount30_u8tp_core_094 = ~(input_a[21] | input_a[10]);
  assign popcount30_u8tp_core_095_not = ~input_a[14];
  assign popcount30_u8tp_core_096 = ~(input_a[9] ^ input_a[21]);
  assign popcount30_u8tp_core_097 = popcount30_u8tp_core_051 ^ popcount30_u8tp_core_087;
  assign popcount30_u8tp_core_098 = popcount30_u8tp_core_051 & popcount30_u8tp_core_087;
  assign popcount30_u8tp_core_100 = input_a[8] | input_a[21];
  assign popcount30_u8tp_core_102 = popcount30_u8tp_core_058 ^ popcount30_u8tp_core_089;
  assign popcount30_u8tp_core_103 = popcount30_u8tp_core_058 & popcount30_u8tp_core_089;
  assign popcount30_u8tp_core_104 = popcount30_u8tp_core_102 ^ popcount30_u8tp_core_098;
  assign popcount30_u8tp_core_105 = popcount30_u8tp_core_102 & popcount30_u8tp_core_098;
  assign popcount30_u8tp_core_106 = popcount30_u8tp_core_103 | popcount30_u8tp_core_105;
  assign popcount30_u8tp_core_108 = input_a[14] & input_a[26];
  assign popcount30_u8tp_core_110 = ~(input_a[16] ^ input_a[12]);
  assign popcount30_u8tp_core_111 = input_a[27] ^ input_a[29];
  assign popcount30_u8tp_core_112 = input_a[16] ^ input_a[17];
  assign popcount30_u8tp_core_113 = input_a[16] & input_a[17];
  assign popcount30_u8tp_core_114 = input_a[15] ^ popcount30_u8tp_core_112;
  assign popcount30_u8tp_core_115 = input_a[15] & popcount30_u8tp_core_112;
  assign popcount30_u8tp_core_116 = popcount30_u8tp_core_113 | popcount30_u8tp_core_115;
  assign popcount30_u8tp_core_119 = input_a[7] & input_a[21];
  assign popcount30_u8tp_core_121 = input_a[27] & input_a[0];
  assign popcount30_u8tp_core_123 = input_a[16] | input_a[20];
  assign popcount30_u8tp_core_125 = input_a[25] ^ input_a[6];
  assign popcount30_u8tp_core_127_not = ~input_a[25];
  assign popcount30_u8tp_core_128 = ~(input_a[18] | input_a[4]);
  assign popcount30_u8tp_core_129 = ~(input_a[13] ^ input_a[14]);
  assign popcount30_u8tp_core_131 = popcount30_u8tp_core_116 ^ popcount30_u8tp_core_119;
  assign popcount30_u8tp_core_132 = popcount30_u8tp_core_116 & popcount30_u8tp_core_119;
  assign popcount30_u8tp_core_133 = popcount30_u8tp_core_131 ^ popcount30_u8tp_core_114;
  assign popcount30_u8tp_core_134 = popcount30_u8tp_core_131 & popcount30_u8tp_core_114;
  assign popcount30_u8tp_core_135 = popcount30_u8tp_core_132 | popcount30_u8tp_core_134;
  assign popcount30_u8tp_core_137 = ~(input_a[20] & input_a[12]);
  assign popcount30_u8tp_core_139 = ~input_a[0];
  assign popcount30_u8tp_core_142 = input_a[22] & input_a[19];
  assign popcount30_u8tp_core_143 = ~(input_a[24] & input_a[25]);
  assign popcount30_u8tp_core_144 = input_a[24] & input_a[25];
  assign popcount30_u8tp_core_147 = popcount30_u8tp_core_142 ^ popcount30_u8tp_core_144;
  assign popcount30_u8tp_core_149 = popcount30_u8tp_core_147 ^ popcount30_u8tp_core_143;
  assign popcount30_u8tp_core_152 = ~(input_a[26] & input_a[27]);
  assign popcount30_u8tp_core_153 = input_a[26] & input_a[27];
  assign popcount30_u8tp_core_157 = popcount30_u8tp_core_152 & input_a[25];
  assign popcount30_u8tp_core_161 = ~(input_a[26] & input_a[19]);
  assign popcount30_u8tp_core_163 = input_a[28] | input_a[2];
  assign popcount30_u8tp_core_165 = popcount30_u8tp_core_149 ^ popcount30_u8tp_core_157;
  assign popcount30_u8tp_core_166 = input_a[25] & popcount30_u8tp_core_157;
  assign popcount30_u8tp_core_168 = input_a[20] ^ input_a[28];
  assign popcount30_u8tp_core_170 = popcount30_u8tp_core_142 ^ popcount30_u8tp_core_153;
  assign popcount30_u8tp_core_171 = popcount30_u8tp_core_142 & popcount30_u8tp_core_153;
  assign popcount30_u8tp_core_172 = popcount30_u8tp_core_170 | popcount30_u8tp_core_166;
  assign popcount30_u8tp_core_173 = input_a[19] | input_a[9];
  assign popcount30_u8tp_core_175 = ~(input_a[21] | input_a[14]);
  assign popcount30_u8tp_core_176 = input_a[0] & input_a[23];
  assign popcount30_u8tp_core_177 = popcount30_u8tp_core_133 ^ popcount30_u8tp_core_165;
  assign popcount30_u8tp_core_178 = popcount30_u8tp_core_133 & popcount30_u8tp_core_165;
  assign popcount30_u8tp_core_179 = popcount30_u8tp_core_177 ^ popcount30_u8tp_core_176;
  assign popcount30_u8tp_core_180 = popcount30_u8tp_core_177 & popcount30_u8tp_core_176;
  assign popcount30_u8tp_core_181 = popcount30_u8tp_core_178 | popcount30_u8tp_core_180;
  assign popcount30_u8tp_core_182 = popcount30_u8tp_core_135 ^ popcount30_u8tp_core_172;
  assign popcount30_u8tp_core_183 = popcount30_u8tp_core_135 & popcount30_u8tp_core_172;
  assign popcount30_u8tp_core_184 = popcount30_u8tp_core_182 ^ popcount30_u8tp_core_181;
  assign popcount30_u8tp_core_185 = popcount30_u8tp_core_182 & popcount30_u8tp_core_181;
  assign popcount30_u8tp_core_186 = popcount30_u8tp_core_183 | popcount30_u8tp_core_185;
  assign popcount30_u8tp_core_189 = popcount30_u8tp_core_171 | popcount30_u8tp_core_186;
  assign popcount30_u8tp_core_190 = input_a[26] & input_a[4];
  assign popcount30_u8tp_core_191 = ~input_a[27];
  assign popcount30_u8tp_core_193 = input_a[28] & input_a[24];
  assign popcount30_u8tp_core_194 = popcount30_u8tp_core_097 | popcount30_u8tp_core_179;
  assign popcount30_u8tp_core_195 = popcount30_u8tp_core_097 & popcount30_u8tp_core_179;
  assign popcount30_u8tp_core_196 = input_a[27] ^ input_a[14];
  assign popcount30_u8tp_core_197 = popcount30_u8tp_core_194 & popcount30_u8tp_core_193;
  assign popcount30_u8tp_core_198 = popcount30_u8tp_core_195 | popcount30_u8tp_core_197;
  assign popcount30_u8tp_core_199 = popcount30_u8tp_core_104 ^ popcount30_u8tp_core_184;
  assign popcount30_u8tp_core_200 = popcount30_u8tp_core_104 & popcount30_u8tp_core_184;
  assign popcount30_u8tp_core_201 = popcount30_u8tp_core_199 ^ popcount30_u8tp_core_198;
  assign popcount30_u8tp_core_202 = popcount30_u8tp_core_199 & popcount30_u8tp_core_198;
  assign popcount30_u8tp_core_203 = popcount30_u8tp_core_200 | popcount30_u8tp_core_202;
  assign popcount30_u8tp_core_204 = popcount30_u8tp_core_106 ^ popcount30_u8tp_core_189;
  assign popcount30_u8tp_core_205 = popcount30_u8tp_core_106 & popcount30_u8tp_core_189;
  assign popcount30_u8tp_core_206 = popcount30_u8tp_core_204 ^ popcount30_u8tp_core_203;
  assign popcount30_u8tp_core_207 = popcount30_u8tp_core_204 & popcount30_u8tp_core_203;
  assign popcount30_u8tp_core_208 = popcount30_u8tp_core_205 | popcount30_u8tp_core_207;
  assign popcount30_u8tp_core_210 = input_a[12] | input_a[17];
  assign popcount30_u8tp_core_213_not = ~input_a[26];

  assign popcount30_u8tp_out[0] = input_a[29];
  assign popcount30_u8tp_out[1] = popcount30_u8tp_core_206;
  assign popcount30_u8tp_out[2] = popcount30_u8tp_core_201;
  assign popcount30_u8tp_out[3] = popcount30_u8tp_core_206;
  assign popcount30_u8tp_out[4] = popcount30_u8tp_core_208;
endmodule