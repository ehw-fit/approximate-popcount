// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.44085
// WCE=17.0
// EP=0.934759%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount19_3csc(input [18:0] input_a, output [4:0] popcount19_3csc_out);
  wire popcount19_3csc_core_022;
  wire popcount19_3csc_core_023;
  wire popcount19_3csc_core_024;
  wire popcount19_3csc_core_025;
  wire popcount19_3csc_core_026;
  wire popcount19_3csc_core_027;
  wire popcount19_3csc_core_028;
  wire popcount19_3csc_core_029;
  wire popcount19_3csc_core_030;
  wire popcount19_3csc_core_033;
  wire popcount19_3csc_core_035;
  wire popcount19_3csc_core_036;
  wire popcount19_3csc_core_038;
  wire popcount19_3csc_core_039;
  wire popcount19_3csc_core_040;
  wire popcount19_3csc_core_041;
  wire popcount19_3csc_core_043;
  wire popcount19_3csc_core_044;
  wire popcount19_3csc_core_045;
  wire popcount19_3csc_core_046;
  wire popcount19_3csc_core_047;
  wire popcount19_3csc_core_050;
  wire popcount19_3csc_core_051;
  wire popcount19_3csc_core_052;
  wire popcount19_3csc_core_053;
  wire popcount19_3csc_core_057;
  wire popcount19_3csc_core_060;
  wire popcount19_3csc_core_062;
  wire popcount19_3csc_core_064;
  wire popcount19_3csc_core_066;
  wire popcount19_3csc_core_069;
  wire popcount19_3csc_core_070;
  wire popcount19_3csc_core_074;
  wire popcount19_3csc_core_076;
  wire popcount19_3csc_core_077;
  wire popcount19_3csc_core_078;
  wire popcount19_3csc_core_080;
  wire popcount19_3csc_core_081;
  wire popcount19_3csc_core_084;
  wire popcount19_3csc_core_085;
  wire popcount19_3csc_core_089;
  wire popcount19_3csc_core_093;
  wire popcount19_3csc_core_094;
  wire popcount19_3csc_core_095;
  wire popcount19_3csc_core_096;
  wire popcount19_3csc_core_097;
  wire popcount19_3csc_core_099;
  wire popcount19_3csc_core_101;
  wire popcount19_3csc_core_103;
  wire popcount19_3csc_core_104;
  wire popcount19_3csc_core_105;
  wire popcount19_3csc_core_106;
  wire popcount19_3csc_core_109;
  wire popcount19_3csc_core_111;
  wire popcount19_3csc_core_112;
  wire popcount19_3csc_core_114;
  wire popcount19_3csc_core_115;
  wire popcount19_3csc_core_116;
  wire popcount19_3csc_core_117;
  wire popcount19_3csc_core_118;
  wire popcount19_3csc_core_119;
  wire popcount19_3csc_core_120;
  wire popcount19_3csc_core_121;
  wire popcount19_3csc_core_122;
  wire popcount19_3csc_core_123;
  wire popcount19_3csc_core_124;
  wire popcount19_3csc_core_126_not;
  wire popcount19_3csc_core_127;
  wire popcount19_3csc_core_129;
  wire popcount19_3csc_core_130;
  wire popcount19_3csc_core_132;
  wire popcount19_3csc_core_135;

  assign popcount19_3csc_core_022 = ~input_a[13];
  assign popcount19_3csc_core_023 = input_a[16] & input_a[2];
  assign popcount19_3csc_core_024 = input_a[15] ^ input_a[2];
  assign popcount19_3csc_core_025 = ~input_a[0];
  assign popcount19_3csc_core_026 = ~input_a[2];
  assign popcount19_3csc_core_027 = input_a[11] ^ input_a[5];
  assign popcount19_3csc_core_028 = ~(input_a[17] & input_a[14]);
  assign popcount19_3csc_core_029 = ~input_a[10];
  assign popcount19_3csc_core_030 = ~(input_a[6] ^ input_a[9]);
  assign popcount19_3csc_core_033 = ~(input_a[1] & input_a[17]);
  assign popcount19_3csc_core_035 = ~(input_a[6] ^ input_a[16]);
  assign popcount19_3csc_core_036 = input_a[17] | input_a[6];
  assign popcount19_3csc_core_038 = ~(input_a[6] | input_a[17]);
  assign popcount19_3csc_core_039 = input_a[8] | input_a[14];
  assign popcount19_3csc_core_040 = input_a[11] & input_a[3];
  assign popcount19_3csc_core_041 = ~(input_a[9] | input_a[4]);
  assign popcount19_3csc_core_043 = ~(input_a[3] ^ input_a[3]);
  assign popcount19_3csc_core_044 = input_a[4] ^ input_a[10];
  assign popcount19_3csc_core_045 = input_a[18] | input_a[17];
  assign popcount19_3csc_core_046 = ~(input_a[12] & input_a[6]);
  assign popcount19_3csc_core_047 = ~(input_a[3] & input_a[7]);
  assign popcount19_3csc_core_050 = ~(input_a[17] ^ input_a[9]);
  assign popcount19_3csc_core_051 = input_a[7] | input_a[14];
  assign popcount19_3csc_core_052 = input_a[18] & input_a[13];
  assign popcount19_3csc_core_053 = ~(input_a[11] ^ input_a[12]);
  assign popcount19_3csc_core_057 = input_a[11] ^ input_a[2];
  assign popcount19_3csc_core_060 = input_a[13] ^ input_a[5];
  assign popcount19_3csc_core_062 = input_a[11] | input_a[8];
  assign popcount19_3csc_core_064 = input_a[0] ^ input_a[4];
  assign popcount19_3csc_core_066 = ~(input_a[7] & input_a[13]);
  assign popcount19_3csc_core_069 = ~(input_a[15] & input_a[16]);
  assign popcount19_3csc_core_070 = input_a[13] & input_a[2];
  assign popcount19_3csc_core_074 = ~(input_a[1] ^ input_a[14]);
  assign popcount19_3csc_core_076 = ~(input_a[3] | input_a[3]);
  assign popcount19_3csc_core_077 = input_a[14] ^ input_a[16];
  assign popcount19_3csc_core_078 = ~input_a[1];
  assign popcount19_3csc_core_080 = ~input_a[9];
  assign popcount19_3csc_core_081 = input_a[11] ^ input_a[2];
  assign popcount19_3csc_core_084 = ~(input_a[3] ^ input_a[7]);
  assign popcount19_3csc_core_085 = ~(input_a[14] | input_a[2]);
  assign popcount19_3csc_core_089 = input_a[18] & input_a[1];
  assign popcount19_3csc_core_093 = ~(input_a[17] & input_a[11]);
  assign popcount19_3csc_core_094 = ~(input_a[16] & input_a[16]);
  assign popcount19_3csc_core_095 = ~(input_a[16] ^ input_a[15]);
  assign popcount19_3csc_core_096 = ~(input_a[8] & input_a[12]);
  assign popcount19_3csc_core_097 = ~(input_a[10] & input_a[11]);
  assign popcount19_3csc_core_099 = input_a[12] & input_a[15];
  assign popcount19_3csc_core_101 = ~input_a[14];
  assign popcount19_3csc_core_103 = input_a[14] & input_a[18];
  assign popcount19_3csc_core_104 = ~(input_a[0] | input_a[1]);
  assign popcount19_3csc_core_105 = ~(input_a[13] | input_a[3]);
  assign popcount19_3csc_core_106 = ~input_a[0];
  assign popcount19_3csc_core_109 = ~(input_a[0] | input_a[11]);
  assign popcount19_3csc_core_111 = input_a[11] & input_a[4];
  assign popcount19_3csc_core_112 = ~input_a[14];
  assign popcount19_3csc_core_114 = ~(input_a[15] | input_a[16]);
  assign popcount19_3csc_core_115 = ~(input_a[12] ^ input_a[8]);
  assign popcount19_3csc_core_116 = input_a[17] & input_a[11];
  assign popcount19_3csc_core_117 = ~(input_a[16] ^ input_a[13]);
  assign popcount19_3csc_core_118 = input_a[13] & input_a[13];
  assign popcount19_3csc_core_119 = ~(input_a[1] ^ input_a[16]);
  assign popcount19_3csc_core_120 = ~input_a[3];
  assign popcount19_3csc_core_121 = ~(input_a[15] | input_a[16]);
  assign popcount19_3csc_core_122 = ~(input_a[14] & input_a[18]);
  assign popcount19_3csc_core_123 = input_a[2] & input_a[6];
  assign popcount19_3csc_core_124 = ~(input_a[10] & input_a[1]);
  assign popcount19_3csc_core_126_not = ~input_a[11];
  assign popcount19_3csc_core_127 = ~input_a[8];
  assign popcount19_3csc_core_129 = ~input_a[2];
  assign popcount19_3csc_core_130 = input_a[8] ^ input_a[15];
  assign popcount19_3csc_core_132 = input_a[10] | input_a[1];
  assign popcount19_3csc_core_135 = input_a[14] ^ input_a[17];

  assign popcount19_3csc_out[0] = input_a[10];
  assign popcount19_3csc_out[1] = input_a[10];
  assign popcount19_3csc_out[2] = input_a[10];
  assign popcount19_3csc_out[3] = input_a[4];
  assign popcount19_3csc_out[4] = 1'b0;
endmodule