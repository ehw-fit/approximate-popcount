// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.30531
// WCE=18.0
// EP=0.952966%
// Printed PDK parameters:
//  Area=55730658.0
//  Delay=83257816.0
//  Power=2068700.0

module popcount36_it2u(input [35:0] input_a, output [5:0] popcount36_it2u_out);
  wire popcount36_it2u_core_038;
  wire popcount36_it2u_core_039;
  wire popcount36_it2u_core_040;
  wire popcount36_it2u_core_042;
  wire popcount36_it2u_core_043;
  wire popcount36_it2u_core_044;
  wire popcount36_it2u_core_045;
  wire popcount36_it2u_core_046;
  wire popcount36_it2u_core_047;
  wire popcount36_it2u_core_049;
  wire popcount36_it2u_core_050;
  wire popcount36_it2u_core_051;
  wire popcount36_it2u_core_052;
  wire popcount36_it2u_core_053;
  wire popcount36_it2u_core_054;
  wire popcount36_it2u_core_055;
  wire popcount36_it2u_core_056;
  wire popcount36_it2u_core_057;
  wire popcount36_it2u_core_059;
  wire popcount36_it2u_core_060;
  wire popcount36_it2u_core_062;
  wire popcount36_it2u_core_064;
  wire popcount36_it2u_core_066;
  wire popcount36_it2u_core_067;
  wire popcount36_it2u_core_069;
  wire popcount36_it2u_core_079;
  wire popcount36_it2u_core_080;
  wire popcount36_it2u_core_081;
  wire popcount36_it2u_core_082;
  wire popcount36_it2u_core_083;
  wire popcount36_it2u_core_084;
  wire popcount36_it2u_core_085;
  wire popcount36_it2u_core_086;
  wire popcount36_it2u_core_087;
  wire popcount36_it2u_core_088;
  wire popcount36_it2u_core_091;
  wire popcount36_it2u_core_092;
  wire popcount36_it2u_core_093;
  wire popcount36_it2u_core_094;
  wire popcount36_it2u_core_095;
  wire popcount36_it2u_core_096;
  wire popcount36_it2u_core_097;
  wire popcount36_it2u_core_099;
  wire popcount36_it2u_core_100;
  wire popcount36_it2u_core_101;
  wire popcount36_it2u_core_102;
  wire popcount36_it2u_core_103;
  wire popcount36_it2u_core_104;
  wire popcount36_it2u_core_105;
  wire popcount36_it2u_core_109;
  wire popcount36_it2u_core_110;
  wire popcount36_it2u_core_111;
  wire popcount36_it2u_core_112;
  wire popcount36_it2u_core_113;
  wire popcount36_it2u_core_114;
  wire popcount36_it2u_core_115;
  wire popcount36_it2u_core_116;
  wire popcount36_it2u_core_117;
  wire popcount36_it2u_core_118;
  wire popcount36_it2u_core_119;
  wire popcount36_it2u_core_122;
  wire popcount36_it2u_core_123;
  wire popcount36_it2u_core_124;
  wire popcount36_it2u_core_125;
  wire popcount36_it2u_core_126;
  wire popcount36_it2u_core_127;
  wire popcount36_it2u_core_128;
  wire popcount36_it2u_core_131;
  wire popcount36_it2u_core_132;
  wire popcount36_it2u_core_134;
  wire popcount36_it2u_core_135;
  wire popcount36_it2u_core_136;
  wire popcount36_it2u_core_137;
  wire popcount36_it2u_core_138;
  wire popcount36_it2u_core_140;
  wire popcount36_it2u_core_142;
  wire popcount36_it2u_core_145;
  wire popcount36_it2u_core_147;
  wire popcount36_it2u_core_149;
  wire popcount36_it2u_core_150;
  wire popcount36_it2u_core_151;
  wire popcount36_it2u_core_155;
  wire popcount36_it2u_core_156;
  wire popcount36_it2u_core_157;
  wire popcount36_it2u_core_159;
  wire popcount36_it2u_core_160;
  wire popcount36_it2u_core_165;
  wire popcount36_it2u_core_166;
  wire popcount36_it2u_core_168;
  wire popcount36_it2u_core_174;
  wire popcount36_it2u_core_175;
  wire popcount36_it2u_core_179;
  wire popcount36_it2u_core_180;
  wire popcount36_it2u_core_181;
  wire popcount36_it2u_core_182;
  wire popcount36_it2u_core_185_not;
  wire popcount36_it2u_core_186;
  wire popcount36_it2u_core_187;
  wire popcount36_it2u_core_188;
  wire popcount36_it2u_core_189;
  wire popcount36_it2u_core_190;
  wire popcount36_it2u_core_192;
  wire popcount36_it2u_core_193;
  wire popcount36_it2u_core_194_not;
  wire popcount36_it2u_core_195;
  wire popcount36_it2u_core_197;
  wire popcount36_it2u_core_199;
  wire popcount36_it2u_core_200;
  wire popcount36_it2u_core_201;
  wire popcount36_it2u_core_205;
  wire popcount36_it2u_core_206;
  wire popcount36_it2u_core_210;
  wire popcount36_it2u_core_215;
  wire popcount36_it2u_core_216;
  wire popcount36_it2u_core_217;
  wire popcount36_it2u_core_218;
  wire popcount36_it2u_core_220;
  wire popcount36_it2u_core_221;
  wire popcount36_it2u_core_222;
  wire popcount36_it2u_core_224;
  wire popcount36_it2u_core_227;
  wire popcount36_it2u_core_228;
  wire popcount36_it2u_core_229;
  wire popcount36_it2u_core_230;
  wire popcount36_it2u_core_231;
  wire popcount36_it2u_core_233;
  wire popcount36_it2u_core_234;
  wire popcount36_it2u_core_235;
  wire popcount36_it2u_core_237;
  wire popcount36_it2u_core_240;
  wire popcount36_it2u_core_241;
  wire popcount36_it2u_core_242;
  wire popcount36_it2u_core_243;
  wire popcount36_it2u_core_244;
  wire popcount36_it2u_core_246;
  wire popcount36_it2u_core_248;
  wire popcount36_it2u_core_249;
  wire popcount36_it2u_core_250;
  wire popcount36_it2u_core_252;
  wire popcount36_it2u_core_253;
  wire popcount36_it2u_core_254;
  wire popcount36_it2u_core_255;
  wire popcount36_it2u_core_256;
  wire popcount36_it2u_core_257;
  wire popcount36_it2u_core_259;
  wire popcount36_it2u_core_260;
  wire popcount36_it2u_core_262;
  wire popcount36_it2u_core_263;
  wire popcount36_it2u_core_265;
  wire popcount36_it2u_core_266;
  wire popcount36_it2u_core_267;
  wire popcount36_it2u_core_268;
  wire popcount36_it2u_core_269;
  wire popcount36_it2u_core_270;
  wire popcount36_it2u_core_271;
  wire popcount36_it2u_core_272;
  wire popcount36_it2u_core_273;
  wire popcount36_it2u_core_275;
  wire popcount36_it2u_core_276_not;

  assign popcount36_it2u_core_038 = input_a[26] ^ input_a[1];
  assign popcount36_it2u_core_039 = input_a[0] & input_a[1];
  assign popcount36_it2u_core_040 = ~(input_a[31] & input_a[1]);
  assign popcount36_it2u_core_042 = ~(input_a[12] | input_a[15]);
  assign popcount36_it2u_core_043 = input_a[22] | input_a[33];
  assign popcount36_it2u_core_044 = input_a[17] & input_a[15];
  assign popcount36_it2u_core_045 = ~(input_a[6] | input_a[12]);
  assign popcount36_it2u_core_046 = ~(input_a[32] | input_a[24]);
  assign popcount36_it2u_core_047 = input_a[10] & input_a[24];
  assign popcount36_it2u_core_049 = ~(input_a[4] & input_a[5]);
  assign popcount36_it2u_core_050 = input_a[4] & input_a[5];
  assign popcount36_it2u_core_051 = ~(input_a[7] & input_a[8]);
  assign popcount36_it2u_core_052 = input_a[7] & input_a[8];
  assign popcount36_it2u_core_053 = input_a[6] ^ popcount36_it2u_core_051;
  assign popcount36_it2u_core_054 = input_a[33] ^ input_a[7];
  assign popcount36_it2u_core_055 = popcount36_it2u_core_052 | input_a[6];
  assign popcount36_it2u_core_056 = popcount36_it2u_core_052 & input_a[6];
  assign popcount36_it2u_core_057 = popcount36_it2u_core_049 ^ popcount36_it2u_core_053;
  assign popcount36_it2u_core_059 = input_a[25] | input_a[4];
  assign popcount36_it2u_core_060 = popcount36_it2u_core_050 & popcount36_it2u_core_055;
  assign popcount36_it2u_core_062 = input_a[15] ^ input_a[33];
  assign popcount36_it2u_core_064 = popcount36_it2u_core_056 | popcount36_it2u_core_060;
  assign popcount36_it2u_core_066 = ~(input_a[19] & popcount36_it2u_core_057);
  assign popcount36_it2u_core_067 = input_a[19] & popcount36_it2u_core_057;
  assign popcount36_it2u_core_069 = input_a[7] | input_a[15];
  assign popcount36_it2u_core_079 = ~(input_a[12] ^ input_a[10]);
  assign popcount36_it2u_core_080 = input_a[9] ^ input_a[10];
  assign popcount36_it2u_core_081 = input_a[9] & input_a[10];
  assign popcount36_it2u_core_082 = input_a[11] ^ input_a[12];
  assign popcount36_it2u_core_083 = input_a[11] & input_a[12];
  assign popcount36_it2u_core_084 = popcount36_it2u_core_080 ^ popcount36_it2u_core_082;
  assign popcount36_it2u_core_085 = popcount36_it2u_core_080 & popcount36_it2u_core_082;
  assign popcount36_it2u_core_086 = popcount36_it2u_core_081 ^ popcount36_it2u_core_083;
  assign popcount36_it2u_core_087 = popcount36_it2u_core_081 & popcount36_it2u_core_083;
  assign popcount36_it2u_core_088 = popcount36_it2u_core_086 | popcount36_it2u_core_085;
  assign popcount36_it2u_core_091 = input_a[13] ^ input_a[14];
  assign popcount36_it2u_core_092 = input_a[13] & input_a[14];
  assign popcount36_it2u_core_093 = input_a[16] ^ input_a[17];
  assign popcount36_it2u_core_094 = input_a[16] & input_a[17];
  assign popcount36_it2u_core_095 = input_a[15] ^ popcount36_it2u_core_093;
  assign popcount36_it2u_core_096 = input_a[15] & popcount36_it2u_core_093;
  assign popcount36_it2u_core_097 = popcount36_it2u_core_094 | popcount36_it2u_core_096;
  assign popcount36_it2u_core_099 = ~input_a[11];
  assign popcount36_it2u_core_100 = popcount36_it2u_core_091 & popcount36_it2u_core_095;
  assign popcount36_it2u_core_101 = popcount36_it2u_core_092 ^ popcount36_it2u_core_097;
  assign popcount36_it2u_core_102 = popcount36_it2u_core_092 & popcount36_it2u_core_097;
  assign popcount36_it2u_core_103 = popcount36_it2u_core_101 ^ popcount36_it2u_core_100;
  assign popcount36_it2u_core_104 = popcount36_it2u_core_101 & popcount36_it2u_core_100;
  assign popcount36_it2u_core_105 = popcount36_it2u_core_102 | popcount36_it2u_core_104;
  assign popcount36_it2u_core_109 = popcount36_it2u_core_084 & input_a[21];
  assign popcount36_it2u_core_110 = popcount36_it2u_core_088 ^ popcount36_it2u_core_103;
  assign popcount36_it2u_core_111 = popcount36_it2u_core_088 & popcount36_it2u_core_103;
  assign popcount36_it2u_core_112 = popcount36_it2u_core_110 ^ popcount36_it2u_core_109;
  assign popcount36_it2u_core_113 = popcount36_it2u_core_110 & popcount36_it2u_core_109;
  assign popcount36_it2u_core_114 = popcount36_it2u_core_111 | popcount36_it2u_core_113;
  assign popcount36_it2u_core_115 = popcount36_it2u_core_087 ^ popcount36_it2u_core_105;
  assign popcount36_it2u_core_116 = popcount36_it2u_core_087 & popcount36_it2u_core_105;
  assign popcount36_it2u_core_117 = popcount36_it2u_core_115 ^ popcount36_it2u_core_114;
  assign popcount36_it2u_core_118 = popcount36_it2u_core_115 & popcount36_it2u_core_114;
  assign popcount36_it2u_core_119 = popcount36_it2u_core_116 | popcount36_it2u_core_118;
  assign popcount36_it2u_core_122 = input_a[28] | input_a[16];
  assign popcount36_it2u_core_123 = popcount36_it2u_core_066 & input_a[18];
  assign popcount36_it2u_core_124 = popcount36_it2u_core_067 | popcount36_it2u_core_112;
  assign popcount36_it2u_core_125 = popcount36_it2u_core_067 & popcount36_it2u_core_112;
  assign popcount36_it2u_core_126 = popcount36_it2u_core_124 ^ popcount36_it2u_core_123;
  assign popcount36_it2u_core_127 = popcount36_it2u_core_124 & popcount36_it2u_core_123;
  assign popcount36_it2u_core_128 = popcount36_it2u_core_125 | popcount36_it2u_core_127;
  assign popcount36_it2u_core_131 = popcount36_it2u_core_117 ^ popcount36_it2u_core_128;
  assign popcount36_it2u_core_132 = popcount36_it2u_core_117 & popcount36_it2u_core_128;
  assign popcount36_it2u_core_134 = popcount36_it2u_core_064 ^ popcount36_it2u_core_119;
  assign popcount36_it2u_core_135 = popcount36_it2u_core_064 & popcount36_it2u_core_119;
  assign popcount36_it2u_core_136 = popcount36_it2u_core_134 ^ popcount36_it2u_core_132;
  assign popcount36_it2u_core_137 = popcount36_it2u_core_134 & popcount36_it2u_core_132;
  assign popcount36_it2u_core_138 = popcount36_it2u_core_135 | popcount36_it2u_core_137;
  assign popcount36_it2u_core_140 = ~input_a[23];
  assign popcount36_it2u_core_142 = ~(input_a[32] ^ input_a[18]);
  assign popcount36_it2u_core_145 = input_a[28] ^ input_a[31];
  assign popcount36_it2u_core_147 = input_a[35] & input_a[22];
  assign popcount36_it2u_core_149 = ~(input_a[33] | input_a[13]);
  assign popcount36_it2u_core_150 = input_a[25] ^ popcount36_it2u_core_147;
  assign popcount36_it2u_core_151 = input_a[25] & popcount36_it2u_core_147;
  assign popcount36_it2u_core_155 = input_a[8] | input_a[12];
  assign popcount36_it2u_core_156 = input_a[31] & input_a[20];
  assign popcount36_it2u_core_157 = ~(input_a[19] | input_a[16]);
  assign popcount36_it2u_core_159 = ~(input_a[2] & input_a[16]);
  assign popcount36_it2u_core_160 = input_a[30] & input_a[34];
  assign popcount36_it2u_core_165 = popcount36_it2u_core_156 | popcount36_it2u_core_160;
  assign popcount36_it2u_core_166 = popcount36_it2u_core_156 & popcount36_it2u_core_160;
  assign popcount36_it2u_core_168 = input_a[29] & input_a[18];
  assign popcount36_it2u_core_174 = input_a[27] ^ input_a[27];
  assign popcount36_it2u_core_175 = popcount36_it2u_core_150 & popcount36_it2u_core_165;
  assign popcount36_it2u_core_179 = popcount36_it2u_core_151 ^ popcount36_it2u_core_166;
  assign popcount36_it2u_core_180 = popcount36_it2u_core_151 & popcount36_it2u_core_166;
  assign popcount36_it2u_core_181 = popcount36_it2u_core_179 | popcount36_it2u_core_175;
  assign popcount36_it2u_core_182 = input_a[7] & input_a[21];
  assign popcount36_it2u_core_185_not = ~input_a[22];
  assign popcount36_it2u_core_186 = input_a[23] | input_a[22];
  assign popcount36_it2u_core_187 = input_a[3] & input_a[33];
  assign popcount36_it2u_core_188 = ~(input_a[28] | input_a[27]);
  assign popcount36_it2u_core_189 = input_a[2] & input_a[23];
  assign popcount36_it2u_core_190 = ~(input_a[32] | input_a[11]);
  assign popcount36_it2u_core_192 = input_a[13] ^ input_a[9];
  assign popcount36_it2u_core_193 = popcount36_it2u_core_187 & popcount36_it2u_core_189;
  assign popcount36_it2u_core_194_not = ~input_a[16];
  assign popcount36_it2u_core_195 = input_a[35] ^ input_a[21];
  assign popcount36_it2u_core_197 = input_a[12] & input_a[12];
  assign popcount36_it2u_core_199 = input_a[31] | input_a[17];
  assign popcount36_it2u_core_200 = input_a[32] & input_a[24];
  assign popcount36_it2u_core_201 = ~input_a[30];
  assign popcount36_it2u_core_205 = ~(input_a[7] | input_a[28]);
  assign popcount36_it2u_core_206 = input_a[29] & input_a[27];
  assign popcount36_it2u_core_210 = popcount36_it2u_core_200 & popcount36_it2u_core_206;
  assign popcount36_it2u_core_215 = ~(input_a[8] ^ input_a[3]);
  assign popcount36_it2u_core_216 = ~(input_a[19] ^ input_a[6]);
  assign popcount36_it2u_core_217 = input_a[21] & input_a[22];
  assign popcount36_it2u_core_218 = ~(input_a[15] & input_a[15]);
  assign popcount36_it2u_core_220 = input_a[2] ^ input_a[9];
  assign popcount36_it2u_core_221 = popcount36_it2u_core_193 ^ popcount36_it2u_core_210;
  assign popcount36_it2u_core_222 = popcount36_it2u_core_193 & popcount36_it2u_core_210;
  assign popcount36_it2u_core_224 = ~(input_a[14] ^ input_a[31]);
  assign popcount36_it2u_core_227 = ~(input_a[1] & input_a[30]);
  assign popcount36_it2u_core_228 = ~(input_a[6] | input_a[0]);
  assign popcount36_it2u_core_229 = input_a[13] | input_a[9];
  assign popcount36_it2u_core_230 = ~(input_a[1] & input_a[0]);
  assign popcount36_it2u_core_231 = ~(input_a[28] & input_a[19]);
  assign popcount36_it2u_core_233 = ~input_a[14];
  assign popcount36_it2u_core_234 = ~(input_a[24] ^ input_a[16]);
  assign popcount36_it2u_core_235 = popcount36_it2u_core_181 | popcount36_it2u_core_221;
  assign popcount36_it2u_core_237 = ~popcount36_it2u_core_235;
  assign popcount36_it2u_core_240 = popcount36_it2u_core_180 ^ popcount36_it2u_core_222;
  assign popcount36_it2u_core_241 = popcount36_it2u_core_180 & popcount36_it2u_core_222;
  assign popcount36_it2u_core_242 = popcount36_it2u_core_240 ^ popcount36_it2u_core_235;
  assign popcount36_it2u_core_243 = popcount36_it2u_core_240 & popcount36_it2u_core_235;
  assign popcount36_it2u_core_244 = popcount36_it2u_core_241 | popcount36_it2u_core_243;
  assign popcount36_it2u_core_246 = input_a[23] | input_a[10];
  assign popcount36_it2u_core_248 = ~input_a[3];
  assign popcount36_it2u_core_249 = ~input_a[12];
  assign popcount36_it2u_core_250 = ~input_a[2];
  assign popcount36_it2u_core_252 = popcount36_it2u_core_126 ^ popcount36_it2u_core_230;
  assign popcount36_it2u_core_253 = popcount36_it2u_core_126 & popcount36_it2u_core_230;
  assign popcount36_it2u_core_254 = popcount36_it2u_core_252 ^ input_a[28];
  assign popcount36_it2u_core_255 = popcount36_it2u_core_252 & input_a[28];
  assign popcount36_it2u_core_256 = popcount36_it2u_core_253 | popcount36_it2u_core_255;
  assign popcount36_it2u_core_257 = popcount36_it2u_core_131 | popcount36_it2u_core_237;
  assign popcount36_it2u_core_259 = ~(input_a[30] ^ input_a[31]);
  assign popcount36_it2u_core_260 = popcount36_it2u_core_257 & popcount36_it2u_core_256;
  assign popcount36_it2u_core_262 = popcount36_it2u_core_136 | popcount36_it2u_core_242;
  assign popcount36_it2u_core_263 = popcount36_it2u_core_136 & popcount36_it2u_core_242;
  assign popcount36_it2u_core_265 = popcount36_it2u_core_262 & popcount36_it2u_core_260;
  assign popcount36_it2u_core_266 = popcount36_it2u_core_263 | popcount36_it2u_core_265;
  assign popcount36_it2u_core_267 = popcount36_it2u_core_138 ^ popcount36_it2u_core_244;
  assign popcount36_it2u_core_268 = popcount36_it2u_core_138 & popcount36_it2u_core_244;
  assign popcount36_it2u_core_269 = popcount36_it2u_core_267 ^ popcount36_it2u_core_266;
  assign popcount36_it2u_core_270 = popcount36_it2u_core_267 & popcount36_it2u_core_266;
  assign popcount36_it2u_core_271 = popcount36_it2u_core_268 | popcount36_it2u_core_270;
  assign popcount36_it2u_core_272 = ~(input_a[24] | input_a[17]);
  assign popcount36_it2u_core_273 = ~(input_a[28] ^ input_a[22]);
  assign popcount36_it2u_core_275 = input_a[26] ^ input_a[6];
  assign popcount36_it2u_core_276_not = ~input_a[11];

  assign popcount36_it2u_out[0] = input_a[26];
  assign popcount36_it2u_out[1] = popcount36_it2u_core_254;
  assign popcount36_it2u_out[2] = popcount36_it2u_core_230;
  assign popcount36_it2u_out[3] = popcount36_it2u_core_039;
  assign popcount36_it2u_out[4] = popcount36_it2u_core_269;
  assign popcount36_it2u_out[5] = popcount36_it2u_core_271;
endmodule