// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.44305
// WCE=8.0
// EP=0.786725%
// Printed PDK parameters:
//  Area=35529853.0
//  Delay=56517156.0
//  Power=1570100.0

module popcount29_khno(input [28:0] input_a, output [4:0] popcount29_khno_out);
  wire popcount29_khno_core_032;
  wire popcount29_khno_core_034;
  wire popcount29_khno_core_035;
  wire popcount29_khno_core_037;
  wire popcount29_khno_core_038;
  wire popcount29_khno_core_039;
  wire popcount29_khno_core_040;
  wire popcount29_khno_core_041;
  wire popcount29_khno_core_043;
  wire popcount29_khno_core_045;
  wire popcount29_khno_core_046;
  wire popcount29_khno_core_048;
  wire popcount29_khno_core_050;
  wire popcount29_khno_core_052;
  wire popcount29_khno_core_053;
  wire popcount29_khno_core_054;
  wire popcount29_khno_core_056;
  wire popcount29_khno_core_057;
  wire popcount29_khno_core_058;
  wire popcount29_khno_core_059;
  wire popcount29_khno_core_061;
  wire popcount29_khno_core_062;
  wire popcount29_khno_core_064;
  wire popcount29_khno_core_065;
  wire popcount29_khno_core_066;
  wire popcount29_khno_core_067;
  wire popcount29_khno_core_068;
  wire popcount29_khno_core_070;
  wire popcount29_khno_core_071;
  wire popcount29_khno_core_074;
  wire popcount29_khno_core_075;
  wire popcount29_khno_core_077;
  wire popcount29_khno_core_078;
  wire popcount29_khno_core_079;
  wire popcount29_khno_core_080;
  wire popcount29_khno_core_082;
  wire popcount29_khno_core_087;
  wire popcount29_khno_core_090;
  wire popcount29_khno_core_091;
  wire popcount29_khno_core_092;
  wire popcount29_khno_core_093;
  wire popcount29_khno_core_094;
  wire popcount29_khno_core_095;
  wire popcount29_khno_core_096;
  wire popcount29_khno_core_097;
  wire popcount29_khno_core_098;
  wire popcount29_khno_core_099;
  wire popcount29_khno_core_100;
  wire popcount29_khno_core_102;
  wire popcount29_khno_core_104;
  wire popcount29_khno_core_105;
  wire popcount29_khno_core_106;
  wire popcount29_khno_core_107;
  wire popcount29_khno_core_108;
  wire popcount29_khno_core_109;
  wire popcount29_khno_core_110;
  wire popcount29_khno_core_113;
  wire popcount29_khno_core_114;
  wire popcount29_khno_core_115;
  wire popcount29_khno_core_116;
  wire popcount29_khno_core_118;
  wire popcount29_khno_core_119;
  wire popcount29_khno_core_121;
  wire popcount29_khno_core_123;
  wire popcount29_khno_core_124;
  wire popcount29_khno_core_125;
  wire popcount29_khno_core_126;
  wire popcount29_khno_core_128;
  wire popcount29_khno_core_131;
  wire popcount29_khno_core_132;
  wire popcount29_khno_core_133;
  wire popcount29_khno_core_134;
  wire popcount29_khno_core_135;
  wire popcount29_khno_core_138;
  wire popcount29_khno_core_142;
  wire popcount29_khno_core_143;
  wire popcount29_khno_core_144;
  wire popcount29_khno_core_145;
  wire popcount29_khno_core_146;
  wire popcount29_khno_core_148;
  wire popcount29_khno_core_150;
  wire popcount29_khno_core_151;
  wire popcount29_khno_core_152;
  wire popcount29_khno_core_154;
  wire popcount29_khno_core_155;
  wire popcount29_khno_core_156;
  wire popcount29_khno_core_159;
  wire popcount29_khno_core_160;
  wire popcount29_khno_core_161;
  wire popcount29_khno_core_162;
  wire popcount29_khno_core_163;
  wire popcount29_khno_core_164;
  wire popcount29_khno_core_168;
  wire popcount29_khno_core_170_not;
  wire popcount29_khno_core_171;
  wire popcount29_khno_core_173;
  wire popcount29_khno_core_175;
  wire popcount29_khno_core_176;
  wire popcount29_khno_core_178;
  wire popcount29_khno_core_179;
  wire popcount29_khno_core_180;
  wire popcount29_khno_core_184;
  wire popcount29_khno_core_185;
  wire popcount29_khno_core_187;
  wire popcount29_khno_core_188;
  wire popcount29_khno_core_189;
  wire popcount29_khno_core_190;
  wire popcount29_khno_core_191;
  wire popcount29_khno_core_192;
  wire popcount29_khno_core_193;
  wire popcount29_khno_core_194;
  wire popcount29_khno_core_195;
  wire popcount29_khno_core_196;
  wire popcount29_khno_core_197;
  wire popcount29_khno_core_198;
  wire popcount29_khno_core_199;
  wire popcount29_khno_core_200;
  wire popcount29_khno_core_201;
  wire popcount29_khno_core_202;
  wire popcount29_khno_core_204;
  wire popcount29_khno_core_205;
  wire popcount29_khno_core_206;

  assign popcount29_khno_core_032 = input_a[23] & input_a[2];
  assign popcount29_khno_core_034 = input_a[0] & input_a[1];
  assign popcount29_khno_core_035 = popcount29_khno_core_032 | popcount29_khno_core_034;
  assign popcount29_khno_core_037 = input_a[3] ^ input_a[4];
  assign popcount29_khno_core_038 = input_a[3] & input_a[4];
  assign popcount29_khno_core_039 = ~(input_a[5] & input_a[6]);
  assign popcount29_khno_core_040 = input_a[5] & input_a[6];
  assign popcount29_khno_core_041 = popcount29_khno_core_037 ^ popcount29_khno_core_039;
  assign popcount29_khno_core_043 = input_a[3] ^ popcount29_khno_core_040;
  assign popcount29_khno_core_045 = popcount29_khno_core_043 | popcount29_khno_core_037;
  assign popcount29_khno_core_046 = ~input_a[22];
  assign popcount29_khno_core_048 = input_a[26] | input_a[1];
  assign popcount29_khno_core_050 = popcount29_khno_core_035 ^ popcount29_khno_core_045;
  assign popcount29_khno_core_052 = popcount29_khno_core_050 ^ popcount29_khno_core_041;
  assign popcount29_khno_core_053 = popcount29_khno_core_050 & popcount29_khno_core_041;
  assign popcount29_khno_core_054 = popcount29_khno_core_035 | popcount29_khno_core_053;
  assign popcount29_khno_core_056 = input_a[3] | input_a[26];
  assign popcount29_khno_core_057 = popcount29_khno_core_038 | popcount29_khno_core_054;
  assign popcount29_khno_core_058 = ~(input_a[18] & input_a[15]);
  assign popcount29_khno_core_059 = input_a[16] ^ input_a[13];
  assign popcount29_khno_core_061 = input_a[17] | input_a[18];
  assign popcount29_khno_core_062 = ~input_a[28];
  assign popcount29_khno_core_064 = input_a[8] | input_a[22];
  assign popcount29_khno_core_065 = ~(input_a[23] & input_a[4]);
  assign popcount29_khno_core_066 = input_a[16] | input_a[21];
  assign popcount29_khno_core_067 = input_a[10] & input_a[11];
  assign popcount29_khno_core_068 = input_a[10] | input_a[11];
  assign popcount29_khno_core_070 = input_a[20] | input_a[27];
  assign popcount29_khno_core_071 = input_a[25] & popcount29_khno_core_068;
  assign popcount29_khno_core_074 = popcount29_khno_core_067 | popcount29_khno_core_071;
  assign popcount29_khno_core_075 = ~(input_a[2] | input_a[13]);
  assign popcount29_khno_core_077 = input_a[16] ^ input_a[27];
  assign popcount29_khno_core_078 = ~(input_a[13] ^ input_a[4]);
  assign popcount29_khno_core_079 = popcount29_khno_core_064 ^ popcount29_khno_core_074;
  assign popcount29_khno_core_080 = popcount29_khno_core_064 & popcount29_khno_core_074;
  assign popcount29_khno_core_082 = ~(input_a[9] & input_a[8]);
  assign popcount29_khno_core_087 = ~(input_a[28] & input_a[25]);
  assign popcount29_khno_core_090 = input_a[26] & input_a[24];
  assign popcount29_khno_core_091 = popcount29_khno_core_052 ^ popcount29_khno_core_079;
  assign popcount29_khno_core_092 = popcount29_khno_core_052 & popcount29_khno_core_079;
  assign popcount29_khno_core_093 = popcount29_khno_core_091 ^ popcount29_khno_core_090;
  assign popcount29_khno_core_094 = popcount29_khno_core_091 & popcount29_khno_core_090;
  assign popcount29_khno_core_095 = popcount29_khno_core_092 | popcount29_khno_core_094;
  assign popcount29_khno_core_096 = popcount29_khno_core_057 ^ popcount29_khno_core_080;
  assign popcount29_khno_core_097 = popcount29_khno_core_057 & popcount29_khno_core_080;
  assign popcount29_khno_core_098 = popcount29_khno_core_096 ^ popcount29_khno_core_095;
  assign popcount29_khno_core_099 = popcount29_khno_core_096 & popcount29_khno_core_095;
  assign popcount29_khno_core_100 = popcount29_khno_core_097 | popcount29_khno_core_099;
  assign popcount29_khno_core_102 = ~(input_a[4] ^ input_a[10]);
  assign popcount29_khno_core_104 = ~(input_a[19] & input_a[20]);
  assign popcount29_khno_core_105 = ~(input_a[23] ^ input_a[14]);
  assign popcount29_khno_core_106 = ~(input_a[20] ^ input_a[13]);
  assign popcount29_khno_core_107 = input_a[12] & input_a[16];
  assign popcount29_khno_core_108 = input_a[3] ^ input_a[1];
  assign popcount29_khno_core_109 = input_a[14] & input_a[15];
  assign popcount29_khno_core_110 = popcount29_khno_core_107 | popcount29_khno_core_109;
  assign popcount29_khno_core_113 = input_a[17] & input_a[9];
  assign popcount29_khno_core_114 = ~input_a[9];
  assign popcount29_khno_core_115 = input_a[20] & input_a[28];
  assign popcount29_khno_core_116 = ~(input_a[4] & input_a[0]);
  assign popcount29_khno_core_118 = popcount29_khno_core_113 ^ popcount29_khno_core_115;
  assign popcount29_khno_core_119 = popcount29_khno_core_113 & popcount29_khno_core_115;
  assign popcount29_khno_core_121 = ~input_a[4];
  assign popcount29_khno_core_123 = ~(input_a[6] & input_a[13]);
  assign popcount29_khno_core_124 = input_a[20] | input_a[20];
  assign popcount29_khno_core_125 = popcount29_khno_core_110 ^ popcount29_khno_core_118;
  assign popcount29_khno_core_126 = popcount29_khno_core_110 & popcount29_khno_core_118;
  assign popcount29_khno_core_128 = ~(input_a[21] & input_a[1]);
  assign popcount29_khno_core_131 = ~(input_a[19] ^ input_a[19]);
  assign popcount29_khno_core_132 = popcount29_khno_core_119 | popcount29_khno_core_126;
  assign popcount29_khno_core_133 = input_a[13] & input_a[28];
  assign popcount29_khno_core_134 = ~input_a[19];
  assign popcount29_khno_core_135 = ~(input_a[2] ^ input_a[21]);
  assign popcount29_khno_core_138 = input_a[2] ^ input_a[7];
  assign popcount29_khno_core_142 = input_a[3] ^ input_a[4];
  assign popcount29_khno_core_143 = ~input_a[21];
  assign popcount29_khno_core_144 = ~(input_a[28] ^ input_a[17]);
  assign popcount29_khno_core_145 = ~(input_a[16] ^ input_a[13]);
  assign popcount29_khno_core_146 = input_a[15] ^ input_a[10];
  assign popcount29_khno_core_148 = ~(input_a[2] | input_a[27]);
  assign popcount29_khno_core_150 = input_a[22] & input_a[11];
  assign popcount29_khno_core_151 = input_a[15] ^ input_a[17];
  assign popcount29_khno_core_152 = input_a[18] & input_a[12];
  assign popcount29_khno_core_154 = ~(input_a[7] & input_a[27]);
  assign popcount29_khno_core_155 = input_a[7] & input_a[27];
  assign popcount29_khno_core_156 = input_a[19] | popcount29_khno_core_155;
  assign popcount29_khno_core_159 = input_a[19] | popcount29_khno_core_154;
  assign popcount29_khno_core_160 = ~(input_a[18] & input_a[3]);
  assign popcount29_khno_core_161 = popcount29_khno_core_159 ^ input_a[19];
  assign popcount29_khno_core_162 = ~(input_a[5] ^ input_a[5]);
  assign popcount29_khno_core_163 = input_a[19] ^ input_a[9];
  assign popcount29_khno_core_164 = input_a[19] | popcount29_khno_core_156;
  assign popcount29_khno_core_168 = input_a[28] ^ input_a[11];
  assign popcount29_khno_core_170_not = ~input_a[12];
  assign popcount29_khno_core_171 = popcount29_khno_core_125 ^ popcount29_khno_core_161;
  assign popcount29_khno_core_173 = ~popcount29_khno_core_171;
  assign popcount29_khno_core_175 = popcount29_khno_core_125 | popcount29_khno_core_171;
  assign popcount29_khno_core_176 = popcount29_khno_core_132 ^ popcount29_khno_core_164;
  assign popcount29_khno_core_178 = popcount29_khno_core_176 ^ popcount29_khno_core_175;
  assign popcount29_khno_core_179 = popcount29_khno_core_176 & popcount29_khno_core_175;
  assign popcount29_khno_core_180 = popcount29_khno_core_132 | popcount29_khno_core_179;
  assign popcount29_khno_core_184 = ~(input_a[27] & input_a[9]);
  assign popcount29_khno_core_185 = ~(input_a[27] ^ input_a[13]);
  assign popcount29_khno_core_187 = input_a[21] & input_a[18];
  assign popcount29_khno_core_188 = popcount29_khno_core_093 ^ popcount29_khno_core_173;
  assign popcount29_khno_core_189 = popcount29_khno_core_093 & popcount29_khno_core_173;
  assign popcount29_khno_core_190 = popcount29_khno_core_188 ^ popcount29_khno_core_187;
  assign popcount29_khno_core_191 = popcount29_khno_core_188 & popcount29_khno_core_187;
  assign popcount29_khno_core_192 = popcount29_khno_core_189 | popcount29_khno_core_191;
  assign popcount29_khno_core_193 = popcount29_khno_core_098 ^ popcount29_khno_core_178;
  assign popcount29_khno_core_194 = popcount29_khno_core_098 & popcount29_khno_core_178;
  assign popcount29_khno_core_195 = popcount29_khno_core_193 ^ popcount29_khno_core_192;
  assign popcount29_khno_core_196 = popcount29_khno_core_193 & popcount29_khno_core_192;
  assign popcount29_khno_core_197 = popcount29_khno_core_194 | popcount29_khno_core_196;
  assign popcount29_khno_core_198 = popcount29_khno_core_100 ^ popcount29_khno_core_180;
  assign popcount29_khno_core_199 = popcount29_khno_core_100 & popcount29_khno_core_180;
  assign popcount29_khno_core_200 = popcount29_khno_core_198 ^ popcount29_khno_core_197;
  assign popcount29_khno_core_201 = popcount29_khno_core_198 & popcount29_khno_core_197;
  assign popcount29_khno_core_202 = popcount29_khno_core_199 | popcount29_khno_core_201;
  assign popcount29_khno_core_204 = input_a[2] | input_a[0];
  assign popcount29_khno_core_205 = ~(input_a[24] ^ input_a[23]);
  assign popcount29_khno_core_206 = input_a[22] ^ input_a[10];

  assign popcount29_khno_out[0] = input_a[13];
  assign popcount29_khno_out[1] = popcount29_khno_core_190;
  assign popcount29_khno_out[2] = popcount29_khno_core_195;
  assign popcount29_khno_out[3] = popcount29_khno_core_200;
  assign popcount29_khno_out[4] = popcount29_khno_core_202;
endmodule