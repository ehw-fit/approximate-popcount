// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.68307
// WCE=47.0
// EP=0.931451%
// Printed PDK parameters:
//  Area=144537987.0
//  Delay=110269552.0
//  Power=7426200.0

module popcount47_8o2d(input [46:0] input_a, output [5:0] popcount47_8o2d_out);
  wire popcount47_8o2d_core_049;
  wire popcount47_8o2d_core_050;
  wire popcount47_8o2d_core_051;
  wire popcount47_8o2d_core_052;
  wire popcount47_8o2d_core_059;
  wire popcount47_8o2d_core_060;
  wire popcount47_8o2d_core_066;
  wire popcount47_8o2d_core_067;
  wire popcount47_8o2d_core_068;
  wire popcount47_8o2d_core_069;
  wire popcount47_8o2d_core_070;
  wire popcount47_8o2d_core_071;
  wire popcount47_8o2d_core_072;
  wire popcount47_8o2d_core_073;
  wire popcount47_8o2d_core_074;
  wire popcount47_8o2d_core_075;
  wire popcount47_8o2d_core_076;
  wire popcount47_8o2d_core_077;
  wire popcount47_8o2d_core_078;
  wire popcount47_8o2d_core_079;
  wire popcount47_8o2d_core_080;
  wire popcount47_8o2d_core_081;
  wire popcount47_8o2d_core_082;
  wire popcount47_8o2d_core_083;
  wire popcount47_8o2d_core_084;
  wire popcount47_8o2d_core_085;
  wire popcount47_8o2d_core_086;
  wire popcount47_8o2d_core_087;
  wire popcount47_8o2d_core_088;
  wire popcount47_8o2d_core_089;
  wire popcount47_8o2d_core_090_not;
  wire popcount47_8o2d_core_091_not;
  wire popcount47_8o2d_core_092;
  wire popcount47_8o2d_core_093;
  wire popcount47_8o2d_core_094;
  wire popcount47_8o2d_core_095;
  wire popcount47_8o2d_core_096;
  wire popcount47_8o2d_core_097;
  wire popcount47_8o2d_core_098;
  wire popcount47_8o2d_core_099;
  wire popcount47_8o2d_core_100;
  wire popcount47_8o2d_core_101;
  wire popcount47_8o2d_core_104;
  wire popcount47_8o2d_core_105;
  wire popcount47_8o2d_core_107;
  wire popcount47_8o2d_core_108;
  wire popcount47_8o2d_core_109;
  wire popcount47_8o2d_core_110;
  wire popcount47_8o2d_core_111;
  wire popcount47_8o2d_core_112;
  wire popcount47_8o2d_core_113;
  wire popcount47_8o2d_core_114;
  wire popcount47_8o2d_core_115;
  wire popcount47_8o2d_core_116;
  wire popcount47_8o2d_core_117;
  wire popcount47_8o2d_core_118;
  wire popcount47_8o2d_core_120;
  wire popcount47_8o2d_core_121;
  wire popcount47_8o2d_core_122;
  wire popcount47_8o2d_core_123;
  wire popcount47_8o2d_core_124;
  wire popcount47_8o2d_core_125;
  wire popcount47_8o2d_core_126;
  wire popcount47_8o2d_core_127;
  wire popcount47_8o2d_core_128;
  wire popcount47_8o2d_core_129;
  wire popcount47_8o2d_core_130;
  wire popcount47_8o2d_core_131;
  wire popcount47_8o2d_core_132;
  wire popcount47_8o2d_core_133;
  wire popcount47_8o2d_core_134;
  wire popcount47_8o2d_core_135;
  wire popcount47_8o2d_core_136;
  wire popcount47_8o2d_core_137;
  wire popcount47_8o2d_core_138;
  wire popcount47_8o2d_core_139;
  wire popcount47_8o2d_core_140;
  wire popcount47_8o2d_core_141;
  wire popcount47_8o2d_core_142;
  wire popcount47_8o2d_core_143;
  wire popcount47_8o2d_core_144;
  wire popcount47_8o2d_core_145;
  wire popcount47_8o2d_core_146;
  wire popcount47_8o2d_core_147;
  wire popcount47_8o2d_core_148;
  wire popcount47_8o2d_core_149;
  wire popcount47_8o2d_core_150;
  wire popcount47_8o2d_core_151;
  wire popcount47_8o2d_core_152;
  wire popcount47_8o2d_core_153;
  wire popcount47_8o2d_core_154;
  wire popcount47_8o2d_core_157;
  wire popcount47_8o2d_core_158;
  wire popcount47_8o2d_core_162;
  wire popcount47_8o2d_core_163;
  wire popcount47_8o2d_core_164;
  wire popcount47_8o2d_core_165;
  wire popcount47_8o2d_core_166;
  wire popcount47_8o2d_core_167;
  wire popcount47_8o2d_core_168;
  wire popcount47_8o2d_core_169;
  wire popcount47_8o2d_core_170;
  wire popcount47_8o2d_core_171;
  wire popcount47_8o2d_core_172_not;
  wire popcount47_8o2d_core_174;
  wire popcount47_8o2d_core_175;
  wire popcount47_8o2d_core_176;
  wire popcount47_8o2d_core_177;
  wire popcount47_8o2d_core_178;
  wire popcount47_8o2d_core_179;
  wire popcount47_8o2d_core_180;
  wire popcount47_8o2d_core_181;
  wire popcount47_8o2d_core_182;
  wire popcount47_8o2d_core_183;
  wire popcount47_8o2d_core_184;
  wire popcount47_8o2d_core_185;
  wire popcount47_8o2d_core_186;
  wire popcount47_8o2d_core_187;
  wire popcount47_8o2d_core_188;
  wire popcount47_8o2d_core_189;
  wire popcount47_8o2d_core_190;
  wire popcount47_8o2d_core_191;
  wire popcount47_8o2d_core_192;
  wire popcount47_8o2d_core_193;
  wire popcount47_8o2d_core_194;
  wire popcount47_8o2d_core_195;
  wire popcount47_8o2d_core_196;
  wire popcount47_8o2d_core_197;
  wire popcount47_8o2d_core_198;
  wire popcount47_8o2d_core_199;
  wire popcount47_8o2d_core_200;
  wire popcount47_8o2d_core_201;
  wire popcount47_8o2d_core_202;
  wire popcount47_8o2d_core_203;
  wire popcount47_8o2d_core_204;
  wire popcount47_8o2d_core_205;
  wire popcount47_8o2d_core_206;
  wire popcount47_8o2d_core_207;
  wire popcount47_8o2d_core_208;
  wire popcount47_8o2d_core_209;
  wire popcount47_8o2d_core_210;
  wire popcount47_8o2d_core_211;
  wire popcount47_8o2d_core_212;
  wire popcount47_8o2d_core_213;
  wire popcount47_8o2d_core_214;
  wire popcount47_8o2d_core_215;
  wire popcount47_8o2d_core_216;
  wire popcount47_8o2d_core_217;
  wire popcount47_8o2d_core_218;
  wire popcount47_8o2d_core_219;
  wire popcount47_8o2d_core_220;
  wire popcount47_8o2d_core_221;
  wire popcount47_8o2d_core_222;
  wire popcount47_8o2d_core_223;
  wire popcount47_8o2d_core_224;
  wire popcount47_8o2d_core_225;
  wire popcount47_8o2d_core_226;
  wire popcount47_8o2d_core_227;
  wire popcount47_8o2d_core_228;
  wire popcount47_8o2d_core_229;
  wire popcount47_8o2d_core_230;
  wire popcount47_8o2d_core_231;
  wire popcount47_8o2d_core_232;
  wire popcount47_8o2d_core_233;
  wire popcount47_8o2d_core_234;
  wire popcount47_8o2d_core_235;
  wire popcount47_8o2d_core_236;
  wire popcount47_8o2d_core_237;
  wire popcount47_8o2d_core_239;
  wire popcount47_8o2d_core_240;
  wire popcount47_8o2d_core_242;
  wire popcount47_8o2d_core_243;
  wire popcount47_8o2d_core_244;
  wire popcount47_8o2d_core_245;
  wire popcount47_8o2d_core_249;
  wire popcount47_8o2d_core_250;
  wire popcount47_8o2d_core_256;
  wire popcount47_8o2d_core_257;
  wire popcount47_8o2d_core_259;
  wire popcount47_8o2d_core_260;
  wire popcount47_8o2d_core_261;
  wire popcount47_8o2d_core_266;
  wire popcount47_8o2d_core_267;
  wire popcount47_8o2d_core_268;
  wire popcount47_8o2d_core_269;
  wire popcount47_8o2d_core_270;
  wire popcount47_8o2d_core_271;
  wire popcount47_8o2d_core_272;
  wire popcount47_8o2d_core_273;
  wire popcount47_8o2d_core_274;
  wire popcount47_8o2d_core_276;
  wire popcount47_8o2d_core_277;
  wire popcount47_8o2d_core_280;
  wire popcount47_8o2d_core_281;
  wire popcount47_8o2d_core_283;
  wire popcount47_8o2d_core_284;
  wire popcount47_8o2d_core_285;
  wire popcount47_8o2d_core_287;
  wire popcount47_8o2d_core_288;
  wire popcount47_8o2d_core_289;
  wire popcount47_8o2d_core_290;
  wire popcount47_8o2d_core_291;
  wire popcount47_8o2d_core_292;
  wire popcount47_8o2d_core_293;
  wire popcount47_8o2d_core_294;
  wire popcount47_8o2d_core_295;
  wire popcount47_8o2d_core_296;
  wire popcount47_8o2d_core_297;
  wire popcount47_8o2d_core_298;
  wire popcount47_8o2d_core_299;
  wire popcount47_8o2d_core_302;
  wire popcount47_8o2d_core_303;
  wire popcount47_8o2d_core_304;
  wire popcount47_8o2d_core_305;
  wire popcount47_8o2d_core_306;
  wire popcount47_8o2d_core_307;
  wire popcount47_8o2d_core_308;
  wire popcount47_8o2d_core_311;
  wire popcount47_8o2d_core_312;
  wire popcount47_8o2d_core_314;
  wire popcount47_8o2d_core_315;
  wire popcount47_8o2d_core_316;
  wire popcount47_8o2d_core_317;
  wire popcount47_8o2d_core_318;
  wire popcount47_8o2d_core_319;
  wire popcount47_8o2d_core_320;
  wire popcount47_8o2d_core_321;
  wire popcount47_8o2d_core_322;
  wire popcount47_8o2d_core_323;
  wire popcount47_8o2d_core_324;
  wire popcount47_8o2d_core_325;
  wire popcount47_8o2d_core_328;
  wire popcount47_8o2d_core_329;
  wire popcount47_8o2d_core_331;
  wire popcount47_8o2d_core_332;
  wire popcount47_8o2d_core_333;
  wire popcount47_8o2d_core_334;
  wire popcount47_8o2d_core_335;
  wire popcount47_8o2d_core_336;
  wire popcount47_8o2d_core_337;
  wire popcount47_8o2d_core_338;
  wire popcount47_8o2d_core_339;
  wire popcount47_8o2d_core_340;
  wire popcount47_8o2d_core_341;
  wire popcount47_8o2d_core_342;
  wire popcount47_8o2d_core_343;
  wire popcount47_8o2d_core_344;
  wire popcount47_8o2d_core_345;
  wire popcount47_8o2d_core_346;
  wire popcount47_8o2d_core_347;
  wire popcount47_8o2d_core_348;
  wire popcount47_8o2d_core_349;
  wire popcount47_8o2d_core_350;
  wire popcount47_8o2d_core_353;
  wire popcount47_8o2d_core_354;
  wire popcount47_8o2d_core_355_not;
  wire popcount47_8o2d_core_357;
  wire popcount47_8o2d_core_358;
  wire popcount47_8o2d_core_359;
  wire popcount47_8o2d_core_360;
  wire popcount47_8o2d_core_361;
  wire popcount47_8o2d_core_362;
  wire popcount47_8o2d_core_363;
  wire popcount47_8o2d_core_364;
  wire popcount47_8o2d_core_365;
  wire popcount47_8o2d_core_366;
  wire popcount47_8o2d_core_367;
  wire popcount47_8o2d_core_368;
  wire popcount47_8o2d_core_369;
  wire popcount47_8o2d_core_370;
  wire popcount47_8o2d_core_371;
  wire popcount47_8o2d_core_372;

  assign popcount47_8o2d_core_049 = input_a[0] ^ input_a[1];
  assign popcount47_8o2d_core_050 = input_a[0] & input_a[1];
  assign popcount47_8o2d_core_051 = input_a[3] ^ input_a[4];
  assign popcount47_8o2d_core_052 = input_a[3] & input_a[4];
  assign popcount47_8o2d_core_059 = popcount47_8o2d_core_050 ^ popcount47_8o2d_core_052;
  assign popcount47_8o2d_core_060 = popcount47_8o2d_core_050 & popcount47_8o2d_core_052;
  assign popcount47_8o2d_core_066 = input_a[6] ^ input_a[7];
  assign popcount47_8o2d_core_067 = input_a[6] & input_a[25];
  assign popcount47_8o2d_core_068 = input_a[5] ^ popcount47_8o2d_core_066;
  assign popcount47_8o2d_core_069 = input_a[11] & popcount47_8o2d_core_066;
  assign popcount47_8o2d_core_070 = popcount47_8o2d_core_067 ^ popcount47_8o2d_core_069;
  assign popcount47_8o2d_core_071 = popcount47_8o2d_core_067 & popcount47_8o2d_core_069;
  assign popcount47_8o2d_core_072 = input_a[9] ^ input_a[10];
  assign popcount47_8o2d_core_073 = ~(input_a[3] & input_a[10]);
  assign popcount47_8o2d_core_074 = input_a[8] ^ popcount47_8o2d_core_072;
  assign popcount47_8o2d_core_075 = input_a[8] & popcount47_8o2d_core_072;
  assign popcount47_8o2d_core_076 = popcount47_8o2d_core_073 ^ popcount47_8o2d_core_075;
  assign popcount47_8o2d_core_077 = popcount47_8o2d_core_073 & popcount47_8o2d_core_075;
  assign popcount47_8o2d_core_078 = input_a[17] ^ popcount47_8o2d_core_074;
  assign popcount47_8o2d_core_079 = popcount47_8o2d_core_068 & popcount47_8o2d_core_074;
  assign popcount47_8o2d_core_080 = popcount47_8o2d_core_070 ^ popcount47_8o2d_core_076;
  assign popcount47_8o2d_core_081 = popcount47_8o2d_core_070 & popcount47_8o2d_core_076;
  assign popcount47_8o2d_core_082 = input_a[29] ^ popcount47_8o2d_core_079;
  assign popcount47_8o2d_core_083 = popcount47_8o2d_core_080 & popcount47_8o2d_core_079;
  assign popcount47_8o2d_core_084 = input_a[43] | popcount47_8o2d_core_083;
  assign popcount47_8o2d_core_085 = popcount47_8o2d_core_071 ^ popcount47_8o2d_core_077;
  assign popcount47_8o2d_core_086 = popcount47_8o2d_core_071 & popcount47_8o2d_core_077;
  assign popcount47_8o2d_core_087 = popcount47_8o2d_core_085 ^ popcount47_8o2d_core_084;
  assign popcount47_8o2d_core_088 = popcount47_8o2d_core_085 & popcount47_8o2d_core_084;
  assign popcount47_8o2d_core_089 = popcount47_8o2d_core_086 | popcount47_8o2d_core_088;
  assign popcount47_8o2d_core_090_not = ~popcount47_8o2d_core_078;
  assign popcount47_8o2d_core_091_not = ~popcount47_8o2d_core_078;
  assign popcount47_8o2d_core_092 = popcount47_8o2d_core_059 | popcount47_8o2d_core_082;
  assign popcount47_8o2d_core_093 = popcount47_8o2d_core_059 & input_a[9];
  assign popcount47_8o2d_core_094 = ~(popcount47_8o2d_core_092 & popcount47_8o2d_core_091_not);
  assign popcount47_8o2d_core_095 = popcount47_8o2d_core_092 & popcount47_8o2d_core_091_not;
  assign popcount47_8o2d_core_096 = popcount47_8o2d_core_093 | popcount47_8o2d_core_095;
  assign popcount47_8o2d_core_097 = popcount47_8o2d_core_060 ^ popcount47_8o2d_core_087;
  assign popcount47_8o2d_core_098 = popcount47_8o2d_core_060 & popcount47_8o2d_core_087;
  assign popcount47_8o2d_core_099 = popcount47_8o2d_core_097 ^ popcount47_8o2d_core_096;
  assign popcount47_8o2d_core_100 = popcount47_8o2d_core_097 & popcount47_8o2d_core_096;
  assign popcount47_8o2d_core_101 = popcount47_8o2d_core_098 | popcount47_8o2d_core_100;
  assign popcount47_8o2d_core_104 = popcount47_8o2d_core_089 ^ popcount47_8o2d_core_101;
  assign popcount47_8o2d_core_105 = popcount47_8o2d_core_089 & popcount47_8o2d_core_101;
  assign popcount47_8o2d_core_107 = input_a[0] ^ input_a[13];
  assign popcount47_8o2d_core_108 = input_a[27] & input_a[13];
  assign popcount47_8o2d_core_109 = input_a[11] ^ popcount47_8o2d_core_107;
  assign popcount47_8o2d_core_110 = input_a[11] & popcount47_8o2d_core_107;
  assign popcount47_8o2d_core_111 = popcount47_8o2d_core_108 ^ popcount47_8o2d_core_110;
  assign popcount47_8o2d_core_112 = input_a[30] & popcount47_8o2d_core_110;
  assign popcount47_8o2d_core_113 = input_a[15] ^ input_a[16];
  assign popcount47_8o2d_core_114 = input_a[15] & input_a[16];
  assign popcount47_8o2d_core_115 = input_a[14] ^ popcount47_8o2d_core_113;
  assign popcount47_8o2d_core_116 = input_a[14] & popcount47_8o2d_core_113;
  assign popcount47_8o2d_core_117 = popcount47_8o2d_core_114 ^ popcount47_8o2d_core_116;
  assign popcount47_8o2d_core_118 = popcount47_8o2d_core_114 & popcount47_8o2d_core_116;
  assign popcount47_8o2d_core_120 = popcount47_8o2d_core_109 & popcount47_8o2d_core_115;
  assign popcount47_8o2d_core_121 = popcount47_8o2d_core_111 ^ input_a[26];
  assign popcount47_8o2d_core_122 = popcount47_8o2d_core_111 & input_a[8];
  assign popcount47_8o2d_core_123 = popcount47_8o2d_core_121 ^ popcount47_8o2d_core_120;
  assign popcount47_8o2d_core_124 = popcount47_8o2d_core_121 & popcount47_8o2d_core_120;
  assign popcount47_8o2d_core_125 = popcount47_8o2d_core_122 | popcount47_8o2d_core_124;
  assign popcount47_8o2d_core_126 = popcount47_8o2d_core_112 ^ popcount47_8o2d_core_118;
  assign popcount47_8o2d_core_127 = popcount47_8o2d_core_112 & popcount47_8o2d_core_118;
  assign popcount47_8o2d_core_128 = popcount47_8o2d_core_126 ^ popcount47_8o2d_core_125;
  assign popcount47_8o2d_core_129 = popcount47_8o2d_core_126 & popcount47_8o2d_core_125;
  assign popcount47_8o2d_core_130 = popcount47_8o2d_core_127 | popcount47_8o2d_core_129;
  assign popcount47_8o2d_core_131 = input_a[18] ^ input_a[19];
  assign popcount47_8o2d_core_132 = input_a[18] & input_a[19];
  assign popcount47_8o2d_core_133 = input_a[17] ^ popcount47_8o2d_core_131;
  assign popcount47_8o2d_core_134 = input_a[17] & popcount47_8o2d_core_131;
  assign popcount47_8o2d_core_135 = popcount47_8o2d_core_132 ^ popcount47_8o2d_core_134;
  assign popcount47_8o2d_core_136 = popcount47_8o2d_core_132 & popcount47_8o2d_core_134;
  assign popcount47_8o2d_core_137 = ~(input_a[21] & input_a[44]);
  assign popcount47_8o2d_core_138 = input_a[21] & input_a[6];
  assign popcount47_8o2d_core_139 = input_a[20] ^ popcount47_8o2d_core_137;
  assign popcount47_8o2d_core_140 = input_a[20] & popcount47_8o2d_core_137;
  assign popcount47_8o2d_core_141 = popcount47_8o2d_core_138 | popcount47_8o2d_core_140;
  assign popcount47_8o2d_core_142 = popcount47_8o2d_core_138 & popcount47_8o2d_core_140;
  assign popcount47_8o2d_core_143 = popcount47_8o2d_core_133 ^ popcount47_8o2d_core_139;
  assign popcount47_8o2d_core_144 = ~popcount47_8o2d_core_133;
  assign popcount47_8o2d_core_145 = input_a[7] ^ popcount47_8o2d_core_141;
  assign popcount47_8o2d_core_146 = popcount47_8o2d_core_135 & popcount47_8o2d_core_141;
  assign popcount47_8o2d_core_147 = popcount47_8o2d_core_145 ^ popcount47_8o2d_core_144;
  assign popcount47_8o2d_core_148 = popcount47_8o2d_core_145 & popcount47_8o2d_core_144;
  assign popcount47_8o2d_core_149 = popcount47_8o2d_core_146 | popcount47_8o2d_core_148;
  assign popcount47_8o2d_core_150 = popcount47_8o2d_core_136 ^ popcount47_8o2d_core_142;
  assign popcount47_8o2d_core_151 = popcount47_8o2d_core_136 & popcount47_8o2d_core_142;
  assign popcount47_8o2d_core_152 = popcount47_8o2d_core_150 ^ popcount47_8o2d_core_149;
  assign popcount47_8o2d_core_153 = popcount47_8o2d_core_150 & popcount47_8o2d_core_149;
  assign popcount47_8o2d_core_154 = popcount47_8o2d_core_151 | popcount47_8o2d_core_153;
  assign popcount47_8o2d_core_157 = popcount47_8o2d_core_123 ^ popcount47_8o2d_core_147;
  assign popcount47_8o2d_core_158 = popcount47_8o2d_core_123 & popcount47_8o2d_core_147;
  assign popcount47_8o2d_core_162 = popcount47_8o2d_core_128 ^ popcount47_8o2d_core_152;
  assign popcount47_8o2d_core_163 = popcount47_8o2d_core_128 & popcount47_8o2d_core_152;
  assign popcount47_8o2d_core_164 = popcount47_8o2d_core_162 ^ popcount47_8o2d_core_158;
  assign popcount47_8o2d_core_165 = popcount47_8o2d_core_162 & popcount47_8o2d_core_158;
  assign popcount47_8o2d_core_166 = popcount47_8o2d_core_163 | popcount47_8o2d_core_165;
  assign popcount47_8o2d_core_167 = popcount47_8o2d_core_130 ^ popcount47_8o2d_core_154;
  assign popcount47_8o2d_core_168 = popcount47_8o2d_core_130 & popcount47_8o2d_core_154;
  assign popcount47_8o2d_core_169 = popcount47_8o2d_core_167 ^ popcount47_8o2d_core_166;
  assign popcount47_8o2d_core_170 = popcount47_8o2d_core_167 & popcount47_8o2d_core_166;
  assign popcount47_8o2d_core_171 = popcount47_8o2d_core_168 | popcount47_8o2d_core_170;
  assign popcount47_8o2d_core_172_not = ~popcount47_8o2d_core_090_not;
  assign popcount47_8o2d_core_174 = popcount47_8o2d_core_094 ^ popcount47_8o2d_core_157;
  assign popcount47_8o2d_core_175 = popcount47_8o2d_core_094 & popcount47_8o2d_core_157;
  assign popcount47_8o2d_core_176 = popcount47_8o2d_core_174 ^ input_a[38];
  assign popcount47_8o2d_core_177 = popcount47_8o2d_core_174 & input_a[38];
  assign popcount47_8o2d_core_178 = popcount47_8o2d_core_175 | input_a[6];
  assign popcount47_8o2d_core_179 = popcount47_8o2d_core_099 ^ popcount47_8o2d_core_164;
  assign popcount47_8o2d_core_180 = popcount47_8o2d_core_099 & popcount47_8o2d_core_164;
  assign popcount47_8o2d_core_181 = popcount47_8o2d_core_179 ^ popcount47_8o2d_core_178;
  assign popcount47_8o2d_core_182 = popcount47_8o2d_core_179 & popcount47_8o2d_core_178;
  assign popcount47_8o2d_core_183 = popcount47_8o2d_core_180 | popcount47_8o2d_core_182;
  assign popcount47_8o2d_core_184 = popcount47_8o2d_core_104 ^ popcount47_8o2d_core_169;
  assign popcount47_8o2d_core_185 = popcount47_8o2d_core_104 & popcount47_8o2d_core_169;
  assign popcount47_8o2d_core_186 = popcount47_8o2d_core_184 ^ popcount47_8o2d_core_183;
  assign popcount47_8o2d_core_187 = popcount47_8o2d_core_184 & popcount47_8o2d_core_183;
  assign popcount47_8o2d_core_188 = popcount47_8o2d_core_185 | popcount47_8o2d_core_187;
  assign popcount47_8o2d_core_189 = popcount47_8o2d_core_105 ^ popcount47_8o2d_core_171;
  assign popcount47_8o2d_core_190 = popcount47_8o2d_core_105 & popcount47_8o2d_core_171;
  assign popcount47_8o2d_core_191 = popcount47_8o2d_core_189 ^ popcount47_8o2d_core_188;
  assign popcount47_8o2d_core_192 = popcount47_8o2d_core_189 & popcount47_8o2d_core_188;
  assign popcount47_8o2d_core_193 = popcount47_8o2d_core_190 | popcount47_8o2d_core_192;
  assign popcount47_8o2d_core_194 = input_a[24] ^ input_a[24];
  assign popcount47_8o2d_core_195 = input_a[24] & input_a[25];
  assign popcount47_8o2d_core_196 = input_a[23] ^ popcount47_8o2d_core_194;
  assign popcount47_8o2d_core_197 = input_a[23] & popcount47_8o2d_core_194;
  assign popcount47_8o2d_core_198 = popcount47_8o2d_core_195 & popcount47_8o2d_core_197;
  assign popcount47_8o2d_core_199 = popcount47_8o2d_core_195 & input_a[36];
  assign popcount47_8o2d_core_200 = input_a[27] ^ input_a[28];
  assign popcount47_8o2d_core_201 = input_a[27] & input_a[28];
  assign popcount47_8o2d_core_202 = input_a[26] ^ popcount47_8o2d_core_200;
  assign popcount47_8o2d_core_203 = input_a[26] & popcount47_8o2d_core_200;
  assign popcount47_8o2d_core_204 = popcount47_8o2d_core_201 ^ popcount47_8o2d_core_203;
  assign popcount47_8o2d_core_205 = popcount47_8o2d_core_201 & popcount47_8o2d_core_203;
  assign popcount47_8o2d_core_206 = popcount47_8o2d_core_196 ^ input_a[29];
  assign popcount47_8o2d_core_207 = popcount47_8o2d_core_196 & popcount47_8o2d_core_202;
  assign popcount47_8o2d_core_208 = popcount47_8o2d_core_198 ^ popcount47_8o2d_core_204;
  assign popcount47_8o2d_core_209 = popcount47_8o2d_core_198 & popcount47_8o2d_core_204;
  assign popcount47_8o2d_core_210 = popcount47_8o2d_core_208 ^ popcount47_8o2d_core_207;
  assign popcount47_8o2d_core_211 = popcount47_8o2d_core_208 & popcount47_8o2d_core_207;
  assign popcount47_8o2d_core_212 = popcount47_8o2d_core_209 | popcount47_8o2d_core_211;
  assign popcount47_8o2d_core_213 = popcount47_8o2d_core_199 ^ popcount47_8o2d_core_205;
  assign popcount47_8o2d_core_214 = popcount47_8o2d_core_199 & popcount47_8o2d_core_205;
  assign popcount47_8o2d_core_215 = popcount47_8o2d_core_213 ^ popcount47_8o2d_core_212;
  assign popcount47_8o2d_core_216 = popcount47_8o2d_core_213 & popcount47_8o2d_core_212;
  assign popcount47_8o2d_core_217 = popcount47_8o2d_core_214 | popcount47_8o2d_core_216;
  assign popcount47_8o2d_core_218 = input_a[30] ^ input_a[31];
  assign popcount47_8o2d_core_219 = input_a[30] & input_a[31];
  assign popcount47_8o2d_core_220 = input_a[29] ^ popcount47_8o2d_core_218;
  assign popcount47_8o2d_core_221 = input_a[29] & popcount47_8o2d_core_218;
  assign popcount47_8o2d_core_222 = popcount47_8o2d_core_219 ^ popcount47_8o2d_core_221;
  assign popcount47_8o2d_core_223 = popcount47_8o2d_core_219 & popcount47_8o2d_core_221;
  assign popcount47_8o2d_core_224 = input_a[33] ^ input_a[34];
  assign popcount47_8o2d_core_225 = input_a[33] & input_a[34];
  assign popcount47_8o2d_core_226 = input_a[32] ^ popcount47_8o2d_core_224;
  assign popcount47_8o2d_core_227 = input_a[15] & popcount47_8o2d_core_224;
  assign popcount47_8o2d_core_228 = popcount47_8o2d_core_225 & input_a[24];
  assign popcount47_8o2d_core_229 = popcount47_8o2d_core_225 & popcount47_8o2d_core_227;
  assign popcount47_8o2d_core_230 = popcount47_8o2d_core_220 ^ popcount47_8o2d_core_226;
  assign popcount47_8o2d_core_231 = popcount47_8o2d_core_220 & popcount47_8o2d_core_226;
  assign popcount47_8o2d_core_232 = popcount47_8o2d_core_222 ^ popcount47_8o2d_core_228;
  assign popcount47_8o2d_core_233 = popcount47_8o2d_core_222 & popcount47_8o2d_core_228;
  assign popcount47_8o2d_core_234 = popcount47_8o2d_core_232 ^ popcount47_8o2d_core_231;
  assign popcount47_8o2d_core_235 = popcount47_8o2d_core_232 & popcount47_8o2d_core_231;
  assign popcount47_8o2d_core_236 = popcount47_8o2d_core_233 | popcount47_8o2d_core_235;
  assign popcount47_8o2d_core_237 = popcount47_8o2d_core_223 ^ popcount47_8o2d_core_229;
  assign popcount47_8o2d_core_239 = popcount47_8o2d_core_237 ^ popcount47_8o2d_core_236;
  assign popcount47_8o2d_core_240 = popcount47_8o2d_core_237 & popcount47_8o2d_core_236;
  assign popcount47_8o2d_core_242 = popcount47_8o2d_core_206 ^ popcount47_8o2d_core_230;
  assign popcount47_8o2d_core_243 = popcount47_8o2d_core_206 & popcount47_8o2d_core_230;
  assign popcount47_8o2d_core_244 = popcount47_8o2d_core_210 ^ popcount47_8o2d_core_234;
  assign popcount47_8o2d_core_245 = popcount47_8o2d_core_210 & popcount47_8o2d_core_234;
  assign popcount47_8o2d_core_249 = popcount47_8o2d_core_215 & popcount47_8o2d_core_239;
  assign popcount47_8o2d_core_250 = popcount47_8o2d_core_215 & popcount47_8o2d_core_239;
  assign popcount47_8o2d_core_256 = popcount47_8o2d_core_217 ^ popcount47_8o2d_core_250;
  assign popcount47_8o2d_core_257 = popcount47_8o2d_core_217 & popcount47_8o2d_core_250;
  assign popcount47_8o2d_core_259 = input_a[36] ^ input_a[37];
  assign popcount47_8o2d_core_260 = input_a[36] & input_a[37];
  assign popcount47_8o2d_core_261 = input_a[38] ^ popcount47_8o2d_core_259;
  assign popcount47_8o2d_core_266 = input_a[39] & input_a[40];
  assign popcount47_8o2d_core_267 = input_a[38] ^ input_a[39];
  assign popcount47_8o2d_core_268 = input_a[38] & input_a[25];
  assign popcount47_8o2d_core_269 = popcount47_8o2d_core_266 ^ popcount47_8o2d_core_268;
  assign popcount47_8o2d_core_270 = popcount47_8o2d_core_266 & popcount47_8o2d_core_268;
  assign popcount47_8o2d_core_271 = popcount47_8o2d_core_261 ^ popcount47_8o2d_core_267;
  assign popcount47_8o2d_core_272 = popcount47_8o2d_core_261 & popcount47_8o2d_core_267;
  assign popcount47_8o2d_core_273 = popcount47_8o2d_core_260 ^ popcount47_8o2d_core_269;
  assign popcount47_8o2d_core_274 = popcount47_8o2d_core_260 & popcount47_8o2d_core_269;
  assign popcount47_8o2d_core_276 = popcount47_8o2d_core_273 & popcount47_8o2d_core_272;
  assign popcount47_8o2d_core_277 = popcount47_8o2d_core_274 | popcount47_8o2d_core_276;
  assign popcount47_8o2d_core_280 = popcount47_8o2d_core_270 ^ popcount47_8o2d_core_277;
  assign popcount47_8o2d_core_281 = popcount47_8o2d_core_270 & popcount47_8o2d_core_277;
  assign popcount47_8o2d_core_283 = input_a[42] ^ input_a[43];
  assign popcount47_8o2d_core_284 = ~(input_a[42] & input_a[43]);
  assign popcount47_8o2d_core_285 = input_a[41] ^ input_a[31];
  assign popcount47_8o2d_core_287 = popcount47_8o2d_core_284 ^ input_a[41];
  assign popcount47_8o2d_core_288 = popcount47_8o2d_core_284 & input_a[41];
  assign popcount47_8o2d_core_289 = input_a[45] ^ input_a[46];
  assign popcount47_8o2d_core_290 = input_a[23] & input_a[46];
  assign popcount47_8o2d_core_291 = input_a[44] ^ popcount47_8o2d_core_289;
  assign popcount47_8o2d_core_292 = input_a[44] & popcount47_8o2d_core_289;
  assign popcount47_8o2d_core_293 = popcount47_8o2d_core_290 ^ popcount47_8o2d_core_292;
  assign popcount47_8o2d_core_294 = popcount47_8o2d_core_290 & popcount47_8o2d_core_292;
  assign popcount47_8o2d_core_295 = popcount47_8o2d_core_285 ^ popcount47_8o2d_core_291;
  assign popcount47_8o2d_core_296 = popcount47_8o2d_core_285 & popcount47_8o2d_core_291;
  assign popcount47_8o2d_core_297 = popcount47_8o2d_core_287 ^ popcount47_8o2d_core_293;
  assign popcount47_8o2d_core_298 = popcount47_8o2d_core_287 & popcount47_8o2d_core_293;
  assign popcount47_8o2d_core_299 = popcount47_8o2d_core_297 ^ popcount47_8o2d_core_296;
  assign popcount47_8o2d_core_302 = popcount47_8o2d_core_288 ^ popcount47_8o2d_core_294;
  assign popcount47_8o2d_core_303 = popcount47_8o2d_core_288 & popcount47_8o2d_core_294;
  assign popcount47_8o2d_core_304 = popcount47_8o2d_core_302 ^ popcount47_8o2d_core_298;
  assign popcount47_8o2d_core_305 = popcount47_8o2d_core_302 & popcount47_8o2d_core_298;
  assign popcount47_8o2d_core_306 = popcount47_8o2d_core_303 | popcount47_8o2d_core_305;
  assign popcount47_8o2d_core_307 = input_a[31] ^ popcount47_8o2d_core_295;
  assign popcount47_8o2d_core_308 = popcount47_8o2d_core_271 & popcount47_8o2d_core_295;
  assign popcount47_8o2d_core_311 = popcount47_8o2d_core_299 ^ popcount47_8o2d_core_308;
  assign popcount47_8o2d_core_312 = popcount47_8o2d_core_299 & popcount47_8o2d_core_308;
  assign popcount47_8o2d_core_314 = popcount47_8o2d_core_280 ^ popcount47_8o2d_core_304;
  assign popcount47_8o2d_core_315 = popcount47_8o2d_core_280 & popcount47_8o2d_core_304;
  assign popcount47_8o2d_core_316 = popcount47_8o2d_core_314 ^ popcount47_8o2d_core_312;
  assign popcount47_8o2d_core_317 = popcount47_8o2d_core_314 & popcount47_8o2d_core_312;
  assign popcount47_8o2d_core_318 = popcount47_8o2d_core_315 | popcount47_8o2d_core_317;
  assign popcount47_8o2d_core_319 = popcount47_8o2d_core_281 ^ popcount47_8o2d_core_306;
  assign popcount47_8o2d_core_320 = popcount47_8o2d_core_281 & popcount47_8o2d_core_306;
  assign popcount47_8o2d_core_321 = popcount47_8o2d_core_319 ^ popcount47_8o2d_core_318;
  assign popcount47_8o2d_core_322 = popcount47_8o2d_core_319 & popcount47_8o2d_core_318;
  assign popcount47_8o2d_core_323 = popcount47_8o2d_core_320 | popcount47_8o2d_core_322;
  assign popcount47_8o2d_core_324 = popcount47_8o2d_core_242 ^ popcount47_8o2d_core_307;
  assign popcount47_8o2d_core_325 = popcount47_8o2d_core_242 & popcount47_8o2d_core_307;
  assign popcount47_8o2d_core_328 = input_a[16] ^ popcount47_8o2d_core_325;
  assign popcount47_8o2d_core_329 = popcount47_8o2d_core_311 & popcount47_8o2d_core_325;
  assign popcount47_8o2d_core_331 = popcount47_8o2d_core_249 ^ popcount47_8o2d_core_316;
  assign popcount47_8o2d_core_332 = popcount47_8o2d_core_249 & popcount47_8o2d_core_316;
  assign popcount47_8o2d_core_333 = popcount47_8o2d_core_331 ^ popcount47_8o2d_core_329;
  assign popcount47_8o2d_core_334 = popcount47_8o2d_core_331 & popcount47_8o2d_core_329;
  assign popcount47_8o2d_core_335 = popcount47_8o2d_core_332 | popcount47_8o2d_core_334;
  assign popcount47_8o2d_core_336 = popcount47_8o2d_core_256 ^ popcount47_8o2d_core_321;
  assign popcount47_8o2d_core_337 = popcount47_8o2d_core_256 & popcount47_8o2d_core_321;
  assign popcount47_8o2d_core_338 = popcount47_8o2d_core_336 ^ popcount47_8o2d_core_335;
  assign popcount47_8o2d_core_339 = popcount47_8o2d_core_336 & popcount47_8o2d_core_335;
  assign popcount47_8o2d_core_340 = popcount47_8o2d_core_337 | popcount47_8o2d_core_339;
  assign popcount47_8o2d_core_341 = popcount47_8o2d_core_257 ^ popcount47_8o2d_core_323;
  assign popcount47_8o2d_core_342 = popcount47_8o2d_core_257 & popcount47_8o2d_core_323;
  assign popcount47_8o2d_core_343 = popcount47_8o2d_core_341 ^ popcount47_8o2d_core_340;
  assign popcount47_8o2d_core_344 = popcount47_8o2d_core_341 & popcount47_8o2d_core_340;
  assign popcount47_8o2d_core_345 = popcount47_8o2d_core_342 | popcount47_8o2d_core_344;
  assign popcount47_8o2d_core_346 = popcount47_8o2d_core_172_not ^ popcount47_8o2d_core_324;
  assign popcount47_8o2d_core_347 = popcount47_8o2d_core_172_not & popcount47_8o2d_core_324;
  assign popcount47_8o2d_core_348 = popcount47_8o2d_core_176 ^ popcount47_8o2d_core_328;
  assign popcount47_8o2d_core_349 = input_a[29] & popcount47_8o2d_core_328;
  assign popcount47_8o2d_core_350 = popcount47_8o2d_core_348 ^ popcount47_8o2d_core_347;
  assign popcount47_8o2d_core_353 = popcount47_8o2d_core_181 ^ popcount47_8o2d_core_333;
  assign popcount47_8o2d_core_354 = popcount47_8o2d_core_181 & popcount47_8o2d_core_333;
  assign popcount47_8o2d_core_355_not = ~popcount47_8o2d_core_353;
  assign popcount47_8o2d_core_357 = popcount47_8o2d_core_354 | popcount47_8o2d_core_353;
  assign popcount47_8o2d_core_358 = popcount47_8o2d_core_186 ^ popcount47_8o2d_core_338;
  assign popcount47_8o2d_core_359 = popcount47_8o2d_core_186 & popcount47_8o2d_core_338;
  assign popcount47_8o2d_core_360 = popcount47_8o2d_core_358 ^ popcount47_8o2d_core_357;
  assign popcount47_8o2d_core_361 = popcount47_8o2d_core_358 & popcount47_8o2d_core_357;
  assign popcount47_8o2d_core_362 = popcount47_8o2d_core_359 | popcount47_8o2d_core_361;
  assign popcount47_8o2d_core_363 = popcount47_8o2d_core_191 ^ popcount47_8o2d_core_343;
  assign popcount47_8o2d_core_364 = popcount47_8o2d_core_191 & popcount47_8o2d_core_343;
  assign popcount47_8o2d_core_365 = popcount47_8o2d_core_363 ^ popcount47_8o2d_core_362;
  assign popcount47_8o2d_core_366 = popcount47_8o2d_core_363 & popcount47_8o2d_core_362;
  assign popcount47_8o2d_core_367 = popcount47_8o2d_core_364 | popcount47_8o2d_core_366;
  assign popcount47_8o2d_core_368 = popcount47_8o2d_core_193 ^ popcount47_8o2d_core_345;
  assign popcount47_8o2d_core_369 = popcount47_8o2d_core_193 & popcount47_8o2d_core_345;
  assign popcount47_8o2d_core_370 = popcount47_8o2d_core_368 ^ popcount47_8o2d_core_367;
  assign popcount47_8o2d_core_371 = popcount47_8o2d_core_368 & popcount47_8o2d_core_367;
  assign popcount47_8o2d_core_372 = ~(popcount47_8o2d_core_369 & popcount47_8o2d_core_371);

  assign popcount47_8o2d_out[0] = popcount47_8o2d_core_346;
  assign popcount47_8o2d_out[1] = popcount47_8o2d_core_350;
  assign popcount47_8o2d_out[2] = popcount47_8o2d_core_355_not;
  assign popcount47_8o2d_out[3] = popcount47_8o2d_core_360;
  assign popcount47_8o2d_out[4] = popcount47_8o2d_core_365;
  assign popcount47_8o2d_out[5] = popcount47_8o2d_core_370;
endmodule