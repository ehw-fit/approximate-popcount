// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.43927
// WCE=8.0
// EP=0.785115%
// Printed PDK parameters:
//  Area=36827327.0
//  Delay=64766356.0
//  Power=1989400.0

module popcount29_b8e8(input [28:0] input_a, output [4:0] popcount29_b8e8_out);
  wire popcount29_b8e8_core_031;
  wire popcount29_b8e8_core_033;
  wire popcount29_b8e8_core_037;
  wire popcount29_b8e8_core_038;
  wire popcount29_b8e8_core_041;
  wire popcount29_b8e8_core_044;
  wire popcount29_b8e8_core_045_not;
  wire popcount29_b8e8_core_047;
  wire popcount29_b8e8_core_048;
  wire popcount29_b8e8_core_049;
  wire popcount29_b8e8_core_053;
  wire popcount29_b8e8_core_054;
  wire popcount29_b8e8_core_055;
  wire popcount29_b8e8_core_059;
  wire popcount29_b8e8_core_061;
  wire popcount29_b8e8_core_062;
  wire popcount29_b8e8_core_063;
  wire popcount29_b8e8_core_066;
  wire popcount29_b8e8_core_067;
  wire popcount29_b8e8_core_069;
  wire popcount29_b8e8_core_070;
  wire popcount29_b8e8_core_071;
  wire popcount29_b8e8_core_072;
  wire popcount29_b8e8_core_073;
  wire popcount29_b8e8_core_074;
  wire popcount29_b8e8_core_075;
  wire popcount29_b8e8_core_078;
  wire popcount29_b8e8_core_079;
  wire popcount29_b8e8_core_080;
  wire popcount29_b8e8_core_081;
  wire popcount29_b8e8_core_082;
  wire popcount29_b8e8_core_083;
  wire popcount29_b8e8_core_085;
  wire popcount29_b8e8_core_086;
  wire popcount29_b8e8_core_087;
  wire popcount29_b8e8_core_089;
  wire popcount29_b8e8_core_090;
  wire popcount29_b8e8_core_093;
  wire popcount29_b8e8_core_094;
  wire popcount29_b8e8_core_096_not;
  wire popcount29_b8e8_core_098;
  wire popcount29_b8e8_core_099;
  wire popcount29_b8e8_core_100;
  wire popcount29_b8e8_core_102;
  wire popcount29_b8e8_core_104;
  wire popcount29_b8e8_core_105;
  wire popcount29_b8e8_core_106;
  wire popcount29_b8e8_core_107;
  wire popcount29_b8e8_core_108;
  wire popcount29_b8e8_core_109;
  wire popcount29_b8e8_core_111;
  wire popcount29_b8e8_core_112;
  wire popcount29_b8e8_core_113;
  wire popcount29_b8e8_core_114;
  wire popcount29_b8e8_core_115;
  wire popcount29_b8e8_core_116;
  wire popcount29_b8e8_core_117;
  wire popcount29_b8e8_core_120;
  wire popcount29_b8e8_core_121;
  wire popcount29_b8e8_core_124;
  wire popcount29_b8e8_core_125;
  wire popcount29_b8e8_core_126;
  wire popcount29_b8e8_core_127;
  wire popcount29_b8e8_core_128;
  wire popcount29_b8e8_core_129;
  wire popcount29_b8e8_core_131;
  wire popcount29_b8e8_core_133;
  wire popcount29_b8e8_core_134;
  wire popcount29_b8e8_core_135;
  wire popcount29_b8e8_core_136;
  wire popcount29_b8e8_core_138;
  wire popcount29_b8e8_core_139;
  wire popcount29_b8e8_core_140;
  wire popcount29_b8e8_core_143;
  wire popcount29_b8e8_core_145;
  wire popcount29_b8e8_core_147;
  wire popcount29_b8e8_core_148;
  wire popcount29_b8e8_core_150;
  wire popcount29_b8e8_core_151;
  wire popcount29_b8e8_core_152;
  wire popcount29_b8e8_core_154;
  wire popcount29_b8e8_core_155;
  wire popcount29_b8e8_core_157;
  wire popcount29_b8e8_core_158;
  wire popcount29_b8e8_core_159;
  wire popcount29_b8e8_core_160;
  wire popcount29_b8e8_core_161;
  wire popcount29_b8e8_core_162;
  wire popcount29_b8e8_core_166;
  wire popcount29_b8e8_core_167;
  wire popcount29_b8e8_core_169;
  wire popcount29_b8e8_core_170;
  wire popcount29_b8e8_core_171;
  wire popcount29_b8e8_core_172;
  wire popcount29_b8e8_core_173;
  wire popcount29_b8e8_core_174;
  wire popcount29_b8e8_core_175;
  wire popcount29_b8e8_core_176;
  wire popcount29_b8e8_core_177;
  wire popcount29_b8e8_core_178;
  wire popcount29_b8e8_core_179;
  wire popcount29_b8e8_core_180;
  wire popcount29_b8e8_core_182;
  wire popcount29_b8e8_core_184;
  wire popcount29_b8e8_core_185;
  wire popcount29_b8e8_core_186;
  wire popcount29_b8e8_core_188;
  wire popcount29_b8e8_core_189;
  wire popcount29_b8e8_core_191;
  wire popcount29_b8e8_core_193;
  wire popcount29_b8e8_core_194;
  wire popcount29_b8e8_core_195;
  wire popcount29_b8e8_core_196;
  wire popcount29_b8e8_core_197;
  wire popcount29_b8e8_core_198;
  wire popcount29_b8e8_core_199;
  wire popcount29_b8e8_core_200;
  wire popcount29_b8e8_core_201;
  wire popcount29_b8e8_core_202;
  wire popcount29_b8e8_core_203;
  wire popcount29_b8e8_core_204;
  wire popcount29_b8e8_core_206;
  wire popcount29_b8e8_core_207;

  assign popcount29_b8e8_core_031 = input_a[0] & input_a[13];
  assign popcount29_b8e8_core_033 = ~(input_a[15] & input_a[25]);
  assign popcount29_b8e8_core_037 = ~input_a[24];
  assign popcount29_b8e8_core_038 = ~(input_a[13] & input_a[16]);
  assign popcount29_b8e8_core_041 = ~input_a[10];
  assign popcount29_b8e8_core_044 = ~(input_a[12] & input_a[7]);
  assign popcount29_b8e8_core_045_not = ~input_a[23];
  assign popcount29_b8e8_core_047 = input_a[10] | input_a[8];
  assign popcount29_b8e8_core_048 = ~(input_a[8] | input_a[10]);
  assign popcount29_b8e8_core_049 = ~input_a[7];
  assign popcount29_b8e8_core_053 = input_a[18] ^ input_a[27];
  assign popcount29_b8e8_core_054 = input_a[0] & input_a[28];
  assign popcount29_b8e8_core_055 = input_a[27] ^ input_a[13];
  assign popcount29_b8e8_core_059 = input_a[20] & input_a[24];
  assign popcount29_b8e8_core_061 = input_a[8] & input_a[15];
  assign popcount29_b8e8_core_062 = input_a[24] | input_a[4];
  assign popcount29_b8e8_core_063 = ~input_a[26];
  assign popcount29_b8e8_core_066 = ~(input_a[7] | input_a[5]);
  assign popcount29_b8e8_core_067 = input_a[10] & input_a[11];
  assign popcount29_b8e8_core_069 = input_a[26] & input_a[28];
  assign popcount29_b8e8_core_070 = ~(input_a[3] | input_a[23]);
  assign popcount29_b8e8_core_071 = input_a[16] & input_a[12];
  assign popcount29_b8e8_core_072 = popcount29_b8e8_core_067 ^ popcount29_b8e8_core_069;
  assign popcount29_b8e8_core_073 = popcount29_b8e8_core_067 & popcount29_b8e8_core_069;
  assign popcount29_b8e8_core_074 = popcount29_b8e8_core_072 | popcount29_b8e8_core_071;
  assign popcount29_b8e8_core_075 = ~input_a[4];
  assign popcount29_b8e8_core_078 = input_a[20] & input_a[7];
  assign popcount29_b8e8_core_079 = popcount29_b8e8_core_061 ^ popcount29_b8e8_core_074;
  assign popcount29_b8e8_core_080 = popcount29_b8e8_core_061 & popcount29_b8e8_core_074;
  assign popcount29_b8e8_core_081 = popcount29_b8e8_core_079 ^ popcount29_b8e8_core_078;
  assign popcount29_b8e8_core_082 = popcount29_b8e8_core_079 & popcount29_b8e8_core_078;
  assign popcount29_b8e8_core_083 = popcount29_b8e8_core_080 | popcount29_b8e8_core_082;
  assign popcount29_b8e8_core_085 = ~(input_a[1] | input_a[4]);
  assign popcount29_b8e8_core_086 = popcount29_b8e8_core_073 | popcount29_b8e8_core_083;
  assign popcount29_b8e8_core_087 = input_a[19] ^ input_a[12];
  assign popcount29_b8e8_core_089 = input_a[6] | input_a[28];
  assign popcount29_b8e8_core_090 = input_a[6] & input_a[14];
  assign popcount29_b8e8_core_093 = popcount29_b8e8_core_081 ^ popcount29_b8e8_core_090;
  assign popcount29_b8e8_core_094 = popcount29_b8e8_core_081 & popcount29_b8e8_core_090;
  assign popcount29_b8e8_core_096_not = ~popcount29_b8e8_core_086;
  assign popcount29_b8e8_core_098 = popcount29_b8e8_core_096_not ^ popcount29_b8e8_core_094;
  assign popcount29_b8e8_core_099 = input_a[14] & popcount29_b8e8_core_094;
  assign popcount29_b8e8_core_100 = popcount29_b8e8_core_086 | popcount29_b8e8_core_099;
  assign popcount29_b8e8_core_102 = ~(input_a[23] & input_a[2]);
  assign popcount29_b8e8_core_104 = ~(input_a[20] | input_a[0]);
  assign popcount29_b8e8_core_105 = ~(input_a[19] ^ input_a[9]);
  assign popcount29_b8e8_core_106 = input_a[17] & input_a[8];
  assign popcount29_b8e8_core_107 = input_a[22] & input_a[24];
  assign popcount29_b8e8_core_108 = ~input_a[24];
  assign popcount29_b8e8_core_109 = input_a[20] ^ input_a[4];
  assign popcount29_b8e8_core_111 = input_a[6] ^ input_a[28];
  assign popcount29_b8e8_core_112 = input_a[17] | input_a[18];
  assign popcount29_b8e8_core_113 = input_a[13] & input_a[5];
  assign popcount29_b8e8_core_114 = input_a[19] | input_a[4];
  assign popcount29_b8e8_core_115 = ~(input_a[3] ^ input_a[3]);
  assign popcount29_b8e8_core_116 = ~(input_a[14] | input_a[9]);
  assign popcount29_b8e8_core_117 = popcount29_b8e8_core_112 & popcount29_b8e8_core_114;
  assign popcount29_b8e8_core_120 = popcount29_b8e8_core_113 | popcount29_b8e8_core_117;
  assign popcount29_b8e8_core_121 = input_a[8] ^ input_a[8];
  assign popcount29_b8e8_core_124 = input_a[23] & input_a[21];
  assign popcount29_b8e8_core_125 = popcount29_b8e8_core_107 ^ popcount29_b8e8_core_120;
  assign popcount29_b8e8_core_126 = popcount29_b8e8_core_107 & popcount29_b8e8_core_120;
  assign popcount29_b8e8_core_127 = popcount29_b8e8_core_125 ^ popcount29_b8e8_core_124;
  assign popcount29_b8e8_core_128 = popcount29_b8e8_core_125 & popcount29_b8e8_core_124;
  assign popcount29_b8e8_core_129 = popcount29_b8e8_core_126 | popcount29_b8e8_core_128;
  assign popcount29_b8e8_core_131 = ~input_a[12];
  assign popcount29_b8e8_core_133 = input_a[13] ^ input_a[14];
  assign popcount29_b8e8_core_134 = ~(input_a[5] ^ input_a[13]);
  assign popcount29_b8e8_core_135 = input_a[20] & input_a[17];
  assign popcount29_b8e8_core_136 = input_a[25] | input_a[27];
  assign popcount29_b8e8_core_138 = input_a[23] ^ input_a[4];
  assign popcount29_b8e8_core_139 = input_a[18] ^ input_a[28];
  assign popcount29_b8e8_core_140 = ~(input_a[5] | input_a[0]);
  assign popcount29_b8e8_core_143 = input_a[25] | input_a[0];
  assign popcount29_b8e8_core_145 = ~input_a[28];
  assign popcount29_b8e8_core_147 = ~(input_a[2] ^ input_a[12]);
  assign popcount29_b8e8_core_148 = input_a[21] & input_a[7];
  assign popcount29_b8e8_core_150 = ~(input_a[4] | input_a[5]);
  assign popcount29_b8e8_core_151 = ~(input_a[21] | input_a[23]);
  assign popcount29_b8e8_core_152 = input_a[1] & input_a[24];
  assign popcount29_b8e8_core_154 = input_a[2] | input_a[27];
  assign popcount29_b8e8_core_155 = input_a[12] | input_a[17];
  assign popcount29_b8e8_core_157 = ~(input_a[1] | input_a[12]);
  assign popcount29_b8e8_core_158 = ~(input_a[9] & input_a[15]);
  assign popcount29_b8e8_core_159 = ~(popcount29_b8e8_core_143 & popcount29_b8e8_core_154);
  assign popcount29_b8e8_core_160 = popcount29_b8e8_core_143 & popcount29_b8e8_core_154;
  assign popcount29_b8e8_core_161 = popcount29_b8e8_core_159 ^ input_a[9];
  assign popcount29_b8e8_core_162 = input_a[4] ^ input_a[8];
  assign popcount29_b8e8_core_166 = input_a[9] | popcount29_b8e8_core_160;
  assign popcount29_b8e8_core_167 = ~input_a[18];
  assign popcount29_b8e8_core_169 = input_a[28] | input_a[7];
  assign popcount29_b8e8_core_170 = input_a[1] & input_a[3];
  assign popcount29_b8e8_core_171 = popcount29_b8e8_core_127 ^ popcount29_b8e8_core_161;
  assign popcount29_b8e8_core_172 = popcount29_b8e8_core_127 & popcount29_b8e8_core_161;
  assign popcount29_b8e8_core_173 = popcount29_b8e8_core_171 ^ popcount29_b8e8_core_170;
  assign popcount29_b8e8_core_174 = popcount29_b8e8_core_171 & popcount29_b8e8_core_170;
  assign popcount29_b8e8_core_175 = popcount29_b8e8_core_172 | popcount29_b8e8_core_174;
  assign popcount29_b8e8_core_176 = popcount29_b8e8_core_129 ^ popcount29_b8e8_core_166;
  assign popcount29_b8e8_core_177 = popcount29_b8e8_core_129 & popcount29_b8e8_core_166;
  assign popcount29_b8e8_core_178 = popcount29_b8e8_core_176 ^ popcount29_b8e8_core_175;
  assign popcount29_b8e8_core_179 = popcount29_b8e8_core_176 & popcount29_b8e8_core_175;
  assign popcount29_b8e8_core_180 = popcount29_b8e8_core_177 | popcount29_b8e8_core_179;
  assign popcount29_b8e8_core_182 = input_a[23] | input_a[23];
  assign popcount29_b8e8_core_184 = ~(input_a[2] | input_a[26]);
  assign popcount29_b8e8_core_185 = ~(input_a[25] & input_a[22]);
  assign popcount29_b8e8_core_186 = input_a[23] | input_a[7];
  assign popcount29_b8e8_core_188 = popcount29_b8e8_core_093 ^ popcount29_b8e8_core_173;
  assign popcount29_b8e8_core_189 = popcount29_b8e8_core_093 & popcount29_b8e8_core_173;
  assign popcount29_b8e8_core_191 = ~input_a[26];
  assign popcount29_b8e8_core_193 = popcount29_b8e8_core_098 ^ popcount29_b8e8_core_178;
  assign popcount29_b8e8_core_194 = popcount29_b8e8_core_098 & popcount29_b8e8_core_178;
  assign popcount29_b8e8_core_195 = popcount29_b8e8_core_193 ^ popcount29_b8e8_core_189;
  assign popcount29_b8e8_core_196 = popcount29_b8e8_core_193 & popcount29_b8e8_core_189;
  assign popcount29_b8e8_core_197 = popcount29_b8e8_core_194 | popcount29_b8e8_core_196;
  assign popcount29_b8e8_core_198 = popcount29_b8e8_core_100 ^ popcount29_b8e8_core_180;
  assign popcount29_b8e8_core_199 = popcount29_b8e8_core_100 & popcount29_b8e8_core_180;
  assign popcount29_b8e8_core_200 = popcount29_b8e8_core_198 ^ popcount29_b8e8_core_197;
  assign popcount29_b8e8_core_201 = popcount29_b8e8_core_198 & popcount29_b8e8_core_197;
  assign popcount29_b8e8_core_202 = popcount29_b8e8_core_199 | popcount29_b8e8_core_201;
  assign popcount29_b8e8_core_203 = ~(input_a[3] ^ input_a[18]);
  assign popcount29_b8e8_core_204 = ~(input_a[3] ^ input_a[11]);
  assign popcount29_b8e8_core_206 = input_a[9] ^ input_a[23];
  assign popcount29_b8e8_core_207 = input_a[9] | input_a[21];

  assign popcount29_b8e8_out[0] = popcount29_b8e8_core_200;
  assign popcount29_b8e8_out[1] = popcount29_b8e8_core_188;
  assign popcount29_b8e8_out[2] = popcount29_b8e8_core_195;
  assign popcount29_b8e8_out[3] = popcount29_b8e8_core_200;
  assign popcount29_b8e8_out[4] = popcount29_b8e8_core_202;
endmodule