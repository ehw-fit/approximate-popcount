
module cmp_pos(input [44:0] input_a, output [5:0] cgp_out);
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_061;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_101;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_111;
  wire cgp_core_114;
  wire cgp_core_115;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_118;
  wire cgp_core_119;
  wire cgp_core_121;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_129;
  wire cgp_core_131;
  wire cgp_core_132;
  wire cgp_core_135;
  wire cgp_core_138;
  wire cgp_core_139;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_147;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_150;
  wire cgp_core_151;
  wire cgp_core_152;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_162;
  wire cgp_core_164;
  wire cgp_core_165;
  wire cgp_core_166;
  wire cgp_core_167;
  wire cgp_core_168;
  wire cgp_core_169;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_181;
  wire cgp_core_183;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_188;
  wire cgp_core_189;
  wire cgp_core_191;
  wire cgp_core_194;
  wire cgp_core_197;
  wire cgp_core_198;
  wire cgp_core_199;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_203;
  wire cgp_core_204;
  wire cgp_core_205;
  wire cgp_core_207;
  wire cgp_core_208;
  wire cgp_core_209;
  wire cgp_core_210;
  wire cgp_core_211;
  wire cgp_core_212;
  wire cgp_core_214;
  wire cgp_core_215;
  wire cgp_core_218;
  wire cgp_core_219;
  wire cgp_core_222;
  wire cgp_core_225;
  wire cgp_core_226;
  wire cgp_core_227;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_230;
  wire cgp_core_231;
  wire cgp_core_232;
  wire cgp_core_235;
  wire cgp_core_236;
  wire cgp_core_237;
  wire cgp_core_238;
  wire cgp_core_239;
  wire cgp_core_241;
  wire cgp_core_242;
  wire cgp_core_243;
  wire cgp_core_244;
  wire cgp_core_246;
  wire cgp_core_247;
  wire cgp_core_248;
  wire cgp_core_250;
  wire cgp_core_252;
  wire cgp_core_254;
  wire cgp_core_255;
  wire cgp_core_256;
  wire cgp_core_258;
  wire cgp_core_260;
  wire cgp_core_261;
  wire cgp_core_262;
  wire cgp_core_263;
  wire cgp_core_266;
  wire cgp_core_267;
  wire cgp_core_268;
  wire cgp_core_269;
  wire cgp_core_272;
  wire cgp_core_273;
  wire cgp_core_274;
  wire cgp_core_275;
  wire cgp_core_276;
  wire cgp_core_277;
  wire cgp_core_278;
  wire cgp_core_279;
  wire cgp_core_280;
  wire cgp_core_282;
  wire cgp_core_286;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_291;
  wire cgp_core_293;
  wire cgp_core_294;
  wire cgp_core_296;
  wire cgp_core_301;
  wire cgp_core_303;
  wire cgp_core_304;
  wire cgp_core_306;
  wire cgp_core_308;
  wire cgp_core_309;
  wire cgp_core_310;
  wire cgp_core_311;
  wire cgp_core_312;
  wire cgp_core_313;
  wire cgp_core_314;
  wire cgp_core_315;
  wire cgp_core_316;
  wire cgp_core_317;
  wire cgp_core_318;
  wire cgp_core_319;
  wire cgp_core_322;
  wire cgp_core_328;
  wire cgp_core_329;
  wire cgp_core_330;
  wire cgp_core_331;
  wire cgp_core_332;
  wire cgp_core_333;
  wire cgp_core_334;
  wire cgp_core_335;
  wire cgp_core_336;
  wire cgp_core_337;
  wire cgp_core_338;
  wire cgp_core_339;
  wire cgp_core_340;
  wire cgp_core_341;
  wire cgp_core_342;
  wire cgp_core_343;
  wire cgp_core_344;
  wire cgp_core_345;
  wire cgp_core_346;
  wire cgp_core_347;
  wire cgp_core_348;
  wire cgp_core_349;
  wire cgp_core_350;
  wire cgp_core_351;
  wire cgp_core_352;
  wire cgp_core_354;
  wire cgp_core_355;

  assign cgp_core_049 = ~input_a[0];
  assign cgp_core_050 = input_a[43] & input_a[37];
  assign cgp_core_051 = input_a[17] & input_a[2];
  assign cgp_core_052 = input_a[44] & input_a[39];
  assign cgp_core_053 = cgp_core_050 | cgp_core_052;
  assign cgp_core_054 = ~input_a[35];
  assign cgp_core_055 = input_a[11] | input_a[37];
  assign cgp_core_056 = ~(input_a[0] ^ input_a[10]);
  assign cgp_core_061 = input_a[39] & input_a[30];
  assign cgp_core_063 = input_a[38] ^ input_a[15];
  assign cgp_core_065 = input_a[6] & input_a[7];
  assign cgp_core_067 = input_a[2] & input_a[36];
  assign cgp_core_068 = cgp_core_065 | cgp_core_067;
  assign cgp_core_070 = input_a[9] ^ input_a[10];
  assign cgp_core_071 = input_a[9] & input_a[10];
  assign cgp_core_072 = input_a[8] ^ cgp_core_070;
  assign cgp_core_073 = input_a[8] & cgp_core_070;
  assign cgp_core_074 = cgp_core_071 | cgp_core_073;
  assign cgp_core_076 = ~(input_a[40] | input_a[6]);
  assign cgp_core_077 = input_a[1] & cgp_core_072;
  assign cgp_core_078 = cgp_core_068 ^ cgp_core_074;
  assign cgp_core_079 = cgp_core_068 & cgp_core_074;
  assign cgp_core_080 = cgp_core_078 ^ cgp_core_077;
  assign cgp_core_081 = cgp_core_078 & cgp_core_077;
  assign cgp_core_082 = cgp_core_079 | cgp_core_081;
  assign cgp_core_084 = input_a[28] & input_a[44];
  assign cgp_core_087 = ~(input_a[18] & input_a[17]);
  assign cgp_core_088 = input_a[10] & input_a[26];
  assign cgp_core_089 = input_a[29] & input_a[18];
  assign cgp_core_090 = cgp_core_053 ^ cgp_core_080;
  assign cgp_core_091 = cgp_core_053 & cgp_core_080;
  assign cgp_core_092 = cgp_core_090 ^ cgp_core_089;
  assign cgp_core_093 = cgp_core_090 & cgp_core_089;
  assign cgp_core_094 = cgp_core_091 | cgp_core_093;
  assign cgp_core_097 = cgp_core_082 ^ cgp_core_094;
  assign cgp_core_098 = cgp_core_082 & cgp_core_094;
  assign cgp_core_101 = ~(input_a[36] & input_a[33]);
  assign cgp_core_103 = input_a[9] | input_a[27];
  assign cgp_core_104 = input_a[27] | input_a[16];
  assign cgp_core_105 = input_a[11] ^ input_a[12];
  assign cgp_core_106 = input_a[11] & input_a[12];
  assign cgp_core_107 = input_a[14] ^ input_a[15];
  assign cgp_core_108 = input_a[14] & input_a[15];
  assign cgp_core_109 = input_a[13] ^ cgp_core_107;
  assign cgp_core_110 = input_a[13] & cgp_core_107;
  assign cgp_core_111 = cgp_core_108 | cgp_core_110;
  assign cgp_core_114 = cgp_core_105 & cgp_core_109;
  assign cgp_core_115 = cgp_core_106 ^ cgp_core_111;
  assign cgp_core_116 = cgp_core_106 & cgp_core_111;
  assign cgp_core_117 = cgp_core_115 ^ cgp_core_114;
  assign cgp_core_118 = cgp_core_115 & cgp_core_114;
  assign cgp_core_119 = cgp_core_116 | cgp_core_118;
  assign cgp_core_121 = ~input_a[30];
  assign cgp_core_123 = ~input_a[36];
  assign cgp_core_124 = input_a[25] ^ input_a[7];
  assign cgp_core_127 = input_a[14] ^ input_a[6];
  assign cgp_core_128 = input_a[20] | input_a[21];
  assign cgp_core_129 = input_a[20] & input_a[21];
  assign cgp_core_131 = input_a[19] & cgp_core_128;
  assign cgp_core_132 = cgp_core_129 | cgp_core_131;
  assign cgp_core_135 = input_a[42] & input_a[24];
  assign cgp_core_138 = cgp_core_132 ^ cgp_core_135;
  assign cgp_core_139 = cgp_core_132 & cgp_core_135;
  assign cgp_core_144 = input_a[42] ^ input_a[23];
  assign cgp_core_145 = ~(input_a[24] | input_a[38]);
  assign cgp_core_147 = input_a[34] & input_a[25];
  assign cgp_core_148 = cgp_core_117 ^ cgp_core_138;
  assign cgp_core_149 = cgp_core_117 & cgp_core_138;
  assign cgp_core_150 = cgp_core_148 ^ cgp_core_147;
  assign cgp_core_151 = cgp_core_148 & cgp_core_147;
  assign cgp_core_152 = cgp_core_149 | cgp_core_151;
  assign cgp_core_153 = cgp_core_119 ^ cgp_core_139;
  assign cgp_core_154 = cgp_core_119 & cgp_core_139;
  assign cgp_core_155 = cgp_core_153 ^ cgp_core_152;
  assign cgp_core_156 = cgp_core_153 & cgp_core_152;
  assign cgp_core_157 = cgp_core_154 | cgp_core_156;
  assign cgp_core_162 = input_a[27] & input_a[19];
  assign cgp_core_164 = input_a[0] & input_a[40];
  assign cgp_core_165 = cgp_core_092 ^ cgp_core_150;
  assign cgp_core_166 = cgp_core_092 & cgp_core_150;
  assign cgp_core_167 = cgp_core_165 ^ cgp_core_164;
  assign cgp_core_168 = cgp_core_165 & cgp_core_164;
  assign cgp_core_169 = cgp_core_166 | cgp_core_168;
  assign cgp_core_170 = cgp_core_097 ^ cgp_core_155;
  assign cgp_core_171 = cgp_core_097 & cgp_core_155;
  assign cgp_core_172 = cgp_core_170 ^ cgp_core_169;
  assign cgp_core_173 = cgp_core_170 & cgp_core_169;
  assign cgp_core_174 = cgp_core_171 | cgp_core_173;
  assign cgp_core_175 = cgp_core_098 ^ cgp_core_157;
  assign cgp_core_176 = cgp_core_098 & cgp_core_157;
  assign cgp_core_177 = cgp_core_175 ^ cgp_core_174;
  assign cgp_core_178 = cgp_core_175 & cgp_core_174;
  assign cgp_core_179 = cgp_core_176 | cgp_core_178;
  assign cgp_core_181 = ~input_a[25];
  assign cgp_core_183 = ~(input_a[37] | input_a[16]);
  assign cgp_core_185 = input_a[43] | input_a[1];
  assign cgp_core_186 = input_a[22] & input_a[4];
  assign cgp_core_187 = ~(input_a[13] | input_a[32]);
  assign cgp_core_188 = ~input_a[32];
  assign cgp_core_189 = input_a[26] | input_a[7];
  assign cgp_core_191 = ~(input_a[29] | input_a[31]);
  assign cgp_core_194 = input_a[5] & input_a[33];
  assign cgp_core_197 = cgp_core_186 | cgp_core_194;
  assign cgp_core_198 = ~input_a[16];
  assign cgp_core_199 = ~(input_a[12] ^ input_a[4]);
  assign cgp_core_201 = input_a[4] & input_a[40];
  assign cgp_core_202 = ~input_a[30];
  assign cgp_core_203 = ~input_a[10];
  assign cgp_core_204 = ~(input_a[20] | input_a[23]);
  assign cgp_core_205 = ~input_a[4];
  assign cgp_core_207 = input_a[18] ^ input_a[1];
  assign cgp_core_208 = input_a[31] ^ input_a[32];
  assign cgp_core_209 = input_a[31] & input_a[32];
  assign cgp_core_210 = input_a[30] ^ cgp_core_208;
  assign cgp_core_211 = input_a[30] & cgp_core_208;
  assign cgp_core_212 = cgp_core_209 | cgp_core_211;
  assign cgp_core_214 = input_a[41] ^ cgp_core_210;
  assign cgp_core_215 = input_a[41] & cgp_core_210;
  assign cgp_core_218 = cgp_core_212 ^ cgp_core_215;
  assign cgp_core_219 = cgp_core_212 & cgp_core_215;
  assign cgp_core_222 = ~(input_a[42] | input_a[24]);
  assign cgp_core_225 = ~(input_a[26] | input_a[32]);
  assign cgp_core_226 = input_a[9] ^ input_a[1];
  assign cgp_core_227 = input_a[17] & cgp_core_214;
  assign cgp_core_228 = cgp_core_197 ^ cgp_core_218;
  assign cgp_core_229 = cgp_core_197 & cgp_core_218;
  assign cgp_core_230 = cgp_core_228 ^ cgp_core_227;
  assign cgp_core_231 = cgp_core_228 & cgp_core_227;
  assign cgp_core_232 = cgp_core_229 | cgp_core_231;
  assign cgp_core_235 = cgp_core_219 | cgp_core_232;
  assign cgp_core_236 = ~(input_a[31] & input_a[14]);
  assign cgp_core_237 = ~(input_a[0] ^ input_a[27]);
  assign cgp_core_238 = ~input_a[13];
  assign cgp_core_239 = ~input_a[5];
  assign cgp_core_241 = input_a[31] | input_a[5];
  assign cgp_core_242 = ~(input_a[15] & input_a[18]);
  assign cgp_core_243 = ~(input_a[11] | input_a[19]);
  assign cgp_core_244 = ~(input_a[29] & input_a[36]);
  assign cgp_core_246 = ~(input_a[17] ^ input_a[12]);
  assign cgp_core_247 = ~(input_a[33] & input_a[6]);
  assign cgp_core_248 = ~input_a[3];
  assign cgp_core_250 = ~(input_a[0] ^ input_a[11]);
  assign cgp_core_252 = ~input_a[42];
  assign cgp_core_254 = ~(input_a[43] | input_a[42]);
  assign cgp_core_255 = ~(input_a[40] ^ input_a[22]);
  assign cgp_core_256 = input_a[16] & input_a[3];
  assign cgp_core_258 = ~(input_a[40] | input_a[40]);
  assign cgp_core_260 = input_a[44] ^ input_a[35];
  assign cgp_core_261 = ~input_a[38];
  assign cgp_core_262 = ~(input_a[33] ^ input_a[34]);
  assign cgp_core_263 = input_a[29] | input_a[9];
  assign cgp_core_266 = ~input_a[17];
  assign cgp_core_267 = ~(input_a[16] ^ input_a[25]);
  assign cgp_core_268 = input_a[41] | input_a[6];
  assign cgp_core_269 = input_a[22] ^ input_a[13];
  assign cgp_core_272 = input_a[33] | input_a[44];
  assign cgp_core_273 = input_a[12] ^ input_a[32];
  assign cgp_core_274 = input_a[6] | input_a[37];
  assign cgp_core_275 = ~(input_a[40] ^ input_a[40]);
  assign cgp_core_276 = ~(input_a[21] & input_a[39]);
  assign cgp_core_277 = ~input_a[6];
  assign cgp_core_278 = ~input_a[9];
  assign cgp_core_279 = ~(input_a[34] & input_a[38]);
  assign cgp_core_280 = input_a[35] & input_a[26];
  assign cgp_core_282 = input_a[30] | input_a[17];
  assign cgp_core_286 = input_a[24] & input_a[44];
  assign cgp_core_287 = input_a[43] | input_a[40];
  assign cgp_core_288 = ~(input_a[16] ^ input_a[5]);
  assign cgp_core_289 = ~(input_a[17] & input_a[41]);
  assign cgp_core_291 = ~(input_a[8] ^ input_a[20]);
  assign cgp_core_293 = cgp_core_256 ^ cgp_core_280;
  assign cgp_core_294 = cgp_core_256 & cgp_core_280;
  assign cgp_core_296 = ~input_a[27];
  assign cgp_core_301 = ~(input_a[20] | input_a[13]);
  assign cgp_core_303 = ~(input_a[4] | input_a[20]);
  assign cgp_core_304 = input_a[3] ^ input_a[20];
  assign cgp_core_306 = ~input_a[11];
  assign cgp_core_308 = ~(input_a[13] ^ input_a[25]);
  assign cgp_core_309 = input_a[37] | input_a[18];
  assign cgp_core_310 = cgp_core_230 ^ cgp_core_293;
  assign cgp_core_311 = cgp_core_230 & cgp_core_293;
  assign cgp_core_312 = cgp_core_310 ^ input_a[28];
  assign cgp_core_313 = cgp_core_310 & input_a[28];
  assign cgp_core_314 = cgp_core_311 | cgp_core_313;
  assign cgp_core_315 = cgp_core_235 ^ cgp_core_294;
  assign cgp_core_316 = cgp_core_235 & cgp_core_294;
  assign cgp_core_317 = cgp_core_315 ^ cgp_core_314;
  assign cgp_core_318 = cgp_core_315 & cgp_core_314;
  assign cgp_core_319 = cgp_core_316 | cgp_core_318;
  assign cgp_core_322 = ~cgp_core_319;
  assign cgp_core_328 = ~(input_a[16] | input_a[34]);
  assign cgp_core_329 = ~(input_a[4] | input_a[8]);
  assign cgp_core_330 = ~input_a[22];
  assign cgp_core_331 = input_a[38] & input_a[27];
  assign cgp_core_332 = cgp_core_167 ^ cgp_core_312;
  assign cgp_core_333 = cgp_core_167 & cgp_core_312;
  assign cgp_core_334 = cgp_core_332 ^ cgp_core_331;
  assign cgp_core_335 = cgp_core_332 & cgp_core_331;
  assign cgp_core_336 = cgp_core_333 | cgp_core_335;
  assign cgp_core_337 = cgp_core_172 ^ cgp_core_317;
  assign cgp_core_338 = cgp_core_172 & cgp_core_317;
  assign cgp_core_339 = cgp_core_337 ^ cgp_core_336;
  assign cgp_core_340 = cgp_core_337 & cgp_core_336;
  assign cgp_core_341 = cgp_core_338 | cgp_core_340;
  assign cgp_core_342 = cgp_core_177 ^ cgp_core_322;
  assign cgp_core_343 = cgp_core_177 & cgp_core_322;
  assign cgp_core_344 = cgp_core_342 ^ cgp_core_341;
  assign cgp_core_345 = cgp_core_342 & cgp_core_341;
  assign cgp_core_346 = cgp_core_343 | cgp_core_345;
  assign cgp_core_347 = cgp_core_179 ^ cgp_core_319;
  assign cgp_core_348 = cgp_core_179 & cgp_core_319;
  assign cgp_core_349 = cgp_core_347 ^ cgp_core_346;
  assign cgp_core_350 = cgp_core_347 & cgp_core_346;
  assign cgp_core_351 = cgp_core_348 | cgp_core_350;
  assign cgp_core_352 = input_a[24] & input_a[18];
  assign cgp_core_354 = ~(input_a[31] & input_a[18]);
  assign cgp_core_355 = ~(input_a[29] | input_a[35]);

  assign cgp_out[0] = input_a[23];
  assign cgp_out[1] = cgp_core_334;
  assign cgp_out[2] = cgp_core_339;
  assign cgp_out[3] = cgp_core_344;
  assign cgp_out[4] = cgp_core_349;
  assign cgp_out[5] = cgp_core_351;
endmodule

module cmp_neg(input [38:0] input_a, output [5:0] cgp_out);
  wire cgp_core_041;
  wire cgp_core_042;
  wire cgp_core_043;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_046;
  wire cgp_core_047;
  wire cgp_core_048;
  wire cgp_core_049;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_060;
  wire cgp_core_062;
  wire cgp_core_066;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_074;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_082;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_099;
  wire cgp_core_101;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_111;
  wire cgp_core_113;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_119;
  wire cgp_core_121;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_127;
  wire cgp_core_128;
  wire cgp_core_133;
  wire cgp_core_134;
  wire cgp_core_136;
  wire cgp_core_138;
  wire cgp_core_140;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_158;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_162;
  wire cgp_core_164;
  wire cgp_core_166;
  wire cgp_core_167;
  wire cgp_core_168;
  wire cgp_core_169;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_189;
  wire cgp_core_190;
  wire cgp_core_193;
  wire cgp_core_197;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_203;
  wire cgp_core_210;
  wire cgp_core_212;
  wire cgp_core_213;
  wire cgp_core_216;
  wire cgp_core_217;
  wire cgp_core_222;
  wire cgp_core_225;
  wire cgp_core_226;
  wire cgp_core_227;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_230;
  wire cgp_core_232;
  wire cgp_core_233;
  wire cgp_core_235;
  wire cgp_core_237;
  wire cgp_core_238;
  wire cgp_core_239;
  wire cgp_core_240;
  wire cgp_core_243;
  wire cgp_core_244;
  wire cgp_core_246;
  wire cgp_core_247;
  wire cgp_core_252;
  wire cgp_core_255;
  wire cgp_core_256;
  wire cgp_core_258;
  wire cgp_core_259;
  wire cgp_core_262;
  wire cgp_core_265;
  wire cgp_core_267;
  wire cgp_core_268;
  wire cgp_core_271;
  wire cgp_core_272;
  wire cgp_core_276;
  wire cgp_core_278;
  wire cgp_core_279;
  wire cgp_core_280;
  wire cgp_core_282;
  wire cgp_core_283;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_290;
  wire cgp_core_291;
  wire cgp_core_292;
  wire cgp_core_293;
  wire cgp_core_294;
  wire cgp_core_295;
  wire cgp_core_296;
  wire cgp_core_298;
  wire cgp_core_299;
  wire cgp_core_302;
  wire cgp_core_303;
  wire cgp_core_305;
  wire cgp_core_306;

  assign cgp_core_041 = input_a[0] ^ input_a[1];
  assign cgp_core_042 = input_a[0] & input_a[1];
  assign cgp_core_043 = ~(input_a[2] & input_a[3]);
  assign cgp_core_044 = input_a[2] & input_a[3];
  assign cgp_core_045 = ~(input_a[23] ^ input_a[1]);
  assign cgp_core_046 = input_a[37] & cgp_core_043;
  assign cgp_core_047 = cgp_core_042 ^ cgp_core_044;
  assign cgp_core_048 = cgp_core_042 & cgp_core_044;
  assign cgp_core_049 = cgp_core_047 | cgp_core_046;
  assign cgp_core_052 = ~(input_a[22] | input_a[35]);
  assign cgp_core_053 = ~(input_a[19] ^ input_a[3]);
  assign cgp_core_055 = ~(input_a[16] & input_a[7]);
  assign cgp_core_057 = input_a[7] ^ input_a[16];
  assign cgp_core_060 = ~input_a[30];
  assign cgp_core_062 = input_a[16] | input_a[30];
  assign cgp_core_066 = ~input_a[2];
  assign cgp_core_068 = input_a[26] ^ input_a[31];
  assign cgp_core_069 = ~(input_a[22] ^ input_a[3]);
  assign cgp_core_071 = cgp_core_049 ^ cgp_core_062;
  assign cgp_core_072 = cgp_core_049 & cgp_core_062;
  assign cgp_core_074 = input_a[21] & input_a[10];
  assign cgp_core_077 = ~(input_a[15] | input_a[20]);
  assign cgp_core_078 = cgp_core_048 | cgp_core_072;
  assign cgp_core_079 = ~input_a[8];
  assign cgp_core_080 = ~(input_a[28] & input_a[32]);
  assign cgp_core_082 = input_a[20] ^ input_a[38];
  assign cgp_core_084 = input_a[5] & input_a[4];
  assign cgp_core_085 = input_a[12] ^ input_a[13];
  assign cgp_core_086 = input_a[12] & input_a[13];
  assign cgp_core_087 = ~(input_a[38] | input_a[36]);
  assign cgp_core_088 = input_a[11] & cgp_core_085;
  assign cgp_core_089 = cgp_core_086 | cgp_core_088;
  assign cgp_core_092 = input_a[32] & input_a[23];
  assign cgp_core_093 = cgp_core_084 ^ cgp_core_089;
  assign cgp_core_094 = cgp_core_084 & cgp_core_089;
  assign cgp_core_095 = cgp_core_093 ^ cgp_core_092;
  assign cgp_core_096 = cgp_core_093 & cgp_core_092;
  assign cgp_core_097 = cgp_core_094 | cgp_core_096;
  assign cgp_core_099 = ~input_a[35];
  assign cgp_core_101 = input_a[20] & input_a[15];
  assign cgp_core_102 = input_a[17] ^ input_a[18];
  assign cgp_core_103 = input_a[17] & input_a[18];
  assign cgp_core_104 = ~(input_a[31] | input_a[15]);
  assign cgp_core_105 = input_a[33] & cgp_core_102;
  assign cgp_core_106 = cgp_core_103 | cgp_core_105;
  assign cgp_core_109 = input_a[4] ^ input_a[34];
  assign cgp_core_110 = cgp_core_101 ^ cgp_core_106;
  assign cgp_core_111 = cgp_core_101 & cgp_core_106;
  assign cgp_core_113 = ~(input_a[4] & input_a[12]);
  assign cgp_core_116 = input_a[19] & input_a[8];
  assign cgp_core_117 = ~input_a[4];
  assign cgp_core_119 = cgp_core_095 ^ cgp_core_110;
  assign cgp_core_121 = ~cgp_core_119;
  assign cgp_core_123 = cgp_core_095 | cgp_core_119;
  assign cgp_core_124 = cgp_core_097 ^ cgp_core_111;
  assign cgp_core_125 = cgp_core_097 & cgp_core_111;
  assign cgp_core_126 = cgp_core_124 ^ cgp_core_123;
  assign cgp_core_127 = cgp_core_124 & cgp_core_123;
  assign cgp_core_128 = cgp_core_125 | cgp_core_127;
  assign cgp_core_133 = ~input_a[5];
  assign cgp_core_134 = ~input_a[5];
  assign cgp_core_136 = cgp_core_071 ^ cgp_core_121;
  assign cgp_core_138 = ~cgp_core_136;
  assign cgp_core_140 = cgp_core_071 | cgp_core_136;
  assign cgp_core_141 = cgp_core_078 ^ cgp_core_126;
  assign cgp_core_142 = cgp_core_078 & cgp_core_126;
  assign cgp_core_143 = cgp_core_141 ^ cgp_core_140;
  assign cgp_core_144 = cgp_core_141 & cgp_core_140;
  assign cgp_core_145 = cgp_core_142 | cgp_core_144;
  assign cgp_core_148 = cgp_core_128 ^ cgp_core_145;
  assign cgp_core_149 = cgp_core_128 & cgp_core_145;
  assign cgp_core_154 = ~(input_a[9] | input_a[25]);
  assign cgp_core_155 = input_a[5] ^ input_a[10];
  assign cgp_core_156 = input_a[19] ^ input_a[36];
  assign cgp_core_157 = input_a[19] & input_a[8];
  assign cgp_core_158 = input_a[17] ^ input_a[10];
  assign cgp_core_159 = input_a[31] & input_a[9];
  assign cgp_core_160 = ~(input_a[2] | input_a[38]);
  assign cgp_core_162 = cgp_core_159 | input_a[35];
  assign cgp_core_164 = ~input_a[7];
  assign cgp_core_166 = cgp_core_157 ^ cgp_core_162;
  assign cgp_core_167 = cgp_core_157 & input_a[35];
  assign cgp_core_168 = cgp_core_166 ^ input_a[14];
  assign cgp_core_169 = cgp_core_166 & input_a[14];
  assign cgp_core_170 = cgp_core_167 | cgp_core_169;
  assign cgp_core_171 = cgp_core_159 | cgp_core_170;
  assign cgp_core_172 = input_a[30] ^ input_a[34];
  assign cgp_core_173 = input_a[24] ^ input_a[25];
  assign cgp_core_174 = input_a[24] & input_a[25];
  assign cgp_core_175 = input_a[27] ^ input_a[28];
  assign cgp_core_176 = input_a[27] & input_a[28];
  assign cgp_core_177 = input_a[26] ^ cgp_core_175;
  assign cgp_core_178 = input_a[26] & cgp_core_175;
  assign cgp_core_179 = cgp_core_176 | cgp_core_178;
  assign cgp_core_182 = cgp_core_173 & cgp_core_177;
  assign cgp_core_183 = cgp_core_174 ^ cgp_core_179;
  assign cgp_core_184 = cgp_core_174 & cgp_core_179;
  assign cgp_core_185 = cgp_core_183 ^ cgp_core_182;
  assign cgp_core_186 = cgp_core_183 & cgp_core_182;
  assign cgp_core_187 = cgp_core_184 | cgp_core_186;
  assign cgp_core_189 = input_a[10] | input_a[1];
  assign cgp_core_190 = input_a[13] ^ input_a[3];
  assign cgp_core_193 = cgp_core_168 & cgp_core_185;
  assign cgp_core_197 = cgp_core_171 ^ cgp_core_187;
  assign cgp_core_199 = cgp_core_197 | cgp_core_193;
  assign cgp_core_200 = input_a[34] & cgp_core_193;
  assign cgp_core_201 = cgp_core_171 | cgp_core_200;
  assign cgp_core_203 = ~input_a[34];
  assign cgp_core_210 = ~(input_a[4] ^ input_a[35]);
  assign cgp_core_212 = input_a[36] | input_a[20];
  assign cgp_core_213 = input_a[38] ^ input_a[37];
  assign cgp_core_216 = ~(input_a[2] ^ input_a[0]);
  assign cgp_core_217 = input_a[18] ^ input_a[18];
  assign cgp_core_222 = input_a[3] | input_a[6];
  assign cgp_core_225 = input_a[38] & input_a[22];
  assign cgp_core_226 = ~(input_a[1] & input_a[36]);
  assign cgp_core_227 = ~(input_a[33] ^ input_a[4]);
  assign cgp_core_228 = input_a[34] ^ input_a[14];
  assign cgp_core_229 = input_a[37] | input_a[13];
  assign cgp_core_230 = ~(input_a[16] | input_a[31]);
  assign cgp_core_232 = ~(input_a[33] | input_a[12]);
  assign cgp_core_233 = input_a[4] | input_a[21];
  assign cgp_core_235 = ~input_a[15];
  assign cgp_core_237 = ~(input_a[19] & input_a[19]);
  assign cgp_core_238 = input_a[33] ^ input_a[38];
  assign cgp_core_239 = ~input_a[38];
  assign cgp_core_240 = ~(input_a[12] ^ input_a[3]);
  assign cgp_core_243 = ~cgp_core_225;
  assign cgp_core_244 = input_a[4] & cgp_core_225;
  assign cgp_core_246 = ~cgp_core_243;
  assign cgp_core_247 = cgp_core_244 | cgp_core_246;
  assign cgp_core_252 = input_a[37] ^ input_a[21];
  assign cgp_core_255 = ~(input_a[30] & input_a[7]);
  assign cgp_core_256 = ~(input_a[5] ^ input_a[7]);
  assign cgp_core_258 = input_a[20] & input_a[22];
  assign cgp_core_259 = input_a[8] & input_a[10];
  assign cgp_core_262 = ~cgp_core_243;
  assign cgp_core_265 = cgp_core_199 ^ cgp_core_247;
  assign cgp_core_267 = cgp_core_265 ^ cgp_core_243;
  assign cgp_core_268 = input_a[20] & input_a[14];
  assign cgp_core_271 = ~(input_a[0] | input_a[37]);
  assign cgp_core_272 = cgp_core_201 | cgp_core_199;
  assign cgp_core_276 = input_a[15] & input_a[6];
  assign cgp_core_278 = ~(input_a[22] ^ input_a[17]);
  assign cgp_core_279 = ~input_a[0];
  assign cgp_core_280 = input_a[27] & input_a[18];
  assign cgp_core_282 = cgp_core_138 ^ cgp_core_262;
  assign cgp_core_283 = cgp_core_138 & cgp_core_262;
  assign cgp_core_287 = cgp_core_143 ^ cgp_core_267;
  assign cgp_core_288 = cgp_core_143 & cgp_core_267;
  assign cgp_core_289 = cgp_core_287 ^ cgp_core_283;
  assign cgp_core_290 = cgp_core_287 & cgp_core_283;
  assign cgp_core_291 = cgp_core_288 | cgp_core_290;
  assign cgp_core_292 = cgp_core_148 ^ cgp_core_272;
  assign cgp_core_293 = cgp_core_148 & cgp_core_272;
  assign cgp_core_294 = cgp_core_292 ^ cgp_core_291;
  assign cgp_core_295 = cgp_core_292 & cgp_core_291;
  assign cgp_core_296 = cgp_core_293 | cgp_core_295;
  assign cgp_core_298 = input_a[10] & input_a[27];
  assign cgp_core_299 = cgp_core_149 ^ cgp_core_296;
  assign cgp_core_302 = ~(input_a[35] ^ input_a[1]);
  assign cgp_core_303 = ~(input_a[30] ^ input_a[35]);
  assign cgp_core_305 = input_a[30] & input_a[15];
  assign cgp_core_306 = input_a[23] ^ input_a[17];

  assign cgp_out[0] = input_a[34];
  assign cgp_out[1] = cgp_core_282;
  assign cgp_out[2] = cgp_core_289;
  assign cgp_out[3] = cgp_core_294;
  assign cgp_out[4] = cgp_core_299;
  assign cgp_out[5] = 1'b0;
endmodule
module pcc(input [44:0] pos, input [38:0] neg, output outval);
    wire [5:0] cnt_pos;
    wire [5:0] cnt_neg;

    cmp_pos ipos(pos, cnt_pos);
    cmp_neg ineg(neg, cnt_neg);

    assign outval = (cnt_pos >= cnt_neg);
endmodule
