// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.09375
// WCE=4.0
// EP=0.726562%
// Printed PDK parameters:
//  Area=34250257.0
//  Delay=62472784.0
//  Power=1710900.0

module popcount19_vq19(input [18:0] input_a, output [4:0] popcount19_vq19_out);
  wire popcount19_vq19_core_021;
  wire popcount19_vq19_core_022;
  wire popcount19_vq19_core_023;
  wire popcount19_vq19_core_024;
  wire popcount19_vq19_core_026;
  wire popcount19_vq19_core_027;
  wire popcount19_vq19_core_028;
  wire popcount19_vq19_core_029;
  wire popcount19_vq19_core_030;
  wire popcount19_vq19_core_031;
  wire popcount19_vq19_core_032;
  wire popcount19_vq19_core_033;
  wire popcount19_vq19_core_034;
  wire popcount19_vq19_core_035;
  wire popcount19_vq19_core_036;
  wire popcount19_vq19_core_037;
  wire popcount19_vq19_core_038;
  wire popcount19_vq19_core_042;
  wire popcount19_vq19_core_043;
  wire popcount19_vq19_core_044;
  wire popcount19_vq19_core_045;
  wire popcount19_vq19_core_046_not;
  wire popcount19_vq19_core_047;
  wire popcount19_vq19_core_048;
  wire popcount19_vq19_core_049;
  wire popcount19_vq19_core_050;
  wire popcount19_vq19_core_051;
  wire popcount19_vq19_core_052;
  wire popcount19_vq19_core_057;
  wire popcount19_vq19_core_058;
  wire popcount19_vq19_core_060;
  wire popcount19_vq19_core_062;
  wire popcount19_vq19_core_063_not;
  wire popcount19_vq19_core_064;
  wire popcount19_vq19_core_065;
  wire popcount19_vq19_core_067;
  wire popcount19_vq19_core_068;
  wire popcount19_vq19_core_069;
  wire popcount19_vq19_core_071;
  wire popcount19_vq19_core_072;
  wire popcount19_vq19_core_073;
  wire popcount19_vq19_core_074;
  wire popcount19_vq19_core_075;
  wire popcount19_vq19_core_076;
  wire popcount19_vq19_core_077;
  wire popcount19_vq19_core_079;
  wire popcount19_vq19_core_080;
  wire popcount19_vq19_core_081;
  wire popcount19_vq19_core_082;
  wire popcount19_vq19_core_083;
  wire popcount19_vq19_core_084;
  wire popcount19_vq19_core_085;
  wire popcount19_vq19_core_086;
  wire popcount19_vq19_core_089;
  wire popcount19_vq19_core_090;
  wire popcount19_vq19_core_091;
  wire popcount19_vq19_core_092;
  wire popcount19_vq19_core_093;
  wire popcount19_vq19_core_094;
  wire popcount19_vq19_core_096;
  wire popcount19_vq19_core_097;
  wire popcount19_vq19_core_099;
  wire popcount19_vq19_core_100;
  wire popcount19_vq19_core_101;
  wire popcount19_vq19_core_102;
  wire popcount19_vq19_core_103;
  wire popcount19_vq19_core_104;
  wire popcount19_vq19_core_105;
  wire popcount19_vq19_core_106;
  wire popcount19_vq19_core_107;
  wire popcount19_vq19_core_108;
  wire popcount19_vq19_core_113;
  wire popcount19_vq19_core_115;
  wire popcount19_vq19_core_116;
  wire popcount19_vq19_core_117;
  wire popcount19_vq19_core_118;
  wire popcount19_vq19_core_119;
  wire popcount19_vq19_core_121;
  wire popcount19_vq19_core_122;
  wire popcount19_vq19_core_123;
  wire popcount19_vq19_core_124;
  wire popcount19_vq19_core_125;
  wire popcount19_vq19_core_127;
  wire popcount19_vq19_core_128;
  wire popcount19_vq19_core_129;
  wire popcount19_vq19_core_130;
  wire popcount19_vq19_core_131;
  wire popcount19_vq19_core_133;
  wire popcount19_vq19_core_134;
  wire popcount19_vq19_core_135;

  assign popcount19_vq19_core_021 = input_a[0] ^ input_a[1];
  assign popcount19_vq19_core_022 = input_a[0] & input_a[1];
  assign popcount19_vq19_core_023 = input_a[4] | input_a[4];
  assign popcount19_vq19_core_024 = input_a[8] & input_a[7];
  assign popcount19_vq19_core_026 = popcount19_vq19_core_021 & input_a[3];
  assign popcount19_vq19_core_027 = popcount19_vq19_core_022 ^ popcount19_vq19_core_024;
  assign popcount19_vq19_core_028 = popcount19_vq19_core_022 & popcount19_vq19_core_024;
  assign popcount19_vq19_core_029 = popcount19_vq19_core_027 ^ popcount19_vq19_core_026;
  assign popcount19_vq19_core_030 = popcount19_vq19_core_027 & popcount19_vq19_core_026;
  assign popcount19_vq19_core_031 = popcount19_vq19_core_028 | popcount19_vq19_core_030;
  assign popcount19_vq19_core_032 = input_a[7] | input_a[10];
  assign popcount19_vq19_core_033 = ~(input_a[13] ^ input_a[18]);
  assign popcount19_vq19_core_034 = ~(input_a[14] | input_a[10]);
  assign popcount19_vq19_core_035 = ~(input_a[14] & input_a[16]);
  assign popcount19_vq19_core_036 = input_a[14] | input_a[14];
  assign popcount19_vq19_core_037 = input_a[11] | input_a[12];
  assign popcount19_vq19_core_038 = ~input_a[5];
  assign popcount19_vq19_core_042 = input_a[11] ^ input_a[15];
  assign popcount19_vq19_core_043 = ~input_a[0];
  assign popcount19_vq19_core_044 = input_a[4] | input_a[5];
  assign popcount19_vq19_core_045 = ~input_a[7];
  assign popcount19_vq19_core_046_not = ~input_a[15];
  assign popcount19_vq19_core_047 = input_a[6] | input_a[4];
  assign popcount19_vq19_core_048 = ~(input_a[12] & input_a[4]);
  assign popcount19_vq19_core_049 = input_a[4] ^ input_a[3];
  assign popcount19_vq19_core_050 = ~(input_a[8] ^ input_a[5]);
  assign popcount19_vq19_core_051 = popcount19_vq19_core_029 ^ popcount19_vq19_core_044;
  assign popcount19_vq19_core_052 = popcount19_vq19_core_029 & popcount19_vq19_core_044;
  assign popcount19_vq19_core_057 = input_a[12] | input_a[8];
  assign popcount19_vq19_core_058 = popcount19_vq19_core_031 | popcount19_vq19_core_052;
  assign popcount19_vq19_core_060 = input_a[1] & input_a[0];
  assign popcount19_vq19_core_062 = ~(input_a[18] | input_a[0]);
  assign popcount19_vq19_core_063_not = ~input_a[2];
  assign popcount19_vq19_core_064 = input_a[9] & input_a[10];
  assign popcount19_vq19_core_065 = input_a[18] ^ input_a[18];
  assign popcount19_vq19_core_067 = ~input_a[2];
  assign popcount19_vq19_core_068 = input_a[0] & input_a[2];
  assign popcount19_vq19_core_069 = input_a[12] | input_a[11];
  assign popcount19_vq19_core_071 = ~input_a[12];
  assign popcount19_vq19_core_072 = input_a[6] & popcount19_vq19_core_067;
  assign popcount19_vq19_core_073 = popcount19_vq19_core_064 ^ popcount19_vq19_core_069;
  assign popcount19_vq19_core_074 = popcount19_vq19_core_064 & popcount19_vq19_core_069;
  assign popcount19_vq19_core_075 = popcount19_vq19_core_073 ^ popcount19_vq19_core_072;
  assign popcount19_vq19_core_076 = popcount19_vq19_core_073 & popcount19_vq19_core_072;
  assign popcount19_vq19_core_077 = popcount19_vq19_core_074 | popcount19_vq19_core_076;
  assign popcount19_vq19_core_079 = input_a[7] ^ input_a[9];
  assign popcount19_vq19_core_080 = input_a[10] | input_a[16];
  assign popcount19_vq19_core_081 = input_a[14] & input_a[15];
  assign popcount19_vq19_core_082 = input_a[17] ^ input_a[18];
  assign popcount19_vq19_core_083 = input_a[17] & input_a[18];
  assign popcount19_vq19_core_084 = input_a[16] ^ popcount19_vq19_core_082;
  assign popcount19_vq19_core_085 = input_a[16] & popcount19_vq19_core_082;
  assign popcount19_vq19_core_086 = popcount19_vq19_core_083 | popcount19_vq19_core_085;
  assign popcount19_vq19_core_089 = input_a[13] & popcount19_vq19_core_084;
  assign popcount19_vq19_core_090 = popcount19_vq19_core_081 ^ popcount19_vq19_core_086;
  assign popcount19_vq19_core_091 = popcount19_vq19_core_081 & popcount19_vq19_core_086;
  assign popcount19_vq19_core_092 = popcount19_vq19_core_090 ^ popcount19_vq19_core_089;
  assign popcount19_vq19_core_093 = popcount19_vq19_core_090 & popcount19_vq19_core_089;
  assign popcount19_vq19_core_094 = popcount19_vq19_core_091 | popcount19_vq19_core_093;
  assign popcount19_vq19_core_096 = input_a[4] ^ input_a[13];
  assign popcount19_vq19_core_097 = ~(input_a[17] ^ input_a[0]);
  assign popcount19_vq19_core_099 = popcount19_vq19_core_075 ^ popcount19_vq19_core_092;
  assign popcount19_vq19_core_100 = popcount19_vq19_core_075 & popcount19_vq19_core_092;
  assign popcount19_vq19_core_101 = popcount19_vq19_core_099 ^ input_a[2];
  assign popcount19_vq19_core_102 = popcount19_vq19_core_099 & input_a[2];
  assign popcount19_vq19_core_103 = popcount19_vq19_core_100 | popcount19_vq19_core_102;
  assign popcount19_vq19_core_104 = popcount19_vq19_core_077 ^ popcount19_vq19_core_094;
  assign popcount19_vq19_core_105 = popcount19_vq19_core_077 & popcount19_vq19_core_094;
  assign popcount19_vq19_core_106 = popcount19_vq19_core_104 ^ popcount19_vq19_core_103;
  assign popcount19_vq19_core_107 = popcount19_vq19_core_104 & popcount19_vq19_core_103;
  assign popcount19_vq19_core_108 = popcount19_vq19_core_105 | popcount19_vq19_core_107;
  assign popcount19_vq19_core_113 = ~(input_a[18] & input_a[1]);
  assign popcount19_vq19_core_115 = input_a[8] | input_a[0];
  assign popcount19_vq19_core_116 = popcount19_vq19_core_051 ^ popcount19_vq19_core_101;
  assign popcount19_vq19_core_117 = popcount19_vq19_core_051 & popcount19_vq19_core_101;
  assign popcount19_vq19_core_118 = ~(input_a[17] ^ input_a[8]);
  assign popcount19_vq19_core_119 = input_a[13] & input_a[12];
  assign popcount19_vq19_core_121 = popcount19_vq19_core_058 ^ popcount19_vq19_core_106;
  assign popcount19_vq19_core_122 = popcount19_vq19_core_058 & popcount19_vq19_core_106;
  assign popcount19_vq19_core_123 = popcount19_vq19_core_121 ^ popcount19_vq19_core_117;
  assign popcount19_vq19_core_124 = popcount19_vq19_core_121 & popcount19_vq19_core_117;
  assign popcount19_vq19_core_125 = popcount19_vq19_core_122 | popcount19_vq19_core_124;
  assign popcount19_vq19_core_127 = input_a[16] ^ input_a[12];
  assign popcount19_vq19_core_128 = popcount19_vq19_core_108 ^ popcount19_vq19_core_125;
  assign popcount19_vq19_core_129 = popcount19_vq19_core_108 & popcount19_vq19_core_125;
  assign popcount19_vq19_core_130 = input_a[8] ^ input_a[14];
  assign popcount19_vq19_core_131 = ~input_a[8];
  assign popcount19_vq19_core_133 = ~(input_a[16] | input_a[11]);
  assign popcount19_vq19_core_134 = ~(input_a[18] | input_a[6]);
  assign popcount19_vq19_core_135 = ~(input_a[9] | input_a[6]);

  assign popcount19_vq19_out[0] = 1'b1;
  assign popcount19_vq19_out[1] = popcount19_vq19_core_116;
  assign popcount19_vq19_out[2] = popcount19_vq19_core_123;
  assign popcount19_vq19_out[3] = popcount19_vq19_core_128;
  assign popcount19_vq19_out[4] = popcount19_vq19_core_129;
endmodule