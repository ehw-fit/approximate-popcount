// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=15.5666
// WCE=43.0
// EP=0.985557%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount32_k31q(input [31:0] input_a, output [5:0] popcount32_k31q_out);
  wire popcount32_k31q_core_036;
  wire popcount32_k31q_core_039;
  wire popcount32_k31q_core_041;
  wire popcount32_k31q_core_042;
  wire popcount32_k31q_core_044;
  wire popcount32_k31q_core_046;
  wire popcount32_k31q_core_051;
  wire popcount32_k31q_core_053;
  wire popcount32_k31q_core_056;
  wire popcount32_k31q_core_057_not;
  wire popcount32_k31q_core_058;
  wire popcount32_k31q_core_059;
  wire popcount32_k31q_core_063;
  wire popcount32_k31q_core_066;
  wire popcount32_k31q_core_067;
  wire popcount32_k31q_core_070;
  wire popcount32_k31q_core_071;
  wire popcount32_k31q_core_075;
  wire popcount32_k31q_core_078;
  wire popcount32_k31q_core_079;
  wire popcount32_k31q_core_080;
  wire popcount32_k31q_core_081_not;
  wire popcount32_k31q_core_083;
  wire popcount32_k31q_core_084;
  wire popcount32_k31q_core_085;
  wire popcount32_k31q_core_089;
  wire popcount32_k31q_core_091;
  wire popcount32_k31q_core_092;
  wire popcount32_k31q_core_094_not;
  wire popcount32_k31q_core_095;
  wire popcount32_k31q_core_096;
  wire popcount32_k31q_core_097;
  wire popcount32_k31q_core_099;
  wire popcount32_k31q_core_101;
  wire popcount32_k31q_core_102;
  wire popcount32_k31q_core_103;
  wire popcount32_k31q_core_104;
  wire popcount32_k31q_core_105;
  wire popcount32_k31q_core_106;
  wire popcount32_k31q_core_109;
  wire popcount32_k31q_core_110;
  wire popcount32_k31q_core_111;
  wire popcount32_k31q_core_112;
  wire popcount32_k31q_core_113;
  wire popcount32_k31q_core_116;
  wire popcount32_k31q_core_117_not;
  wire popcount32_k31q_core_118;
  wire popcount32_k31q_core_119;
  wire popcount32_k31q_core_120;
  wire popcount32_k31q_core_121;
  wire popcount32_k31q_core_123;
  wire popcount32_k31q_core_124;
  wire popcount32_k31q_core_126;
  wire popcount32_k31q_core_130;
  wire popcount32_k31q_core_131;
  wire popcount32_k31q_core_132;
  wire popcount32_k31q_core_134;
  wire popcount32_k31q_core_135;
  wire popcount32_k31q_core_136;
  wire popcount32_k31q_core_140;
  wire popcount32_k31q_core_142;
  wire popcount32_k31q_core_144;
  wire popcount32_k31q_core_145;
  wire popcount32_k31q_core_147;
  wire popcount32_k31q_core_148;
  wire popcount32_k31q_core_156;
  wire popcount32_k31q_core_158;
  wire popcount32_k31q_core_159;
  wire popcount32_k31q_core_160;
  wire popcount32_k31q_core_161;
  wire popcount32_k31q_core_162;
  wire popcount32_k31q_core_163;
  wire popcount32_k31q_core_166;
  wire popcount32_k31q_core_167;
  wire popcount32_k31q_core_168;
  wire popcount32_k31q_core_169;
  wire popcount32_k31q_core_170;
  wire popcount32_k31q_core_171;
  wire popcount32_k31q_core_176;
  wire popcount32_k31q_core_177;
  wire popcount32_k31q_core_178;
  wire popcount32_k31q_core_179_not;
  wire popcount32_k31q_core_180;
  wire popcount32_k31q_core_182;
  wire popcount32_k31q_core_184;
  wire popcount32_k31q_core_185;
  wire popcount32_k31q_core_186;
  wire popcount32_k31q_core_187;
  wire popcount32_k31q_core_188;
  wire popcount32_k31q_core_189;
  wire popcount32_k31q_core_190;
  wire popcount32_k31q_core_194;
  wire popcount32_k31q_core_195;
  wire popcount32_k31q_core_196;
  wire popcount32_k31q_core_197;
  wire popcount32_k31q_core_198;
  wire popcount32_k31q_core_199;
  wire popcount32_k31q_core_200;
  wire popcount32_k31q_core_201;
  wire popcount32_k31q_core_202;
  wire popcount32_k31q_core_204;
  wire popcount32_k31q_core_206;
  wire popcount32_k31q_core_208;
  wire popcount32_k31q_core_209;
  wire popcount32_k31q_core_211;
  wire popcount32_k31q_core_212;
  wire popcount32_k31q_core_213;
  wire popcount32_k31q_core_215;
  wire popcount32_k31q_core_216;
  wire popcount32_k31q_core_218;
  wire popcount32_k31q_core_219;
  wire popcount32_k31q_core_220;
  wire popcount32_k31q_core_223;
  wire popcount32_k31q_core_224;
  wire popcount32_k31q_core_225;

  assign popcount32_k31q_core_036 = ~(input_a[27] & input_a[2]);
  assign popcount32_k31q_core_039 = ~(input_a[16] & input_a[28]);
  assign popcount32_k31q_core_041 = ~(input_a[11] ^ input_a[30]);
  assign popcount32_k31q_core_042 = input_a[13] & input_a[26];
  assign popcount32_k31q_core_044 = input_a[11] ^ input_a[14];
  assign popcount32_k31q_core_046 = input_a[7] ^ input_a[9];
  assign popcount32_k31q_core_051 = input_a[5] | input_a[9];
  assign popcount32_k31q_core_053 = ~(input_a[15] & input_a[20]);
  assign popcount32_k31q_core_056 = input_a[30] | input_a[13];
  assign popcount32_k31q_core_057_not = ~input_a[7];
  assign popcount32_k31q_core_058 = input_a[19] ^ input_a[15];
  assign popcount32_k31q_core_059 = ~(input_a[18] ^ input_a[1]);
  assign popcount32_k31q_core_063 = ~input_a[20];
  assign popcount32_k31q_core_066 = ~(input_a[0] | input_a[24]);
  assign popcount32_k31q_core_067 = ~(input_a[29] & input_a[21]);
  assign popcount32_k31q_core_070 = ~(input_a[31] ^ input_a[4]);
  assign popcount32_k31q_core_071 = input_a[3] ^ input_a[21];
  assign popcount32_k31q_core_075 = ~(input_a[7] | input_a[14]);
  assign popcount32_k31q_core_078 = ~(input_a[8] | input_a[24]);
  assign popcount32_k31q_core_079 = ~(input_a[1] | input_a[4]);
  assign popcount32_k31q_core_080 = ~(input_a[15] ^ input_a[14]);
  assign popcount32_k31q_core_081_not = ~input_a[7];
  assign popcount32_k31q_core_083 = ~(input_a[16] | input_a[19]);
  assign popcount32_k31q_core_084 = ~(input_a[29] | input_a[1]);
  assign popcount32_k31q_core_085 = input_a[18] & input_a[11];
  assign popcount32_k31q_core_089 = input_a[24] ^ input_a[13];
  assign popcount32_k31q_core_091 = ~(input_a[22] | input_a[23]);
  assign popcount32_k31q_core_092 = ~(input_a[20] | input_a[12]);
  assign popcount32_k31q_core_094_not = ~input_a[10];
  assign popcount32_k31q_core_095 = input_a[5] ^ input_a[2];
  assign popcount32_k31q_core_096 = input_a[1] | input_a[13];
  assign popcount32_k31q_core_097 = input_a[4] ^ input_a[21];
  assign popcount32_k31q_core_099 = ~(input_a[12] | input_a[8]);
  assign popcount32_k31q_core_101 = ~(input_a[3] & input_a[28]);
  assign popcount32_k31q_core_102 = input_a[15] | input_a[29];
  assign popcount32_k31q_core_103 = ~(input_a[14] ^ input_a[12]);
  assign popcount32_k31q_core_104 = input_a[3] & input_a[6];
  assign popcount32_k31q_core_105 = ~(input_a[4] & input_a[23]);
  assign popcount32_k31q_core_106 = ~(input_a[1] ^ input_a[28]);
  assign popcount32_k31q_core_109 = ~input_a[12];
  assign popcount32_k31q_core_110 = input_a[7] | input_a[5];
  assign popcount32_k31q_core_111 = input_a[4] ^ input_a[16];
  assign popcount32_k31q_core_112 = ~(input_a[29] ^ input_a[23]);
  assign popcount32_k31q_core_113 = ~(input_a[24] & input_a[18]);
  assign popcount32_k31q_core_116 = input_a[23] & input_a[20];
  assign popcount32_k31q_core_117_not = ~input_a[4];
  assign popcount32_k31q_core_118 = ~input_a[6];
  assign popcount32_k31q_core_119 = input_a[18] | input_a[15];
  assign popcount32_k31q_core_120 = input_a[29] | input_a[22];
  assign popcount32_k31q_core_121 = ~(input_a[9] ^ input_a[0]);
  assign popcount32_k31q_core_123 = ~(input_a[17] & input_a[23]);
  assign popcount32_k31q_core_124 = ~(input_a[23] | input_a[17]);
  assign popcount32_k31q_core_126 = ~(input_a[20] ^ input_a[8]);
  assign popcount32_k31q_core_130 = ~(input_a[22] ^ input_a[28]);
  assign popcount32_k31q_core_131 = input_a[4] & input_a[31];
  assign popcount32_k31q_core_132 = input_a[15] & input_a[24];
  assign popcount32_k31q_core_134 = ~input_a[10];
  assign popcount32_k31q_core_135 = input_a[7] & input_a[8];
  assign popcount32_k31q_core_136 = input_a[4] | input_a[22];
  assign popcount32_k31q_core_140 = input_a[25] ^ input_a[22];
  assign popcount32_k31q_core_142 = input_a[8] ^ input_a[11];
  assign popcount32_k31q_core_144 = ~(input_a[15] & input_a[11]);
  assign popcount32_k31q_core_145 = ~(input_a[5] & input_a[12]);
  assign popcount32_k31q_core_147 = ~input_a[6];
  assign popcount32_k31q_core_148 = ~(input_a[30] ^ input_a[7]);
  assign popcount32_k31q_core_156 = ~input_a[8];
  assign popcount32_k31q_core_158 = ~(input_a[27] | input_a[4]);
  assign popcount32_k31q_core_159 = ~(input_a[1] | input_a[3]);
  assign popcount32_k31q_core_160 = ~input_a[30];
  assign popcount32_k31q_core_161 = ~(input_a[11] ^ input_a[3]);
  assign popcount32_k31q_core_162 = input_a[15] & input_a[17];
  assign popcount32_k31q_core_163 = ~(input_a[7] & input_a[27]);
  assign popcount32_k31q_core_166 = ~(input_a[22] ^ input_a[15]);
  assign popcount32_k31q_core_167 = ~input_a[8];
  assign popcount32_k31q_core_168 = ~(input_a[26] & input_a[19]);
  assign popcount32_k31q_core_169 = ~(input_a[21] ^ input_a[19]);
  assign popcount32_k31q_core_170 = input_a[27] ^ input_a[26];
  assign popcount32_k31q_core_171 = ~(input_a[8] | input_a[15]);
  assign popcount32_k31q_core_176 = input_a[14] ^ input_a[25];
  assign popcount32_k31q_core_177 = input_a[16] | input_a[31];
  assign popcount32_k31q_core_178 = input_a[12] | input_a[31];
  assign popcount32_k31q_core_179_not = ~input_a[5];
  assign popcount32_k31q_core_180 = input_a[26] & input_a[4];
  assign popcount32_k31q_core_182 = ~(input_a[17] | input_a[0]);
  assign popcount32_k31q_core_184 = input_a[15] ^ input_a[23];
  assign popcount32_k31q_core_185 = ~(input_a[20] & input_a[28]);
  assign popcount32_k31q_core_186 = ~(input_a[14] | input_a[28]);
  assign popcount32_k31q_core_187 = ~(input_a[10] & input_a[31]);
  assign popcount32_k31q_core_188 = ~(input_a[19] | input_a[26]);
  assign popcount32_k31q_core_189 = input_a[13] & input_a[10];
  assign popcount32_k31q_core_190 = ~(input_a[19] | input_a[1]);
  assign popcount32_k31q_core_194 = ~(input_a[24] & input_a[25]);
  assign popcount32_k31q_core_195 = ~(input_a[11] | input_a[5]);
  assign popcount32_k31q_core_196 = ~(input_a[28] ^ input_a[27]);
  assign popcount32_k31q_core_197 = input_a[13] | input_a[10];
  assign popcount32_k31q_core_198 = ~(input_a[6] ^ input_a[10]);
  assign popcount32_k31q_core_199 = input_a[1] ^ input_a[5];
  assign popcount32_k31q_core_200 = ~(input_a[23] ^ input_a[11]);
  assign popcount32_k31q_core_201 = ~input_a[20];
  assign popcount32_k31q_core_202 = ~(input_a[7] & input_a[9]);
  assign popcount32_k31q_core_204 = ~(input_a[2] ^ input_a[17]);
  assign popcount32_k31q_core_206 = ~input_a[5];
  assign popcount32_k31q_core_208 = ~(input_a[14] & input_a[26]);
  assign popcount32_k31q_core_209 = input_a[25] | input_a[5];
  assign popcount32_k31q_core_211 = ~(input_a[26] ^ input_a[24]);
  assign popcount32_k31q_core_212 = input_a[25] & input_a[5];
  assign popcount32_k31q_core_213 = input_a[20] | input_a[24];
  assign popcount32_k31q_core_215 = ~(input_a[20] & input_a[9]);
  assign popcount32_k31q_core_216 = ~(input_a[12] & input_a[8]);
  assign popcount32_k31q_core_218 = input_a[12] | input_a[29];
  assign popcount32_k31q_core_219 = input_a[14] & input_a[22];
  assign popcount32_k31q_core_220 = ~(input_a[1] ^ input_a[10]);
  assign popcount32_k31q_core_223 = ~(input_a[1] | input_a[25]);
  assign popcount32_k31q_core_224 = ~(input_a[27] ^ input_a[28]);
  assign popcount32_k31q_core_225 = ~input_a[18];

  assign popcount32_k31q_out[0] = 1'b1;
  assign popcount32_k31q_out[1] = input_a[4];
  assign popcount32_k31q_out[2] = input_a[20];
  assign popcount32_k31q_out[3] = input_a[14];
  assign popcount32_k31q_out[4] = 1'b0;
  assign popcount32_k31q_out[5] = input_a[11];
endmodule