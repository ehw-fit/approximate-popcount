// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=7.73467
// WCE=31.0
// EP=0.968517%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount39_m5xf(input [38:0] input_a, output [5:0] popcount39_m5xf_out);
  wire popcount39_m5xf_core_042;
  wire popcount39_m5xf_core_044;
  wire popcount39_m5xf_core_049;
  wire popcount39_m5xf_core_051;
  wire popcount39_m5xf_core_052;
  wire popcount39_m5xf_core_053;
  wire popcount39_m5xf_core_054;
  wire popcount39_m5xf_core_057;
  wire popcount39_m5xf_core_058;
  wire popcount39_m5xf_core_059;
  wire popcount39_m5xf_core_060;
  wire popcount39_m5xf_core_061;
  wire popcount39_m5xf_core_062;
  wire popcount39_m5xf_core_063;
  wire popcount39_m5xf_core_066;
  wire popcount39_m5xf_core_067;
  wire popcount39_m5xf_core_068;
  wire popcount39_m5xf_core_071;
  wire popcount39_m5xf_core_073;
  wire popcount39_m5xf_core_074;
  wire popcount39_m5xf_core_075;
  wire popcount39_m5xf_core_076;
  wire popcount39_m5xf_core_077;
  wire popcount39_m5xf_core_079;
  wire popcount39_m5xf_core_081;
  wire popcount39_m5xf_core_084;
  wire popcount39_m5xf_core_085;
  wire popcount39_m5xf_core_086;
  wire popcount39_m5xf_core_087;
  wire popcount39_m5xf_core_089;
  wire popcount39_m5xf_core_091;
  wire popcount39_m5xf_core_092;
  wire popcount39_m5xf_core_093;
  wire popcount39_m5xf_core_094;
  wire popcount39_m5xf_core_096;
  wire popcount39_m5xf_core_097;
  wire popcount39_m5xf_core_098;
  wire popcount39_m5xf_core_099;
  wire popcount39_m5xf_core_100;
  wire popcount39_m5xf_core_101;
  wire popcount39_m5xf_core_102;
  wire popcount39_m5xf_core_103;
  wire popcount39_m5xf_core_104_not;
  wire popcount39_m5xf_core_105;
  wire popcount39_m5xf_core_106;
  wire popcount39_m5xf_core_107;
  wire popcount39_m5xf_core_109;
  wire popcount39_m5xf_core_112;
  wire popcount39_m5xf_core_113;
  wire popcount39_m5xf_core_115;
  wire popcount39_m5xf_core_116;
  wire popcount39_m5xf_core_117;
  wire popcount39_m5xf_core_118;
  wire popcount39_m5xf_core_119;
  wire popcount39_m5xf_core_121;
  wire popcount39_m5xf_core_122;
  wire popcount39_m5xf_core_124;
  wire popcount39_m5xf_core_125;
  wire popcount39_m5xf_core_128;
  wire popcount39_m5xf_core_129;
  wire popcount39_m5xf_core_131_not;
  wire popcount39_m5xf_core_132;
  wire popcount39_m5xf_core_133;
  wire popcount39_m5xf_core_134;
  wire popcount39_m5xf_core_136;
  wire popcount39_m5xf_core_137;
  wire popcount39_m5xf_core_138;
  wire popcount39_m5xf_core_141;
  wire popcount39_m5xf_core_142_not;
  wire popcount39_m5xf_core_143;
  wire popcount39_m5xf_core_144;
  wire popcount39_m5xf_core_145;
  wire popcount39_m5xf_core_146;
  wire popcount39_m5xf_core_147;
  wire popcount39_m5xf_core_148;
  wire popcount39_m5xf_core_149;
  wire popcount39_m5xf_core_150;
  wire popcount39_m5xf_core_151;
  wire popcount39_m5xf_core_152;
  wire popcount39_m5xf_core_153;
  wire popcount39_m5xf_core_154;
  wire popcount39_m5xf_core_156;
  wire popcount39_m5xf_core_157;
  wire popcount39_m5xf_core_159;
  wire popcount39_m5xf_core_161;
  wire popcount39_m5xf_core_164;
  wire popcount39_m5xf_core_165;
  wire popcount39_m5xf_core_166;
  wire popcount39_m5xf_core_169;
  wire popcount39_m5xf_core_177;
  wire popcount39_m5xf_core_178;
  wire popcount39_m5xf_core_179;
  wire popcount39_m5xf_core_182;
  wire popcount39_m5xf_core_183;
  wire popcount39_m5xf_core_185;
  wire popcount39_m5xf_core_187;
  wire popcount39_m5xf_core_188;
  wire popcount39_m5xf_core_190;
  wire popcount39_m5xf_core_192;
  wire popcount39_m5xf_core_193;
  wire popcount39_m5xf_core_197;
  wire popcount39_m5xf_core_198;
  wire popcount39_m5xf_core_201;
  wire popcount39_m5xf_core_203_not;
  wire popcount39_m5xf_core_204;
  wire popcount39_m5xf_core_205;
  wire popcount39_m5xf_core_208;
  wire popcount39_m5xf_core_209;
  wire popcount39_m5xf_core_210;
  wire popcount39_m5xf_core_214;
  wire popcount39_m5xf_core_215;
  wire popcount39_m5xf_core_218;
  wire popcount39_m5xf_core_219;
  wire popcount39_m5xf_core_220;
  wire popcount39_m5xf_core_222;
  wire popcount39_m5xf_core_223_not;
  wire popcount39_m5xf_core_224;
  wire popcount39_m5xf_core_225;
  wire popcount39_m5xf_core_226;
  wire popcount39_m5xf_core_227;
  wire popcount39_m5xf_core_228;
  wire popcount39_m5xf_core_229;
  wire popcount39_m5xf_core_232;
  wire popcount39_m5xf_core_233;
  wire popcount39_m5xf_core_235;
  wire popcount39_m5xf_core_236;
  wire popcount39_m5xf_core_238;
  wire popcount39_m5xf_core_240;
  wire popcount39_m5xf_core_244;
  wire popcount39_m5xf_core_245;
  wire popcount39_m5xf_core_246;
  wire popcount39_m5xf_core_247;
  wire popcount39_m5xf_core_250;
  wire popcount39_m5xf_core_252_not;
  wire popcount39_m5xf_core_253;
  wire popcount39_m5xf_core_255;
  wire popcount39_m5xf_core_257;
  wire popcount39_m5xf_core_259;
  wire popcount39_m5xf_core_262;
  wire popcount39_m5xf_core_264_not;
  wire popcount39_m5xf_core_267;
  wire popcount39_m5xf_core_268;
  wire popcount39_m5xf_core_269;
  wire popcount39_m5xf_core_271;
  wire popcount39_m5xf_core_272;
  wire popcount39_m5xf_core_273;
  wire popcount39_m5xf_core_274;
  wire popcount39_m5xf_core_276;
  wire popcount39_m5xf_core_277;
  wire popcount39_m5xf_core_278;
  wire popcount39_m5xf_core_280;
  wire popcount39_m5xf_core_282;
  wire popcount39_m5xf_core_283;
  wire popcount39_m5xf_core_284;
  wire popcount39_m5xf_core_286;
  wire popcount39_m5xf_core_288;
  wire popcount39_m5xf_core_291;
  wire popcount39_m5xf_core_292;
  wire popcount39_m5xf_core_294;
  wire popcount39_m5xf_core_295;
  wire popcount39_m5xf_core_296;
  wire popcount39_m5xf_core_298;
  wire popcount39_m5xf_core_299;
  wire popcount39_m5xf_core_300;
  wire popcount39_m5xf_core_303;
  wire popcount39_m5xf_core_304;

  assign popcount39_m5xf_core_042 = input_a[21] ^ input_a[4];
  assign popcount39_m5xf_core_044 = input_a[21] & input_a[26];
  assign popcount39_m5xf_core_049 = ~input_a[20];
  assign popcount39_m5xf_core_051 = input_a[26] & input_a[26];
  assign popcount39_m5xf_core_052 = ~input_a[14];
  assign popcount39_m5xf_core_053 = ~input_a[9];
  assign popcount39_m5xf_core_054 = ~input_a[27];
  assign popcount39_m5xf_core_057 = ~(input_a[36] & input_a[18]);
  assign popcount39_m5xf_core_058 = ~input_a[27];
  assign popcount39_m5xf_core_059 = ~(input_a[20] ^ input_a[0]);
  assign popcount39_m5xf_core_060 = ~(input_a[36] & input_a[16]);
  assign popcount39_m5xf_core_061 = input_a[3] | input_a[23];
  assign popcount39_m5xf_core_062 = ~input_a[12];
  assign popcount39_m5xf_core_063 = input_a[9] & input_a[16];
  assign popcount39_m5xf_core_066 = ~(input_a[30] & input_a[8]);
  assign popcount39_m5xf_core_067 = input_a[30] & input_a[21];
  assign popcount39_m5xf_core_068 = ~(input_a[4] ^ input_a[12]);
  assign popcount39_m5xf_core_071 = input_a[34] ^ input_a[10];
  assign popcount39_m5xf_core_073 = ~(input_a[19] ^ input_a[26]);
  assign popcount39_m5xf_core_074 = input_a[28] ^ input_a[25];
  assign popcount39_m5xf_core_075 = ~(input_a[10] & input_a[32]);
  assign popcount39_m5xf_core_076 = ~input_a[24];
  assign popcount39_m5xf_core_077 = input_a[38] | input_a[34];
  assign popcount39_m5xf_core_079 = input_a[2] & input_a[30];
  assign popcount39_m5xf_core_081 = ~input_a[33];
  assign popcount39_m5xf_core_084 = ~(input_a[29] & input_a[18]);
  assign popcount39_m5xf_core_085 = ~(input_a[23] ^ input_a[21]);
  assign popcount39_m5xf_core_086 = ~input_a[12];
  assign popcount39_m5xf_core_087 = ~(input_a[22] | input_a[28]);
  assign popcount39_m5xf_core_089 = ~(input_a[30] | input_a[8]);
  assign popcount39_m5xf_core_091 = ~(input_a[6] & input_a[9]);
  assign popcount39_m5xf_core_092 = input_a[3] & input_a[2];
  assign popcount39_m5xf_core_093 = input_a[27] & input_a[29];
  assign popcount39_m5xf_core_094 = ~(input_a[37] & input_a[34]);
  assign popcount39_m5xf_core_096 = input_a[16] | input_a[16];
  assign popcount39_m5xf_core_097 = input_a[23] | input_a[31];
  assign popcount39_m5xf_core_098 = ~(input_a[18] & input_a[18]);
  assign popcount39_m5xf_core_099 = ~input_a[24];
  assign popcount39_m5xf_core_100 = ~(input_a[30] | input_a[3]);
  assign popcount39_m5xf_core_101 = input_a[8] & input_a[36];
  assign popcount39_m5xf_core_102 = input_a[6] | input_a[19];
  assign popcount39_m5xf_core_103 = input_a[32] & input_a[25];
  assign popcount39_m5xf_core_104_not = ~input_a[32];
  assign popcount39_m5xf_core_105 = ~(input_a[11] & input_a[30]);
  assign popcount39_m5xf_core_106 = ~(input_a[30] | input_a[29]);
  assign popcount39_m5xf_core_107 = input_a[22] ^ input_a[16];
  assign popcount39_m5xf_core_109 = ~(input_a[5] ^ input_a[29]);
  assign popcount39_m5xf_core_112 = ~(input_a[36] | input_a[24]);
  assign popcount39_m5xf_core_113 = input_a[5] | input_a[8];
  assign popcount39_m5xf_core_115 = input_a[6] ^ input_a[23];
  assign popcount39_m5xf_core_116 = ~(input_a[30] | input_a[31]);
  assign popcount39_m5xf_core_117 = ~input_a[29];
  assign popcount39_m5xf_core_118 = ~(input_a[2] | input_a[3]);
  assign popcount39_m5xf_core_119 = input_a[7] | input_a[37];
  assign popcount39_m5xf_core_121 = ~input_a[19];
  assign popcount39_m5xf_core_122 = ~(input_a[20] ^ input_a[24]);
  assign popcount39_m5xf_core_124 = input_a[3] | input_a[26];
  assign popcount39_m5xf_core_125 = ~(input_a[1] & input_a[31]);
  assign popcount39_m5xf_core_128 = ~(input_a[2] ^ input_a[15]);
  assign popcount39_m5xf_core_129 = input_a[23] | input_a[10];
  assign popcount39_m5xf_core_131_not = ~input_a[38];
  assign popcount39_m5xf_core_132 = ~(input_a[30] ^ input_a[29]);
  assign popcount39_m5xf_core_133 = input_a[5] | input_a[37];
  assign popcount39_m5xf_core_134 = ~input_a[2];
  assign popcount39_m5xf_core_136 = ~input_a[32];
  assign popcount39_m5xf_core_137 = input_a[18] | input_a[0];
  assign popcount39_m5xf_core_138 = ~(input_a[30] | input_a[29]);
  assign popcount39_m5xf_core_141 = ~input_a[25];
  assign popcount39_m5xf_core_142_not = ~input_a[30];
  assign popcount39_m5xf_core_143 = ~(input_a[6] | input_a[25]);
  assign popcount39_m5xf_core_144 = ~(input_a[12] ^ input_a[1]);
  assign popcount39_m5xf_core_145 = ~(input_a[36] | input_a[38]);
  assign popcount39_m5xf_core_146 = ~(input_a[1] ^ input_a[14]);
  assign popcount39_m5xf_core_147 = input_a[19] & input_a[21];
  assign popcount39_m5xf_core_148 = input_a[30] | input_a[26];
  assign popcount39_m5xf_core_149 = input_a[16] ^ input_a[7];
  assign popcount39_m5xf_core_150 = input_a[1] & input_a[5];
  assign popcount39_m5xf_core_151 = ~input_a[27];
  assign popcount39_m5xf_core_152 = ~(input_a[13] ^ input_a[21]);
  assign popcount39_m5xf_core_153 = input_a[11] | input_a[13];
  assign popcount39_m5xf_core_154 = input_a[8] ^ input_a[37];
  assign popcount39_m5xf_core_156 = input_a[38] ^ input_a[7];
  assign popcount39_m5xf_core_157 = input_a[3] | input_a[37];
  assign popcount39_m5xf_core_159 = input_a[14] & input_a[8];
  assign popcount39_m5xf_core_161 = ~input_a[8];
  assign popcount39_m5xf_core_164 = input_a[36] & input_a[2];
  assign popcount39_m5xf_core_165 = input_a[26] ^ input_a[36];
  assign popcount39_m5xf_core_166 = ~input_a[28];
  assign popcount39_m5xf_core_169 = input_a[2] | input_a[15];
  assign popcount39_m5xf_core_177 = ~input_a[1];
  assign popcount39_m5xf_core_178 = input_a[14] | input_a[18];
  assign popcount39_m5xf_core_179 = ~(input_a[25] ^ input_a[37]);
  assign popcount39_m5xf_core_182 = input_a[16] & input_a[38];
  assign popcount39_m5xf_core_183 = ~(input_a[13] & input_a[14]);
  assign popcount39_m5xf_core_185 = input_a[28] & input_a[34];
  assign popcount39_m5xf_core_187 = input_a[12] | input_a[24];
  assign popcount39_m5xf_core_188 = input_a[15] & input_a[16];
  assign popcount39_m5xf_core_190 = ~(input_a[9] & input_a[8]);
  assign popcount39_m5xf_core_192 = ~(input_a[15] ^ input_a[33]);
  assign popcount39_m5xf_core_193 = ~(input_a[38] | input_a[6]);
  assign popcount39_m5xf_core_197 = input_a[9] ^ input_a[3];
  assign popcount39_m5xf_core_198 = ~(input_a[2] ^ input_a[17]);
  assign popcount39_m5xf_core_201 = ~(input_a[24] ^ input_a[2]);
  assign popcount39_m5xf_core_203_not = ~input_a[23];
  assign popcount39_m5xf_core_204 = ~(input_a[32] & input_a[25]);
  assign popcount39_m5xf_core_205 = input_a[23] ^ input_a[3];
  assign popcount39_m5xf_core_208 = input_a[26] | input_a[28];
  assign popcount39_m5xf_core_209 = ~input_a[5];
  assign popcount39_m5xf_core_210 = input_a[9] | input_a[26];
  assign popcount39_m5xf_core_214 = ~input_a[28];
  assign popcount39_m5xf_core_215 = input_a[6] & input_a[18];
  assign popcount39_m5xf_core_218 = ~(input_a[27] & input_a[5]);
  assign popcount39_m5xf_core_219 = ~(input_a[12] | input_a[21]);
  assign popcount39_m5xf_core_220 = ~input_a[26];
  assign popcount39_m5xf_core_222 = input_a[37] | input_a[19];
  assign popcount39_m5xf_core_223_not = ~input_a[36];
  assign popcount39_m5xf_core_224 = ~(input_a[5] & input_a[5]);
  assign popcount39_m5xf_core_225 = input_a[13] ^ input_a[28];
  assign popcount39_m5xf_core_226 = input_a[38] | input_a[8];
  assign popcount39_m5xf_core_227 = ~(input_a[17] & input_a[24]);
  assign popcount39_m5xf_core_228 = input_a[4] & input_a[31];
  assign popcount39_m5xf_core_229 = input_a[26] | input_a[20];
  assign popcount39_m5xf_core_232 = input_a[29] | input_a[27];
  assign popcount39_m5xf_core_233 = ~(input_a[35] ^ input_a[1]);
  assign popcount39_m5xf_core_235 = ~(input_a[3] & input_a[15]);
  assign popcount39_m5xf_core_236 = ~(input_a[26] ^ input_a[25]);
  assign popcount39_m5xf_core_238 = input_a[5] | input_a[7];
  assign popcount39_m5xf_core_240 = input_a[9] ^ input_a[28];
  assign popcount39_m5xf_core_244 = input_a[10] | input_a[18];
  assign popcount39_m5xf_core_245 = ~input_a[36];
  assign popcount39_m5xf_core_246 = ~(input_a[1] | input_a[14]);
  assign popcount39_m5xf_core_247 = input_a[36] ^ input_a[17];
  assign popcount39_m5xf_core_250 = ~input_a[21];
  assign popcount39_m5xf_core_252_not = ~input_a[17];
  assign popcount39_m5xf_core_253 = input_a[15] & input_a[31];
  assign popcount39_m5xf_core_255 = input_a[30] & input_a[6];
  assign popcount39_m5xf_core_257 = input_a[32] & input_a[15];
  assign popcount39_m5xf_core_259 = input_a[33] | input_a[1];
  assign popcount39_m5xf_core_262 = ~(input_a[18] | input_a[25]);
  assign popcount39_m5xf_core_264_not = ~input_a[3];
  assign popcount39_m5xf_core_267 = ~(input_a[27] & input_a[24]);
  assign popcount39_m5xf_core_268 = ~input_a[19];
  assign popcount39_m5xf_core_269 = input_a[31] | input_a[23];
  assign popcount39_m5xf_core_271 = input_a[9] & input_a[17];
  assign popcount39_m5xf_core_272 = input_a[26] | input_a[9];
  assign popcount39_m5xf_core_273 = ~(input_a[36] | input_a[35]);
  assign popcount39_m5xf_core_274 = input_a[4] & input_a[7];
  assign popcount39_m5xf_core_276 = input_a[11] | input_a[0];
  assign popcount39_m5xf_core_277 = ~(input_a[34] & input_a[8]);
  assign popcount39_m5xf_core_278 = input_a[17] | input_a[15];
  assign popcount39_m5xf_core_280 = ~(input_a[34] ^ input_a[23]);
  assign popcount39_m5xf_core_282 = input_a[33] & input_a[28];
  assign popcount39_m5xf_core_283 = input_a[18] | input_a[10];
  assign popcount39_m5xf_core_284 = input_a[5] & input_a[0];
  assign popcount39_m5xf_core_286 = ~(input_a[8] & input_a[14]);
  assign popcount39_m5xf_core_288 = ~(input_a[16] & input_a[11]);
  assign popcount39_m5xf_core_291 = ~(input_a[1] ^ input_a[15]);
  assign popcount39_m5xf_core_292 = input_a[1] | input_a[19];
  assign popcount39_m5xf_core_294 = ~input_a[10];
  assign popcount39_m5xf_core_295 = ~(input_a[27] ^ input_a[36]);
  assign popcount39_m5xf_core_296 = ~(input_a[14] & input_a[24]);
  assign popcount39_m5xf_core_298 = input_a[9] | input_a[0];
  assign popcount39_m5xf_core_299 = ~(input_a[22] ^ input_a[13]);
  assign popcount39_m5xf_core_300 = input_a[37] & input_a[37];
  assign popcount39_m5xf_core_303 = input_a[29] & input_a[38];
  assign popcount39_m5xf_core_304 = input_a[1] | input_a[31];

  assign popcount39_m5xf_out[0] = input_a[29];
  assign popcount39_m5xf_out[1] = input_a[7];
  assign popcount39_m5xf_out[2] = 1'b1;
  assign popcount39_m5xf_out[3] = input_a[8];
  assign popcount39_m5xf_out[4] = input_a[14];
  assign popcount39_m5xf_out[5] = 1'b0;
endmodule