// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.39972
// WCE=10.0
// EP=0.78055%
// Printed PDK parameters:
//  Area=47229198.0
//  Delay=59015508.0
//  Power=2207000.0

module popcount28_jvgw(input [27:0] input_a, output [4:0] popcount28_jvgw_out);
  wire popcount28_jvgw_core_030_not;
  wire popcount28_jvgw_core_031;
  wire popcount28_jvgw_core_032;
  wire popcount28_jvgw_core_033;
  wire popcount28_jvgw_core_036;
  wire popcount28_jvgw_core_037;
  wire popcount28_jvgw_core_038;
  wire popcount28_jvgw_core_039;
  wire popcount28_jvgw_core_041;
  wire popcount28_jvgw_core_042;
  wire popcount28_jvgw_core_044;
  wire popcount28_jvgw_core_045;
  wire popcount28_jvgw_core_047;
  wire popcount28_jvgw_core_048;
  wire popcount28_jvgw_core_049;
  wire popcount28_jvgw_core_050;
  wire popcount28_jvgw_core_052;
  wire popcount28_jvgw_core_055;
  wire popcount28_jvgw_core_056;
  wire popcount28_jvgw_core_057;
  wire popcount28_jvgw_core_058;
  wire popcount28_jvgw_core_059;
  wire popcount28_jvgw_core_060;
  wire popcount28_jvgw_core_061;
  wire popcount28_jvgw_core_062;
  wire popcount28_jvgw_core_063;
  wire popcount28_jvgw_core_065;
  wire popcount28_jvgw_core_066;
  wire popcount28_jvgw_core_067;
  wire popcount28_jvgw_core_068;
  wire popcount28_jvgw_core_070;
  wire popcount28_jvgw_core_071;
  wire popcount28_jvgw_core_072;
  wire popcount28_jvgw_core_073;
  wire popcount28_jvgw_core_074;
  wire popcount28_jvgw_core_077;
  wire popcount28_jvgw_core_078;
  wire popcount28_jvgw_core_079;
  wire popcount28_jvgw_core_081;
  wire popcount28_jvgw_core_084;
  wire popcount28_jvgw_core_085;
  wire popcount28_jvgw_core_088;
  wire popcount28_jvgw_core_089;
  wire popcount28_jvgw_core_090;
  wire popcount28_jvgw_core_091;
  wire popcount28_jvgw_core_092;
  wire popcount28_jvgw_core_093;
  wire popcount28_jvgw_core_094;
  wire popcount28_jvgw_core_095;
  wire popcount28_jvgw_core_096;
  wire popcount28_jvgw_core_097;
  wire popcount28_jvgw_core_098;
  wire popcount28_jvgw_core_099;
  wire popcount28_jvgw_core_101;
  wire popcount28_jvgw_core_103_not;
  wire popcount28_jvgw_core_104;
  wire popcount28_jvgw_core_105;
  wire popcount28_jvgw_core_106;
  wire popcount28_jvgw_core_107;
  wire popcount28_jvgw_core_108;
  wire popcount28_jvgw_core_111;
  wire popcount28_jvgw_core_112;
  wire popcount28_jvgw_core_113;
  wire popcount28_jvgw_core_114;
  wire popcount28_jvgw_core_116;
  wire popcount28_jvgw_core_117;
  wire popcount28_jvgw_core_118;
  wire popcount28_jvgw_core_119;
  wire popcount28_jvgw_core_122;
  wire popcount28_jvgw_core_123;
  wire popcount28_jvgw_core_124;
  wire popcount28_jvgw_core_126;
  wire popcount28_jvgw_core_128;
  wire popcount28_jvgw_core_131;
  wire popcount28_jvgw_core_135;
  wire popcount28_jvgw_core_138;
  wire popcount28_jvgw_core_139;
  wire popcount28_jvgw_core_141;
  wire popcount28_jvgw_core_142;
  wire popcount28_jvgw_core_144;
  wire popcount28_jvgw_core_146;
  wire popcount28_jvgw_core_148_not;
  wire popcount28_jvgw_core_150;
  wire popcount28_jvgw_core_151;
  wire popcount28_jvgw_core_152;
  wire popcount28_jvgw_core_153;
  wire popcount28_jvgw_core_155;
  wire popcount28_jvgw_core_159;
  wire popcount28_jvgw_core_160;
  wire popcount28_jvgw_core_161;
  wire popcount28_jvgw_core_163;
  wire popcount28_jvgw_core_164;
  wire popcount28_jvgw_core_165;
  wire popcount28_jvgw_core_166;
  wire popcount28_jvgw_core_167;
  wire popcount28_jvgw_core_168;
  wire popcount28_jvgw_core_169;
  wire popcount28_jvgw_core_170;
  wire popcount28_jvgw_core_171;
  wire popcount28_jvgw_core_172;
  wire popcount28_jvgw_core_173;
  wire popcount28_jvgw_core_174;
  wire popcount28_jvgw_core_176;
  wire popcount28_jvgw_core_177;
  wire popcount28_jvgw_core_178;
  wire popcount28_jvgw_core_179;
  wire popcount28_jvgw_core_181_not;
  wire popcount28_jvgw_core_182;
  wire popcount28_jvgw_core_183;
  wire popcount28_jvgw_core_185;
  wire popcount28_jvgw_core_187;
  wire popcount28_jvgw_core_188;
  wire popcount28_jvgw_core_189;
  wire popcount28_jvgw_core_190;
  wire popcount28_jvgw_core_191;
  wire popcount28_jvgw_core_192;
  wire popcount28_jvgw_core_193;
  wire popcount28_jvgw_core_194;
  wire popcount28_jvgw_core_195;
  wire popcount28_jvgw_core_196;
  wire popcount28_jvgw_core_198;

  assign popcount28_jvgw_core_030_not = ~input_a[6];
  assign popcount28_jvgw_core_031 = input_a[25] & input_a[2];
  assign popcount28_jvgw_core_032 = input_a[9] & input_a[26];
  assign popcount28_jvgw_core_033 = ~(input_a[20] & input_a[1]);
  assign popcount28_jvgw_core_036 = ~input_a[21];
  assign popcount28_jvgw_core_037 = input_a[3] & input_a[4];
  assign popcount28_jvgw_core_038 = ~(input_a[12] | input_a[14]);
  assign popcount28_jvgw_core_039 = input_a[0] & input_a[1];
  assign popcount28_jvgw_core_041 = input_a[25] & input_a[15];
  assign popcount28_jvgw_core_042 = popcount28_jvgw_core_037 | popcount28_jvgw_core_039;
  assign popcount28_jvgw_core_044 = popcount28_jvgw_core_042 ^ input_a[6];
  assign popcount28_jvgw_core_045 = popcount28_jvgw_core_042 & input_a[6];
  assign popcount28_jvgw_core_047 = input_a[8] | input_a[24];
  assign popcount28_jvgw_core_048 = ~(input_a[26] & input_a[12]);
  assign popcount28_jvgw_core_049 = popcount28_jvgw_core_031 ^ popcount28_jvgw_core_044;
  assign popcount28_jvgw_core_050 = popcount28_jvgw_core_031 & popcount28_jvgw_core_044;
  assign popcount28_jvgw_core_052 = ~input_a[25];
  assign popcount28_jvgw_core_055 = input_a[11] & input_a[13];
  assign popcount28_jvgw_core_056 = popcount28_jvgw_core_045 | popcount28_jvgw_core_050;
  assign popcount28_jvgw_core_057 = input_a[8] & input_a[5];
  assign popcount28_jvgw_core_058 = ~(input_a[5] ^ input_a[16]);
  assign popcount28_jvgw_core_059 = input_a[8] | input_a[9];
  assign popcount28_jvgw_core_060 = input_a[8] & input_a[9];
  assign popcount28_jvgw_core_061 = ~input_a[27];
  assign popcount28_jvgw_core_062 = input_a[7] & popcount28_jvgw_core_059;
  assign popcount28_jvgw_core_063 = popcount28_jvgw_core_060 | popcount28_jvgw_core_062;
  assign popcount28_jvgw_core_065 = input_a[10] | input_a[11];
  assign popcount28_jvgw_core_066 = input_a[10] & input_a[11];
  assign popcount28_jvgw_core_067 = input_a[12] ^ input_a[13];
  assign popcount28_jvgw_core_068 = input_a[12] & input_a[13];
  assign popcount28_jvgw_core_070 = popcount28_jvgw_core_065 & popcount28_jvgw_core_067;
  assign popcount28_jvgw_core_071 = popcount28_jvgw_core_066 ^ popcount28_jvgw_core_068;
  assign popcount28_jvgw_core_072 = popcount28_jvgw_core_066 & popcount28_jvgw_core_068;
  assign popcount28_jvgw_core_073 = popcount28_jvgw_core_071 | popcount28_jvgw_core_070;
  assign popcount28_jvgw_core_074 = ~(input_a[7] ^ input_a[26]);
  assign popcount28_jvgw_core_077 = ~(input_a[21] ^ input_a[8]);
  assign popcount28_jvgw_core_078 = popcount28_jvgw_core_063 ^ popcount28_jvgw_core_073;
  assign popcount28_jvgw_core_079 = popcount28_jvgw_core_063 & popcount28_jvgw_core_073;
  assign popcount28_jvgw_core_081 = ~input_a[17];
  assign popcount28_jvgw_core_084 = input_a[6] & input_a[5];
  assign popcount28_jvgw_core_085 = popcount28_jvgw_core_072 | popcount28_jvgw_core_079;
  assign popcount28_jvgw_core_088 = input_a[23] & input_a[16];
  assign popcount28_jvgw_core_089 = input_a[27] & input_a[20];
  assign popcount28_jvgw_core_090 = popcount28_jvgw_core_049 ^ popcount28_jvgw_core_078;
  assign popcount28_jvgw_core_091 = popcount28_jvgw_core_049 & popcount28_jvgw_core_078;
  assign popcount28_jvgw_core_092 = popcount28_jvgw_core_090 ^ popcount28_jvgw_core_089;
  assign popcount28_jvgw_core_093 = popcount28_jvgw_core_090 & popcount28_jvgw_core_089;
  assign popcount28_jvgw_core_094 = popcount28_jvgw_core_091 | popcount28_jvgw_core_093;
  assign popcount28_jvgw_core_095 = popcount28_jvgw_core_056 ^ popcount28_jvgw_core_085;
  assign popcount28_jvgw_core_096 = popcount28_jvgw_core_056 & popcount28_jvgw_core_085;
  assign popcount28_jvgw_core_097 = popcount28_jvgw_core_095 ^ popcount28_jvgw_core_094;
  assign popcount28_jvgw_core_098 = popcount28_jvgw_core_095 & popcount28_jvgw_core_094;
  assign popcount28_jvgw_core_099 = popcount28_jvgw_core_096 | popcount28_jvgw_core_098;
  assign popcount28_jvgw_core_101 = input_a[27] | input_a[5];
  assign popcount28_jvgw_core_103_not = ~input_a[3];
  assign popcount28_jvgw_core_104 = input_a[0] | input_a[5];
  assign popcount28_jvgw_core_105 = ~(input_a[5] | input_a[13]);
  assign popcount28_jvgw_core_106 = input_a[15] & input_a[16];
  assign popcount28_jvgw_core_107 = input_a[16] | input_a[3];
  assign popcount28_jvgw_core_108 = ~(input_a[25] ^ input_a[27]);
  assign popcount28_jvgw_core_111 = input_a[17] ^ input_a[18];
  assign popcount28_jvgw_core_112 = input_a[17] & input_a[18];
  assign popcount28_jvgw_core_113 = input_a[19] | input_a[14];
  assign popcount28_jvgw_core_114 = input_a[19] & input_a[14];
  assign popcount28_jvgw_core_116 = popcount28_jvgw_core_111 & popcount28_jvgw_core_113;
  assign popcount28_jvgw_core_117 = popcount28_jvgw_core_112 ^ popcount28_jvgw_core_114;
  assign popcount28_jvgw_core_118 = popcount28_jvgw_core_112 & popcount28_jvgw_core_114;
  assign popcount28_jvgw_core_119 = popcount28_jvgw_core_117 | popcount28_jvgw_core_116;
  assign popcount28_jvgw_core_122 = ~(input_a[7] & input_a[5]);
  assign popcount28_jvgw_core_123 = input_a[3] & input_a[6];
  assign popcount28_jvgw_core_124 = popcount28_jvgw_core_106 ^ popcount28_jvgw_core_119;
  assign popcount28_jvgw_core_126 = ~popcount28_jvgw_core_124;
  assign popcount28_jvgw_core_128 = popcount28_jvgw_core_106 | popcount28_jvgw_core_124;
  assign popcount28_jvgw_core_131 = popcount28_jvgw_core_118 ^ popcount28_jvgw_core_128;
  assign popcount28_jvgw_core_135 = input_a[22] & input_a[23];
  assign popcount28_jvgw_core_138 = popcount28_jvgw_core_135 | input_a[5];
  assign popcount28_jvgw_core_139 = ~(input_a[10] | input_a[18]);
  assign popcount28_jvgw_core_141 = ~input_a[8];
  assign popcount28_jvgw_core_142 = ~(input_a[12] & input_a[12]);
  assign popcount28_jvgw_core_144 = ~(input_a[17] & input_a[0]);
  assign popcount28_jvgw_core_146 = ~input_a[22];
  assign popcount28_jvgw_core_148_not = ~input_a[15];
  assign popcount28_jvgw_core_150 = input_a[16] ^ input_a[9];
  assign popcount28_jvgw_core_151 = ~(input_a[4] | input_a[18]);
  assign popcount28_jvgw_core_152 = ~(input_a[8] ^ input_a[1]);
  assign popcount28_jvgw_core_153 = ~popcount28_jvgw_core_138;
  assign popcount28_jvgw_core_155 = popcount28_jvgw_core_153 ^ input_a[26];
  assign popcount28_jvgw_core_159 = input_a[27] & input_a[19];
  assign popcount28_jvgw_core_160 = input_a[26] | popcount28_jvgw_core_138;
  assign popcount28_jvgw_core_161 = ~(input_a[10] ^ input_a[20]);
  assign popcount28_jvgw_core_163 = input_a[17] ^ input_a[1];
  assign popcount28_jvgw_core_164 = input_a[24] & input_a[21];
  assign popcount28_jvgw_core_165 = popcount28_jvgw_core_126 ^ popcount28_jvgw_core_155;
  assign popcount28_jvgw_core_166 = popcount28_jvgw_core_126 & popcount28_jvgw_core_155;
  assign popcount28_jvgw_core_167 = popcount28_jvgw_core_165 ^ popcount28_jvgw_core_164;
  assign popcount28_jvgw_core_168 = popcount28_jvgw_core_165 & popcount28_jvgw_core_164;
  assign popcount28_jvgw_core_169 = popcount28_jvgw_core_166 | popcount28_jvgw_core_168;
  assign popcount28_jvgw_core_170 = popcount28_jvgw_core_131 ^ popcount28_jvgw_core_160;
  assign popcount28_jvgw_core_171 = popcount28_jvgw_core_131 & popcount28_jvgw_core_160;
  assign popcount28_jvgw_core_172 = popcount28_jvgw_core_170 ^ popcount28_jvgw_core_169;
  assign popcount28_jvgw_core_173 = popcount28_jvgw_core_170 & popcount28_jvgw_core_169;
  assign popcount28_jvgw_core_174 = popcount28_jvgw_core_171 | popcount28_jvgw_core_173;
  assign popcount28_jvgw_core_176 = ~(input_a[8] & input_a[19]);
  assign popcount28_jvgw_core_177 = popcount28_jvgw_core_118 | popcount28_jvgw_core_174;
  assign popcount28_jvgw_core_178 = input_a[17] | input_a[25];
  assign popcount28_jvgw_core_179 = input_a[8] | input_a[8];
  assign popcount28_jvgw_core_181_not = ~input_a[18];
  assign popcount28_jvgw_core_182 = popcount28_jvgw_core_092 ^ popcount28_jvgw_core_167;
  assign popcount28_jvgw_core_183 = popcount28_jvgw_core_092 & popcount28_jvgw_core_167;
  assign popcount28_jvgw_core_185 = ~(input_a[12] & input_a[17]);
  assign popcount28_jvgw_core_187 = popcount28_jvgw_core_097 ^ popcount28_jvgw_core_172;
  assign popcount28_jvgw_core_188 = popcount28_jvgw_core_097 & popcount28_jvgw_core_172;
  assign popcount28_jvgw_core_189 = popcount28_jvgw_core_187 ^ popcount28_jvgw_core_183;
  assign popcount28_jvgw_core_190 = popcount28_jvgw_core_187 & popcount28_jvgw_core_183;
  assign popcount28_jvgw_core_191 = popcount28_jvgw_core_188 | popcount28_jvgw_core_190;
  assign popcount28_jvgw_core_192 = popcount28_jvgw_core_099 ^ popcount28_jvgw_core_177;
  assign popcount28_jvgw_core_193 = popcount28_jvgw_core_099 & popcount28_jvgw_core_177;
  assign popcount28_jvgw_core_194 = popcount28_jvgw_core_192 ^ popcount28_jvgw_core_191;
  assign popcount28_jvgw_core_195 = popcount28_jvgw_core_192 & popcount28_jvgw_core_191;
  assign popcount28_jvgw_core_196 = popcount28_jvgw_core_193 | popcount28_jvgw_core_195;
  assign popcount28_jvgw_core_198 = input_a[9] | input_a[21];

  assign popcount28_jvgw_out[0] = 1'b0;
  assign popcount28_jvgw_out[1] = popcount28_jvgw_core_182;
  assign popcount28_jvgw_out[2] = popcount28_jvgw_core_189;
  assign popcount28_jvgw_out[3] = popcount28_jvgw_core_194;
  assign popcount28_jvgw_out[4] = popcount28_jvgw_core_196;
endmodule