// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.59396
// WCE=8.0
// EP=0.806483%
// Printed PDK parameters:
//  Area=70706684.0
//  Delay=74744840.0
//  Power=3592000.0

module popcount36_2fox(input [35:0] input_a, output [5:0] popcount36_2fox_out);
  wire popcount36_2fox_core_038;
  wire popcount36_2fox_core_039;
  wire popcount36_2fox_core_040;
  wire popcount36_2fox_core_041;
  wire popcount36_2fox_core_042;
  wire popcount36_2fox_core_043;
  wire popcount36_2fox_core_044;
  wire popcount36_2fox_core_045;
  wire popcount36_2fox_core_046;
  wire popcount36_2fox_core_050;
  wire popcount36_2fox_core_051;
  wire popcount36_2fox_core_052;
  wire popcount36_2fox_core_053_not;
  wire popcount36_2fox_core_054;
  wire popcount36_2fox_core_057;
  wire popcount36_2fox_core_058;
  wire popcount36_2fox_core_059;
  wire popcount36_2fox_core_060;
  wire popcount36_2fox_core_066;
  wire popcount36_2fox_core_067;
  wire popcount36_2fox_core_068;
  wire popcount36_2fox_core_069;
  wire popcount36_2fox_core_070;
  wire popcount36_2fox_core_071;
  wire popcount36_2fox_core_072;
  wire popcount36_2fox_core_073;
  wire popcount36_2fox_core_074;
  wire popcount36_2fox_core_075;
  wire popcount36_2fox_core_076;
  wire popcount36_2fox_core_079;
  wire popcount36_2fox_core_080;
  wire popcount36_2fox_core_081;
  wire popcount36_2fox_core_082;
  wire popcount36_2fox_core_083;
  wire popcount36_2fox_core_084;
  wire popcount36_2fox_core_085;
  wire popcount36_2fox_core_086;
  wire popcount36_2fox_core_087;
  wire popcount36_2fox_core_088;
  wire popcount36_2fox_core_093;
  wire popcount36_2fox_core_094;
  wire popcount36_2fox_core_096;
  wire popcount36_2fox_core_097;
  wire popcount36_2fox_core_098;
  wire popcount36_2fox_core_099;
  wire popcount36_2fox_core_100;
  wire popcount36_2fox_core_102;
  wire popcount36_2fox_core_103;
  wire popcount36_2fox_core_104;
  wire popcount36_2fox_core_106;
  wire popcount36_2fox_core_108;
  wire popcount36_2fox_core_109;
  wire popcount36_2fox_core_111;
  wire popcount36_2fox_core_113;
  wire popcount36_2fox_core_114;
  wire popcount36_2fox_core_118;
  wire popcount36_2fox_core_119;
  wire popcount36_2fox_core_120;
  wire popcount36_2fox_core_122;
  wire popcount36_2fox_core_123;
  wire popcount36_2fox_core_124;
  wire popcount36_2fox_core_125;
  wire popcount36_2fox_core_126;
  wire popcount36_2fox_core_127;
  wire popcount36_2fox_core_128;
  wire popcount36_2fox_core_129;
  wire popcount36_2fox_core_130;
  wire popcount36_2fox_core_131;
  wire popcount36_2fox_core_132;
  wire popcount36_2fox_core_133;
  wire popcount36_2fox_core_135;
  wire popcount36_2fox_core_136;
  wire popcount36_2fox_core_139;
  wire popcount36_2fox_core_140;
  wire popcount36_2fox_core_142;
  wire popcount36_2fox_core_143;
  wire popcount36_2fox_core_144;
  wire popcount36_2fox_core_145;
  wire popcount36_2fox_core_147;
  wire popcount36_2fox_core_149;
  wire popcount36_2fox_core_150;
  wire popcount36_2fox_core_151;
  wire popcount36_2fox_core_152;
  wire popcount36_2fox_core_156;
  wire popcount36_2fox_core_157;
  wire popcount36_2fox_core_158;
  wire popcount36_2fox_core_160;
  wire popcount36_2fox_core_163;
  wire popcount36_2fox_core_164;
  wire popcount36_2fox_core_165;
  wire popcount36_2fox_core_166;
  wire popcount36_2fox_core_167;
  wire popcount36_2fox_core_168;
  wire popcount36_2fox_core_169;
  wire popcount36_2fox_core_172;
  wire popcount36_2fox_core_173;
  wire popcount36_2fox_core_174;
  wire popcount36_2fox_core_175;
  wire popcount36_2fox_core_177;
  wire popcount36_2fox_core_179_not;
  wire popcount36_2fox_core_181;
  wire popcount36_2fox_core_182;
  wire popcount36_2fox_core_183;
  wire popcount36_2fox_core_185;
  wire popcount36_2fox_core_187;
  wire popcount36_2fox_core_188;
  wire popcount36_2fox_core_189;
  wire popcount36_2fox_core_190;
  wire popcount36_2fox_core_191;
  wire popcount36_2fox_core_192;
  wire popcount36_2fox_core_193;
  wire popcount36_2fox_core_194;
  wire popcount36_2fox_core_195;
  wire popcount36_2fox_core_196;
  wire popcount36_2fox_core_197;
  wire popcount36_2fox_core_198;
  wire popcount36_2fox_core_199;
  wire popcount36_2fox_core_200;
  wire popcount36_2fox_core_201;
  wire popcount36_2fox_core_202;
  wire popcount36_2fox_core_203;
  wire popcount36_2fox_core_205;
  wire popcount36_2fox_core_206;
  wire popcount36_2fox_core_207;
  wire popcount36_2fox_core_208;
  wire popcount36_2fox_core_209;
  wire popcount36_2fox_core_210;
  wire popcount36_2fox_core_211;
  wire popcount36_2fox_core_216;
  wire popcount36_2fox_core_217;
  wire popcount36_2fox_core_221;
  wire popcount36_2fox_core_222;
  wire popcount36_2fox_core_223;
  wire popcount36_2fox_core_227;
  wire popcount36_2fox_core_228;
  wire popcount36_2fox_core_230;
  wire popcount36_2fox_core_231;
  wire popcount36_2fox_core_232;
  wire popcount36_2fox_core_233;
  wire popcount36_2fox_core_234;
  wire popcount36_2fox_core_235;
  wire popcount36_2fox_core_236;
  wire popcount36_2fox_core_237;
  wire popcount36_2fox_core_238;
  wire popcount36_2fox_core_239;
  wire popcount36_2fox_core_240;
  wire popcount36_2fox_core_241;
  wire popcount36_2fox_core_242;
  wire popcount36_2fox_core_243;
  wire popcount36_2fox_core_244;
  wire popcount36_2fox_core_249;
  wire popcount36_2fox_core_251;
  wire popcount36_2fox_core_252;
  wire popcount36_2fox_core_253;
  wire popcount36_2fox_core_254;
  wire popcount36_2fox_core_255;
  wire popcount36_2fox_core_256;
  wire popcount36_2fox_core_257;
  wire popcount36_2fox_core_258;
  wire popcount36_2fox_core_259;
  wire popcount36_2fox_core_260;
  wire popcount36_2fox_core_261;
  wire popcount36_2fox_core_262;
  wire popcount36_2fox_core_263;
  wire popcount36_2fox_core_264;
  wire popcount36_2fox_core_265;
  wire popcount36_2fox_core_266;
  wire popcount36_2fox_core_269;
  wire popcount36_2fox_core_270;
  wire popcount36_2fox_core_272;
  wire popcount36_2fox_core_274;
  wire popcount36_2fox_core_275;

  assign popcount36_2fox_core_038 = input_a[0] ^ input_a[1];
  assign popcount36_2fox_core_039 = input_a[0] & input_a[1];
  assign popcount36_2fox_core_040 = input_a[2] ^ input_a[3];
  assign popcount36_2fox_core_041 = input_a[2] & input_a[3];
  assign popcount36_2fox_core_042 = popcount36_2fox_core_038 ^ popcount36_2fox_core_040;
  assign popcount36_2fox_core_043 = popcount36_2fox_core_038 & popcount36_2fox_core_040;
  assign popcount36_2fox_core_044 = popcount36_2fox_core_039 ^ popcount36_2fox_core_041;
  assign popcount36_2fox_core_045 = popcount36_2fox_core_039 & popcount36_2fox_core_041;
  assign popcount36_2fox_core_046 = popcount36_2fox_core_044 | popcount36_2fox_core_043;
  assign popcount36_2fox_core_050 = ~(input_a[32] ^ input_a[28]);
  assign popcount36_2fox_core_051 = ~(input_a[22] & input_a[6]);
  assign popcount36_2fox_core_052 = ~(input_a[14] | input_a[4]);
  assign popcount36_2fox_core_053_not = ~input_a[17];
  assign popcount36_2fox_core_054 = ~(input_a[11] & input_a[2]);
  assign popcount36_2fox_core_057 = ~input_a[4];
  assign popcount36_2fox_core_058 = ~(input_a[33] | input_a[16]);
  assign popcount36_2fox_core_059 = input_a[4] ^ input_a[7];
  assign popcount36_2fox_core_060 = input_a[4] & input_a[7];
  assign popcount36_2fox_core_066 = popcount36_2fox_core_042 ^ popcount36_2fox_core_057;
  assign popcount36_2fox_core_067 = popcount36_2fox_core_042 & popcount36_2fox_core_057;
  assign popcount36_2fox_core_068 = popcount36_2fox_core_046 ^ popcount36_2fox_core_059;
  assign popcount36_2fox_core_069 = popcount36_2fox_core_046 & popcount36_2fox_core_059;
  assign popcount36_2fox_core_070 = popcount36_2fox_core_068 ^ popcount36_2fox_core_067;
  assign popcount36_2fox_core_071 = popcount36_2fox_core_068 & popcount36_2fox_core_067;
  assign popcount36_2fox_core_072 = popcount36_2fox_core_069 | popcount36_2fox_core_071;
  assign popcount36_2fox_core_073 = popcount36_2fox_core_045 ^ popcount36_2fox_core_060;
  assign popcount36_2fox_core_074 = popcount36_2fox_core_045 & popcount36_2fox_core_060;
  assign popcount36_2fox_core_075 = popcount36_2fox_core_073 | popcount36_2fox_core_072;
  assign popcount36_2fox_core_076 = ~(input_a[32] | input_a[7]);
  assign popcount36_2fox_core_079 = ~(input_a[3] ^ input_a[17]);
  assign popcount36_2fox_core_080 = input_a[18] & input_a[19];
  assign popcount36_2fox_core_081 = input_a[9] & input_a[10];
  assign popcount36_2fox_core_082 = input_a[29] ^ input_a[7];
  assign popcount36_2fox_core_083 = input_a[11] & input_a[12];
  assign popcount36_2fox_core_084 = input_a[0] | input_a[21];
  assign popcount36_2fox_core_085 = input_a[5] & input_a[33];
  assign popcount36_2fox_core_086 = popcount36_2fox_core_081 ^ popcount36_2fox_core_083;
  assign popcount36_2fox_core_087 = popcount36_2fox_core_081 & popcount36_2fox_core_083;
  assign popcount36_2fox_core_088 = popcount36_2fox_core_086 | popcount36_2fox_core_085;
  assign popcount36_2fox_core_093 = ~(input_a[1] & input_a[18]);
  assign popcount36_2fox_core_094 = ~(input_a[27] & input_a[10]);
  assign popcount36_2fox_core_096 = input_a[2] & input_a[17];
  assign popcount36_2fox_core_097 = ~(input_a[18] & input_a[1]);
  assign popcount36_2fox_core_098 = ~(input_a[21] | input_a[11]);
  assign popcount36_2fox_core_099 = ~(input_a[34] ^ input_a[5]);
  assign popcount36_2fox_core_100 = ~(input_a[20] ^ input_a[26]);
  assign popcount36_2fox_core_102 = ~input_a[18];
  assign popcount36_2fox_core_103 = input_a[22] & input_a[11];
  assign popcount36_2fox_core_104 = input_a[22] | input_a[7];
  assign popcount36_2fox_core_106 = ~(input_a[31] & input_a[19]);
  assign popcount36_2fox_core_108 = ~(input_a[1] & input_a[2]);
  assign popcount36_2fox_core_109 = ~input_a[8];
  assign popcount36_2fox_core_111 = ~(input_a[14] ^ input_a[6]);
  assign popcount36_2fox_core_113 = ~(input_a[31] ^ input_a[26]);
  assign popcount36_2fox_core_114 = input_a[1] & input_a[19];
  assign popcount36_2fox_core_118 = ~input_a[20];
  assign popcount36_2fox_core_119 = input_a[0] | input_a[10];
  assign popcount36_2fox_core_120 = input_a[9] | input_a[29];
  assign popcount36_2fox_core_122 = input_a[32] ^ input_a[10];
  assign popcount36_2fox_core_123 = popcount36_2fox_core_066 & input_a[22];
  assign popcount36_2fox_core_124 = popcount36_2fox_core_070 ^ popcount36_2fox_core_088;
  assign popcount36_2fox_core_125 = popcount36_2fox_core_070 & popcount36_2fox_core_088;
  assign popcount36_2fox_core_126 = popcount36_2fox_core_124 ^ popcount36_2fox_core_123;
  assign popcount36_2fox_core_127 = popcount36_2fox_core_124 & popcount36_2fox_core_123;
  assign popcount36_2fox_core_128 = popcount36_2fox_core_125 | popcount36_2fox_core_127;
  assign popcount36_2fox_core_129 = popcount36_2fox_core_075 ^ popcount36_2fox_core_087;
  assign popcount36_2fox_core_130 = popcount36_2fox_core_075 & popcount36_2fox_core_087;
  assign popcount36_2fox_core_131 = popcount36_2fox_core_129 ^ popcount36_2fox_core_128;
  assign popcount36_2fox_core_132 = popcount36_2fox_core_129 & popcount36_2fox_core_128;
  assign popcount36_2fox_core_133 = popcount36_2fox_core_130 | popcount36_2fox_core_132;
  assign popcount36_2fox_core_135 = ~(input_a[11] ^ input_a[23]);
  assign popcount36_2fox_core_136 = popcount36_2fox_core_074 | popcount36_2fox_core_133;
  assign popcount36_2fox_core_139 = input_a[35] | input_a[22];
  assign popcount36_2fox_core_140 = ~(input_a[0] & input_a[10]);
  assign popcount36_2fox_core_142 = input_a[23] ^ input_a[34];
  assign popcount36_2fox_core_143 = input_a[4] & input_a[15];
  assign popcount36_2fox_core_144 = ~(input_a[22] ^ input_a[0]);
  assign popcount36_2fox_core_145 = ~(input_a[23] ^ input_a[29]);
  assign popcount36_2fox_core_147 = ~input_a[3];
  assign popcount36_2fox_core_149 = ~(input_a[13] & input_a[13]);
  assign popcount36_2fox_core_150 = input_a[7] | input_a[26];
  assign popcount36_2fox_core_151 = ~(input_a[11] ^ input_a[32]);
  assign popcount36_2fox_core_152 = ~input_a[1];
  assign popcount36_2fox_core_156 = input_a[20] & input_a[24];
  assign popcount36_2fox_core_157 = input_a[4] ^ input_a[30];
  assign popcount36_2fox_core_158 = input_a[14] & input_a[26];
  assign popcount36_2fox_core_160 = input_a[14] | input_a[21];
  assign popcount36_2fox_core_163 = ~(input_a[6] | input_a[27]);
  assign popcount36_2fox_core_164 = input_a[6] & input_a[18];
  assign popcount36_2fox_core_165 = popcount36_2fox_core_156 ^ popcount36_2fox_core_158;
  assign popcount36_2fox_core_166 = popcount36_2fox_core_156 & popcount36_2fox_core_158;
  assign popcount36_2fox_core_167 = popcount36_2fox_core_165 ^ popcount36_2fox_core_164;
  assign popcount36_2fox_core_168 = popcount36_2fox_core_165 & popcount36_2fox_core_164;
  assign popcount36_2fox_core_169 = popcount36_2fox_core_166 | popcount36_2fox_core_168;
  assign popcount36_2fox_core_172 = ~(input_a[35] | input_a[33]);
  assign popcount36_2fox_core_173 = ~(input_a[31] | input_a[0]);
  assign popcount36_2fox_core_174 = input_a[27] ^ popcount36_2fox_core_167;
  assign popcount36_2fox_core_175 = input_a[27] & popcount36_2fox_core_167;
  assign popcount36_2fox_core_177 = ~(input_a[4] | input_a[8]);
  assign popcount36_2fox_core_179_not = ~popcount36_2fox_core_169;
  assign popcount36_2fox_core_181 = popcount36_2fox_core_179_not ^ popcount36_2fox_core_175;
  assign popcount36_2fox_core_182 = input_a[27] & popcount36_2fox_core_175;
  assign popcount36_2fox_core_183 = popcount36_2fox_core_169 | popcount36_2fox_core_182;
  assign popcount36_2fox_core_185 = ~input_a[14];
  assign popcount36_2fox_core_187 = input_a[15] & input_a[21];
  assign popcount36_2fox_core_188 = input_a[29] ^ input_a[30];
  assign popcount36_2fox_core_189 = input_a[29] & input_a[30];
  assign popcount36_2fox_core_190 = ~(input_a[3] | input_a[17]);
  assign popcount36_2fox_core_191 = input_a[8] & popcount36_2fox_core_188;
  assign popcount36_2fox_core_192 = popcount36_2fox_core_187 ^ popcount36_2fox_core_189;
  assign popcount36_2fox_core_193 = popcount36_2fox_core_187 & popcount36_2fox_core_189;
  assign popcount36_2fox_core_194 = popcount36_2fox_core_192 ^ popcount36_2fox_core_191;
  assign popcount36_2fox_core_195 = popcount36_2fox_core_192 & popcount36_2fox_core_191;
  assign popcount36_2fox_core_196 = popcount36_2fox_core_193 | popcount36_2fox_core_195;
  assign popcount36_2fox_core_197 = input_a[31] ^ input_a[32];
  assign popcount36_2fox_core_198 = input_a[31] & input_a[32];
  assign popcount36_2fox_core_199 = input_a[31] & input_a[17];
  assign popcount36_2fox_core_200 = input_a[19] & input_a[28];
  assign popcount36_2fox_core_201 = ~(input_a[28] ^ input_a[30]);
  assign popcount36_2fox_core_202 = input_a[16] & input_a[34];
  assign popcount36_2fox_core_203 = popcount36_2fox_core_200 | popcount36_2fox_core_202;
  assign popcount36_2fox_core_205 = ~(input_a[1] ^ input_a[14]);
  assign popcount36_2fox_core_206 = popcount36_2fox_core_197 & input_a[13];
  assign popcount36_2fox_core_207 = popcount36_2fox_core_198 ^ popcount36_2fox_core_203;
  assign popcount36_2fox_core_208 = popcount36_2fox_core_198 & popcount36_2fox_core_203;
  assign popcount36_2fox_core_209 = popcount36_2fox_core_207 ^ popcount36_2fox_core_206;
  assign popcount36_2fox_core_210 = popcount36_2fox_core_207 & popcount36_2fox_core_206;
  assign popcount36_2fox_core_211 = popcount36_2fox_core_208 | popcount36_2fox_core_210;
  assign popcount36_2fox_core_216 = popcount36_2fox_core_194 ^ popcount36_2fox_core_209;
  assign popcount36_2fox_core_217 = popcount36_2fox_core_194 & popcount36_2fox_core_209;
  assign popcount36_2fox_core_221 = popcount36_2fox_core_196 ^ popcount36_2fox_core_211;
  assign popcount36_2fox_core_222 = popcount36_2fox_core_196 & popcount36_2fox_core_211;
  assign popcount36_2fox_core_223 = popcount36_2fox_core_221 | popcount36_2fox_core_217;
  assign popcount36_2fox_core_227 = input_a[5] | input_a[6];
  assign popcount36_2fox_core_228 = ~(input_a[13] ^ input_a[25]);
  assign popcount36_2fox_core_230 = popcount36_2fox_core_174 ^ popcount36_2fox_core_216;
  assign popcount36_2fox_core_231 = popcount36_2fox_core_174 & popcount36_2fox_core_216;
  assign popcount36_2fox_core_232 = popcount36_2fox_core_230 ^ input_a[17];
  assign popcount36_2fox_core_233 = popcount36_2fox_core_230 & input_a[17];
  assign popcount36_2fox_core_234 = popcount36_2fox_core_231 | popcount36_2fox_core_233;
  assign popcount36_2fox_core_235 = popcount36_2fox_core_181 ^ popcount36_2fox_core_223;
  assign popcount36_2fox_core_236 = popcount36_2fox_core_181 & popcount36_2fox_core_223;
  assign popcount36_2fox_core_237 = popcount36_2fox_core_235 ^ popcount36_2fox_core_234;
  assign popcount36_2fox_core_238 = popcount36_2fox_core_235 & popcount36_2fox_core_234;
  assign popcount36_2fox_core_239 = popcount36_2fox_core_236 | popcount36_2fox_core_238;
  assign popcount36_2fox_core_240 = popcount36_2fox_core_183 ^ popcount36_2fox_core_222;
  assign popcount36_2fox_core_241 = popcount36_2fox_core_183 & popcount36_2fox_core_222;
  assign popcount36_2fox_core_242 = popcount36_2fox_core_240 ^ popcount36_2fox_core_239;
  assign popcount36_2fox_core_243 = popcount36_2fox_core_240 & popcount36_2fox_core_239;
  assign popcount36_2fox_core_244 = popcount36_2fox_core_241 | popcount36_2fox_core_243;
  assign popcount36_2fox_core_249 = ~(input_a[10] | input_a[0]);
  assign popcount36_2fox_core_251 = input_a[35] & input_a[23];
  assign popcount36_2fox_core_252 = popcount36_2fox_core_126 ^ popcount36_2fox_core_232;
  assign popcount36_2fox_core_253 = popcount36_2fox_core_126 & popcount36_2fox_core_232;
  assign popcount36_2fox_core_254 = popcount36_2fox_core_252 ^ popcount36_2fox_core_251;
  assign popcount36_2fox_core_255 = popcount36_2fox_core_252 & popcount36_2fox_core_251;
  assign popcount36_2fox_core_256 = popcount36_2fox_core_253 | popcount36_2fox_core_255;
  assign popcount36_2fox_core_257 = popcount36_2fox_core_131 ^ popcount36_2fox_core_237;
  assign popcount36_2fox_core_258 = popcount36_2fox_core_131 & popcount36_2fox_core_237;
  assign popcount36_2fox_core_259 = popcount36_2fox_core_257 ^ popcount36_2fox_core_256;
  assign popcount36_2fox_core_260 = popcount36_2fox_core_257 & popcount36_2fox_core_256;
  assign popcount36_2fox_core_261 = popcount36_2fox_core_258 | popcount36_2fox_core_260;
  assign popcount36_2fox_core_262 = popcount36_2fox_core_136 ^ popcount36_2fox_core_242;
  assign popcount36_2fox_core_263 = popcount36_2fox_core_136 & popcount36_2fox_core_242;
  assign popcount36_2fox_core_264 = popcount36_2fox_core_262 ^ popcount36_2fox_core_261;
  assign popcount36_2fox_core_265 = popcount36_2fox_core_262 & popcount36_2fox_core_261;
  assign popcount36_2fox_core_266 = popcount36_2fox_core_263 | popcount36_2fox_core_265;
  assign popcount36_2fox_core_269 = popcount36_2fox_core_244 ^ popcount36_2fox_core_266;
  assign popcount36_2fox_core_270 = popcount36_2fox_core_244 & popcount36_2fox_core_266;
  assign popcount36_2fox_core_272 = ~(input_a[4] | input_a[24]);
  assign popcount36_2fox_core_274 = input_a[17] | input_a[33];
  assign popcount36_2fox_core_275 = ~input_a[6];

  assign popcount36_2fox_out[0] = input_a[25];
  assign popcount36_2fox_out[1] = popcount36_2fox_core_254;
  assign popcount36_2fox_out[2] = popcount36_2fox_core_259;
  assign popcount36_2fox_out[3] = popcount36_2fox_core_264;
  assign popcount36_2fox_out[4] = popcount36_2fox_core_269;
  assign popcount36_2fox_out[5] = popcount36_2fox_core_270;
endmodule