// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.39029
// WCE=9.0
// EP=0.77816%
// Printed PDK parameters:
//  Area=43174938.0
//  Delay=67363560.0
//  Power=2061500.0

module popcount28_n6yf(input [27:0] input_a, output [4:0] popcount28_n6yf_out);
  wire popcount28_n6yf_core_031;
  wire popcount28_n6yf_core_032;
  wire popcount28_n6yf_core_033;
  wire popcount28_n6yf_core_034;
  wire popcount28_n6yf_core_036;
  wire popcount28_n6yf_core_037;
  wire popcount28_n6yf_core_039;
  wire popcount28_n6yf_core_040;
  wire popcount28_n6yf_core_041;
  wire popcount28_n6yf_core_042;
  wire popcount28_n6yf_core_043;
  wire popcount28_n6yf_core_044;
  wire popcount28_n6yf_core_046;
  wire popcount28_n6yf_core_047;
  wire popcount28_n6yf_core_048;
  wire popcount28_n6yf_core_049;
  wire popcount28_n6yf_core_050;
  wire popcount28_n6yf_core_051;
  wire popcount28_n6yf_core_052;
  wire popcount28_n6yf_core_053;
  wire popcount28_n6yf_core_055;
  wire popcount28_n6yf_core_057;
  wire popcount28_n6yf_core_058;
  wire popcount28_n6yf_core_060;
  wire popcount28_n6yf_core_062;
  wire popcount28_n6yf_core_063;
  wire popcount28_n6yf_core_064;
  wire popcount28_n6yf_core_066;
  wire popcount28_n6yf_core_067;
  wire popcount28_n6yf_core_068;
  wire popcount28_n6yf_core_069;
  wire popcount28_n6yf_core_070;
  wire popcount28_n6yf_core_071;
  wire popcount28_n6yf_core_073;
  wire popcount28_n6yf_core_074;
  wire popcount28_n6yf_core_076;
  wire popcount28_n6yf_core_077;
  wire popcount28_n6yf_core_078;
  wire popcount28_n6yf_core_079;
  wire popcount28_n6yf_core_084;
  wire popcount28_n6yf_core_085;
  wire popcount28_n6yf_core_086;
  wire popcount28_n6yf_core_087;
  wire popcount28_n6yf_core_088;
  wire popcount28_n6yf_core_089;
  wire popcount28_n6yf_core_090;
  wire popcount28_n6yf_core_091;
  wire popcount28_n6yf_core_095;
  wire popcount28_n6yf_core_096;
  wire popcount28_n6yf_core_097;
  wire popcount28_n6yf_core_098;
  wire popcount28_n6yf_core_099;
  wire popcount28_n6yf_core_103;
  wire popcount28_n6yf_core_106;
  wire popcount28_n6yf_core_108;
  wire popcount28_n6yf_core_109;
  wire popcount28_n6yf_core_111;
  wire popcount28_n6yf_core_112;
  wire popcount28_n6yf_core_113;
  wire popcount28_n6yf_core_114;
  wire popcount28_n6yf_core_115;
  wire popcount28_n6yf_core_116;
  wire popcount28_n6yf_core_117;
  wire popcount28_n6yf_core_118;
  wire popcount28_n6yf_core_119;
  wire popcount28_n6yf_core_120;
  wire popcount28_n6yf_core_123;
  wire popcount28_n6yf_core_124;
  wire popcount28_n6yf_core_125;
  wire popcount28_n6yf_core_126;
  wire popcount28_n6yf_core_127;
  wire popcount28_n6yf_core_128;
  wire popcount28_n6yf_core_130;
  wire popcount28_n6yf_core_131;
  wire popcount28_n6yf_core_132_not;
  wire popcount28_n6yf_core_133;
  wire popcount28_n6yf_core_135;
  wire popcount28_n6yf_core_136;
  wire popcount28_n6yf_core_137;
  wire popcount28_n6yf_core_139;
  wire popcount28_n6yf_core_140;
  wire popcount28_n6yf_core_143;
  wire popcount28_n6yf_core_144;
  wire popcount28_n6yf_core_146;
  wire popcount28_n6yf_core_147;
  wire popcount28_n6yf_core_148;
  wire popcount28_n6yf_core_149;
  wire popcount28_n6yf_core_150;
  wire popcount28_n6yf_core_152;
  wire popcount28_n6yf_core_155;
  wire popcount28_n6yf_core_156;
  wire popcount28_n6yf_core_162;
  wire popcount28_n6yf_core_163;
  wire popcount28_n6yf_core_164;
  wire popcount28_n6yf_core_165;
  wire popcount28_n6yf_core_166;
  wire popcount28_n6yf_core_167;
  wire popcount28_n6yf_core_168;
  wire popcount28_n6yf_core_169;
  wire popcount28_n6yf_core_170;
  wire popcount28_n6yf_core_171;
  wire popcount28_n6yf_core_172;
  wire popcount28_n6yf_core_173;
  wire popcount28_n6yf_core_174;
  wire popcount28_n6yf_core_176;
  wire popcount28_n6yf_core_178;
  wire popcount28_n6yf_core_179;
  wire popcount28_n6yf_core_180;
  wire popcount28_n6yf_core_182;
  wire popcount28_n6yf_core_183;
  wire popcount28_n6yf_core_184;
  wire popcount28_n6yf_core_185;
  wire popcount28_n6yf_core_186;
  wire popcount28_n6yf_core_187;
  wire popcount28_n6yf_core_188;
  wire popcount28_n6yf_core_189;
  wire popcount28_n6yf_core_190;
  wire popcount28_n6yf_core_191;
  wire popcount28_n6yf_core_192;
  wire popcount28_n6yf_core_193;
  wire popcount28_n6yf_core_194;
  wire popcount28_n6yf_core_195;
  wire popcount28_n6yf_core_196;
  wire popcount28_n6yf_core_197_not;
  wire popcount28_n6yf_core_199;
  wire popcount28_n6yf_core_201;

  assign popcount28_n6yf_core_031 = input_a[23] & input_a[24];
  assign popcount28_n6yf_core_032 = ~(input_a[21] | input_a[6]);
  assign popcount28_n6yf_core_033 = input_a[12] ^ input_a[2];
  assign popcount28_n6yf_core_034 = popcount28_n6yf_core_031 | input_a[13];
  assign popcount28_n6yf_core_036 = input_a[3] | input_a[4];
  assign popcount28_n6yf_core_037 = input_a[3] & input_a[4];
  assign popcount28_n6yf_core_039 = input_a[5] & input_a[6];
  assign popcount28_n6yf_core_040 = ~(input_a[22] & input_a[7]);
  assign popcount28_n6yf_core_041 = popcount28_n6yf_core_036 & input_a[8];
  assign popcount28_n6yf_core_042 = popcount28_n6yf_core_037 | popcount28_n6yf_core_039;
  assign popcount28_n6yf_core_043 = ~(input_a[19] ^ input_a[11]);
  assign popcount28_n6yf_core_044 = popcount28_n6yf_core_042 | popcount28_n6yf_core_041;
  assign popcount28_n6yf_core_046 = ~(input_a[9] & input_a[14]);
  assign popcount28_n6yf_core_047 = ~(input_a[10] | input_a[0]);
  assign popcount28_n6yf_core_048 = input_a[25] & input_a[0];
  assign popcount28_n6yf_core_049 = popcount28_n6yf_core_034 ^ popcount28_n6yf_core_044;
  assign popcount28_n6yf_core_050 = popcount28_n6yf_core_034 & popcount28_n6yf_core_044;
  assign popcount28_n6yf_core_051 = popcount28_n6yf_core_049 ^ popcount28_n6yf_core_048;
  assign popcount28_n6yf_core_052 = popcount28_n6yf_core_049 & popcount28_n6yf_core_048;
  assign popcount28_n6yf_core_053 = popcount28_n6yf_core_050 | popcount28_n6yf_core_052;
  assign popcount28_n6yf_core_055 = input_a[14] ^ input_a[11];
  assign popcount28_n6yf_core_057 = input_a[14] & input_a[23];
  assign popcount28_n6yf_core_058 = ~(input_a[21] ^ input_a[12]);
  assign popcount28_n6yf_core_060 = input_a[9] & input_a[19];
  assign popcount28_n6yf_core_062 = ~(input_a[15] | input_a[27]);
  assign popcount28_n6yf_core_063 = input_a[21] ^ input_a[7];
  assign popcount28_n6yf_core_064 = ~(input_a[12] ^ input_a[6]);
  assign popcount28_n6yf_core_066 = input_a[24] & input_a[1];
  assign popcount28_n6yf_core_067 = ~input_a[26];
  assign popcount28_n6yf_core_068 = input_a[15] ^ input_a[27];
  assign popcount28_n6yf_core_069 = input_a[2] & input_a[5];
  assign popcount28_n6yf_core_070 = input_a[0] ^ input_a[27];
  assign popcount28_n6yf_core_071 = ~(input_a[19] & input_a[5]);
  assign popcount28_n6yf_core_073 = input_a[7] | input_a[18];
  assign popcount28_n6yf_core_074 = input_a[1] | input_a[20];
  assign popcount28_n6yf_core_076 = ~input_a[22];
  assign popcount28_n6yf_core_077 = input_a[12] ^ input_a[13];
  assign popcount28_n6yf_core_078 = ~(popcount28_n6yf_core_063 & popcount28_n6yf_core_073);
  assign popcount28_n6yf_core_079 = input_a[21] & input_a[18];
  assign popcount28_n6yf_core_084 = input_a[9] | input_a[20];
  assign popcount28_n6yf_core_085 = input_a[7] | popcount28_n6yf_core_079;
  assign popcount28_n6yf_core_086 = ~input_a[23];
  assign popcount28_n6yf_core_087 = ~(input_a[6] ^ input_a[15]);
  assign popcount28_n6yf_core_088 = ~input_a[7];
  assign popcount28_n6yf_core_089 = ~(input_a[16] ^ input_a[14]);
  assign popcount28_n6yf_core_090 = popcount28_n6yf_core_051 ^ popcount28_n6yf_core_078;
  assign popcount28_n6yf_core_091 = popcount28_n6yf_core_051 & popcount28_n6yf_core_078;
  assign popcount28_n6yf_core_095 = popcount28_n6yf_core_053 ^ popcount28_n6yf_core_085;
  assign popcount28_n6yf_core_096 = popcount28_n6yf_core_053 & popcount28_n6yf_core_085;
  assign popcount28_n6yf_core_097 = popcount28_n6yf_core_095 ^ popcount28_n6yf_core_091;
  assign popcount28_n6yf_core_098 = popcount28_n6yf_core_095 & popcount28_n6yf_core_091;
  assign popcount28_n6yf_core_099 = popcount28_n6yf_core_096 | popcount28_n6yf_core_098;
  assign popcount28_n6yf_core_103 = ~input_a[1];
  assign popcount28_n6yf_core_106 = input_a[22] & input_a[11];
  assign popcount28_n6yf_core_108 = input_a[1] & input_a[9];
  assign popcount28_n6yf_core_109 = popcount28_n6yf_core_106 | popcount28_n6yf_core_108;
  assign popcount28_n6yf_core_111 = ~(input_a[18] ^ input_a[26]);
  assign popcount28_n6yf_core_112 = input_a[16] & input_a[27];
  assign popcount28_n6yf_core_113 = input_a[19] | input_a[20];
  assign popcount28_n6yf_core_114 = input_a[19] & input_a[20];
  assign popcount28_n6yf_core_115 = ~(input_a[1] & input_a[11]);
  assign popcount28_n6yf_core_116 = input_a[10] & popcount28_n6yf_core_113;
  assign popcount28_n6yf_core_117 = popcount28_n6yf_core_112 ^ popcount28_n6yf_core_114;
  assign popcount28_n6yf_core_118 = popcount28_n6yf_core_112 & popcount28_n6yf_core_114;
  assign popcount28_n6yf_core_119 = popcount28_n6yf_core_117 | popcount28_n6yf_core_116;
  assign popcount28_n6yf_core_120 = ~(input_a[17] ^ input_a[19]);
  assign popcount28_n6yf_core_123 = input_a[12] & input_a[2];
  assign popcount28_n6yf_core_124 = popcount28_n6yf_core_109 ^ popcount28_n6yf_core_119;
  assign popcount28_n6yf_core_125 = popcount28_n6yf_core_109 & popcount28_n6yf_core_119;
  assign popcount28_n6yf_core_126 = popcount28_n6yf_core_124 ^ popcount28_n6yf_core_123;
  assign popcount28_n6yf_core_127 = popcount28_n6yf_core_124 & popcount28_n6yf_core_123;
  assign popcount28_n6yf_core_128 = popcount28_n6yf_core_125 | popcount28_n6yf_core_127;
  assign popcount28_n6yf_core_130 = ~input_a[20];
  assign popcount28_n6yf_core_131 = popcount28_n6yf_core_118 | popcount28_n6yf_core_128;
  assign popcount28_n6yf_core_132_not = ~input_a[10];
  assign popcount28_n6yf_core_133 = ~input_a[5];
  assign popcount28_n6yf_core_135 = ~input_a[19];
  assign popcount28_n6yf_core_136 = input_a[2] | input_a[24];
  assign popcount28_n6yf_core_137 = ~(input_a[16] ^ input_a[9]);
  assign popcount28_n6yf_core_139 = ~(input_a[11] | input_a[11]);
  assign popcount28_n6yf_core_140 = ~(input_a[14] & input_a[26]);
  assign popcount28_n6yf_core_143 = ~(input_a[13] & input_a[9]);
  assign popcount28_n6yf_core_144 = ~(input_a[14] ^ input_a[22]);
  assign popcount28_n6yf_core_146 = input_a[9] ^ input_a[16];
  assign popcount28_n6yf_core_147 = input_a[2] | input_a[11];
  assign popcount28_n6yf_core_148 = input_a[20] | input_a[7];
  assign popcount28_n6yf_core_149 = input_a[13] & input_a[15];
  assign popcount28_n6yf_core_150 = ~(input_a[4] & input_a[3]);
  assign popcount28_n6yf_core_152 = ~(input_a[5] | input_a[27]);
  assign popcount28_n6yf_core_155 = ~(input_a[17] & input_a[26]);
  assign popcount28_n6yf_core_156 = input_a[17] & input_a[26];
  assign popcount28_n6yf_core_162 = ~(input_a[19] & input_a[3]);
  assign popcount28_n6yf_core_163 = ~input_a[5];
  assign popcount28_n6yf_core_164 = input_a[15] & input_a[14];
  assign popcount28_n6yf_core_165 = popcount28_n6yf_core_126 ^ popcount28_n6yf_core_155;
  assign popcount28_n6yf_core_166 = popcount28_n6yf_core_126 & popcount28_n6yf_core_155;
  assign popcount28_n6yf_core_167 = popcount28_n6yf_core_165 ^ popcount28_n6yf_core_164;
  assign popcount28_n6yf_core_168 = popcount28_n6yf_core_165 & popcount28_n6yf_core_164;
  assign popcount28_n6yf_core_169 = popcount28_n6yf_core_166 | popcount28_n6yf_core_168;
  assign popcount28_n6yf_core_170 = popcount28_n6yf_core_131 ^ popcount28_n6yf_core_156;
  assign popcount28_n6yf_core_171 = popcount28_n6yf_core_131 & popcount28_n6yf_core_156;
  assign popcount28_n6yf_core_172 = popcount28_n6yf_core_170 ^ popcount28_n6yf_core_169;
  assign popcount28_n6yf_core_173 = popcount28_n6yf_core_170 & popcount28_n6yf_core_169;
  assign popcount28_n6yf_core_174 = popcount28_n6yf_core_171 | popcount28_n6yf_core_173;
  assign popcount28_n6yf_core_176 = ~(input_a[9] & input_a[4]);
  assign popcount28_n6yf_core_178 = ~(input_a[21] & input_a[2]);
  assign popcount28_n6yf_core_179 = ~(input_a[26] | input_a[16]);
  assign popcount28_n6yf_core_180 = ~input_a[16];
  assign popcount28_n6yf_core_182 = popcount28_n6yf_core_090 ^ popcount28_n6yf_core_167;
  assign popcount28_n6yf_core_183 = popcount28_n6yf_core_090 & popcount28_n6yf_core_167;
  assign popcount28_n6yf_core_184 = popcount28_n6yf_core_182 ^ popcount28_n6yf_core_088;
  assign popcount28_n6yf_core_185 = popcount28_n6yf_core_182 & popcount28_n6yf_core_088;
  assign popcount28_n6yf_core_186 = popcount28_n6yf_core_183 | popcount28_n6yf_core_185;
  assign popcount28_n6yf_core_187 = popcount28_n6yf_core_097 ^ popcount28_n6yf_core_172;
  assign popcount28_n6yf_core_188 = popcount28_n6yf_core_097 & popcount28_n6yf_core_172;
  assign popcount28_n6yf_core_189 = popcount28_n6yf_core_187 ^ popcount28_n6yf_core_186;
  assign popcount28_n6yf_core_190 = popcount28_n6yf_core_187 & popcount28_n6yf_core_186;
  assign popcount28_n6yf_core_191 = popcount28_n6yf_core_188 | popcount28_n6yf_core_190;
  assign popcount28_n6yf_core_192 = popcount28_n6yf_core_099 ^ popcount28_n6yf_core_174;
  assign popcount28_n6yf_core_193 = popcount28_n6yf_core_099 & popcount28_n6yf_core_174;
  assign popcount28_n6yf_core_194 = popcount28_n6yf_core_192 ^ popcount28_n6yf_core_191;
  assign popcount28_n6yf_core_195 = popcount28_n6yf_core_192 & popcount28_n6yf_core_191;
  assign popcount28_n6yf_core_196 = popcount28_n6yf_core_193 | popcount28_n6yf_core_195;
  assign popcount28_n6yf_core_197_not = ~input_a[9];
  assign popcount28_n6yf_core_199 = input_a[5] & input_a[12];
  assign popcount28_n6yf_core_201 = ~(input_a[20] ^ input_a[15]);

  assign popcount28_n6yf_out[0] = popcount28_n6yf_core_194;
  assign popcount28_n6yf_out[1] = popcount28_n6yf_core_184;
  assign popcount28_n6yf_out[2] = popcount28_n6yf_core_189;
  assign popcount28_n6yf_out[3] = popcount28_n6yf_core_194;
  assign popcount28_n6yf_out[4] = popcount28_n6yf_core_196;
endmodule