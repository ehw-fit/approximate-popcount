// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.51395
// WCE=6.0
// EP=0.800797%
// Printed PDK parameters:
//  Area=54066298.0
//  Delay=70794392.0
//  Power=2896400.0

module popcount29_7rcu(input [28:0] input_a, output [4:0] popcount29_7rcu_out);
  wire popcount29_7rcu_core_031;
  wire popcount29_7rcu_core_032;
  wire popcount29_7rcu_core_033;
  wire popcount29_7rcu_core_034;
  wire popcount29_7rcu_core_035;
  wire popcount29_7rcu_core_037;
  wire popcount29_7rcu_core_038;
  wire popcount29_7rcu_core_039;
  wire popcount29_7rcu_core_040;
  wire popcount29_7rcu_core_041;
  wire popcount29_7rcu_core_042;
  wire popcount29_7rcu_core_043;
  wire popcount29_7rcu_core_044;
  wire popcount29_7rcu_core_045;
  wire popcount29_7rcu_core_046;
  wire popcount29_7rcu_core_049;
  wire popcount29_7rcu_core_050;
  wire popcount29_7rcu_core_051;
  wire popcount29_7rcu_core_053;
  wire popcount29_7rcu_core_054;
  wire popcount29_7rcu_core_057;
  wire popcount29_7rcu_core_058;
  wire popcount29_7rcu_core_061;
  wire popcount29_7rcu_core_062;
  wire popcount29_7rcu_core_063;
  wire popcount29_7rcu_core_064;
  wire popcount29_7rcu_core_066;
  wire popcount29_7rcu_core_067;
  wire popcount29_7rcu_core_068;
  wire popcount29_7rcu_core_069;
  wire popcount29_7rcu_core_070;
  wire popcount29_7rcu_core_071;
  wire popcount29_7rcu_core_072;
  wire popcount29_7rcu_core_073;
  wire popcount29_7rcu_core_075;
  wire popcount29_7rcu_core_078;
  wire popcount29_7rcu_core_079;
  wire popcount29_7rcu_core_080;
  wire popcount29_7rcu_core_082;
  wire popcount29_7rcu_core_086;
  wire popcount29_7rcu_core_088;
  wire popcount29_7rcu_core_089;
  wire popcount29_7rcu_core_090;
  wire popcount29_7rcu_core_093;
  wire popcount29_7rcu_core_094;
  wire popcount29_7rcu_core_096;
  wire popcount29_7rcu_core_097;
  wire popcount29_7rcu_core_098;
  wire popcount29_7rcu_core_099;
  wire popcount29_7rcu_core_100;
  wire popcount29_7rcu_core_102;
  wire popcount29_7rcu_core_104;
  wire popcount29_7rcu_core_108;
  wire popcount29_7rcu_core_112;
  wire popcount29_7rcu_core_113;
  wire popcount29_7rcu_core_114;
  wire popcount29_7rcu_core_115;
  wire popcount29_7rcu_core_116;
  wire popcount29_7rcu_core_117;
  wire popcount29_7rcu_core_118;
  wire popcount29_7rcu_core_119;
  wire popcount29_7rcu_core_120;
  wire popcount29_7rcu_core_122;
  wire popcount29_7rcu_core_123;
  wire popcount29_7rcu_core_125;
  wire popcount29_7rcu_core_126;
  wire popcount29_7rcu_core_127;
  wire popcount29_7rcu_core_131;
  wire popcount29_7rcu_core_132;
  wire popcount29_7rcu_core_133;
  wire popcount29_7rcu_core_135;
  wire popcount29_7rcu_core_136;
  wire popcount29_7rcu_core_137;
  wire popcount29_7rcu_core_138;
  wire popcount29_7rcu_core_139;
  wire popcount29_7rcu_core_140;
  wire popcount29_7rcu_core_141;
  wire popcount29_7rcu_core_142;
  wire popcount29_7rcu_core_143;
  wire popcount29_7rcu_core_146;
  wire popcount29_7rcu_core_149;
  wire popcount29_7rcu_core_150;
  wire popcount29_7rcu_core_151;
  wire popcount29_7rcu_core_152;
  wire popcount29_7rcu_core_153;
  wire popcount29_7rcu_core_154;
  wire popcount29_7rcu_core_156;
  wire popcount29_7rcu_core_157;
  wire popcount29_7rcu_core_158;
  wire popcount29_7rcu_core_159;
  wire popcount29_7rcu_core_160;
  wire popcount29_7rcu_core_161;
  wire popcount29_7rcu_core_162;
  wire popcount29_7rcu_core_163;
  wire popcount29_7rcu_core_164;
  wire popcount29_7rcu_core_166;
  wire popcount29_7rcu_core_167;
  wire popcount29_7rcu_core_168;
  wire popcount29_7rcu_core_169;
  wire popcount29_7rcu_core_170;
  wire popcount29_7rcu_core_171;
  wire popcount29_7rcu_core_172;
  wire popcount29_7rcu_core_174;
  wire popcount29_7rcu_core_176;
  wire popcount29_7rcu_core_177;
  wire popcount29_7rcu_core_178;
  wire popcount29_7rcu_core_179;
  wire popcount29_7rcu_core_180;
  wire popcount29_7rcu_core_183;
  wire popcount29_7rcu_core_185;
  wire popcount29_7rcu_core_186;
  wire popcount29_7rcu_core_187;
  wire popcount29_7rcu_core_188;
  wire popcount29_7rcu_core_189;
  wire popcount29_7rcu_core_190;
  wire popcount29_7rcu_core_191;
  wire popcount29_7rcu_core_192;
  wire popcount29_7rcu_core_193;
  wire popcount29_7rcu_core_194;
  wire popcount29_7rcu_core_195;
  wire popcount29_7rcu_core_196;
  wire popcount29_7rcu_core_197;
  wire popcount29_7rcu_core_198;
  wire popcount29_7rcu_core_199;
  wire popcount29_7rcu_core_200;
  wire popcount29_7rcu_core_201;
  wire popcount29_7rcu_core_202;
  wire popcount29_7rcu_core_203;
  wire popcount29_7rcu_core_205;

  assign popcount29_7rcu_core_031 = input_a[1] ^ input_a[2];
  assign popcount29_7rcu_core_032 = input_a[1] & input_a[2];
  assign popcount29_7rcu_core_033 = input_a[0] ^ popcount29_7rcu_core_031;
  assign popcount29_7rcu_core_034 = input_a[0] & popcount29_7rcu_core_031;
  assign popcount29_7rcu_core_035 = popcount29_7rcu_core_032 | popcount29_7rcu_core_034;
  assign popcount29_7rcu_core_037 = input_a[3] ^ input_a[4];
  assign popcount29_7rcu_core_038 = input_a[3] & input_a[4];
  assign popcount29_7rcu_core_039 = input_a[5] ^ input_a[6];
  assign popcount29_7rcu_core_040 = input_a[5] & input_a[6];
  assign popcount29_7rcu_core_041 = popcount29_7rcu_core_037 ^ popcount29_7rcu_core_039;
  assign popcount29_7rcu_core_042 = popcount29_7rcu_core_037 & popcount29_7rcu_core_039;
  assign popcount29_7rcu_core_043 = popcount29_7rcu_core_038 | popcount29_7rcu_core_040;
  assign popcount29_7rcu_core_044 = popcount29_7rcu_core_038 & popcount29_7rcu_core_040;
  assign popcount29_7rcu_core_045 = popcount29_7rcu_core_043 | popcount29_7rcu_core_042;
  assign popcount29_7rcu_core_046 = ~(input_a[4] ^ input_a[27]);
  assign popcount29_7rcu_core_049 = popcount29_7rcu_core_033 & popcount29_7rcu_core_041;
  assign popcount29_7rcu_core_050 = popcount29_7rcu_core_035 | popcount29_7rcu_core_045;
  assign popcount29_7rcu_core_051 = popcount29_7rcu_core_035 & popcount29_7rcu_core_045;
  assign popcount29_7rcu_core_053 = popcount29_7rcu_core_050 & popcount29_7rcu_core_049;
  assign popcount29_7rcu_core_054 = popcount29_7rcu_core_051 | popcount29_7rcu_core_053;
  assign popcount29_7rcu_core_057 = popcount29_7rcu_core_044 | popcount29_7rcu_core_054;
  assign popcount29_7rcu_core_058 = ~(input_a[17] | input_a[18]);
  assign popcount29_7rcu_core_061 = input_a[8] & input_a[9];
  assign popcount29_7rcu_core_062 = input_a[28] & input_a[18];
  assign popcount29_7rcu_core_063 = input_a[13] & input_a[11];
  assign popcount29_7rcu_core_064 = popcount29_7rcu_core_061 | popcount29_7rcu_core_063;
  assign popcount29_7rcu_core_066 = input_a[19] | input_a[26];
  assign popcount29_7rcu_core_067 = input_a[10] & input_a[27];
  assign popcount29_7rcu_core_068 = ~(input_a[22] ^ input_a[8]);
  assign popcount29_7rcu_core_069 = input_a[16] & input_a[15];
  assign popcount29_7rcu_core_070 = input_a[20] | input_a[17];
  assign popcount29_7rcu_core_071 = ~(input_a[2] & input_a[25]);
  assign popcount29_7rcu_core_072 = popcount29_7rcu_core_067 ^ popcount29_7rcu_core_069;
  assign popcount29_7rcu_core_073 = popcount29_7rcu_core_067 & popcount29_7rcu_core_069;
  assign popcount29_7rcu_core_075 = ~(input_a[20] ^ input_a[25]);
  assign popcount29_7rcu_core_078 = ~(input_a[10] | input_a[13]);
  assign popcount29_7rcu_core_079 = popcount29_7rcu_core_064 ^ popcount29_7rcu_core_072;
  assign popcount29_7rcu_core_080 = popcount29_7rcu_core_064 & popcount29_7rcu_core_072;
  assign popcount29_7rcu_core_082 = ~(input_a[21] | input_a[2]);
  assign popcount29_7rcu_core_086 = popcount29_7rcu_core_073 | popcount29_7rcu_core_080;
  assign popcount29_7rcu_core_088 = input_a[11] | input_a[17];
  assign popcount29_7rcu_core_089 = ~(input_a[23] ^ input_a[14]);
  assign popcount29_7rcu_core_090 = ~input_a[18];
  assign popcount29_7rcu_core_093 = popcount29_7rcu_core_079 ^ input_a[26];
  assign popcount29_7rcu_core_094 = popcount29_7rcu_core_079 & input_a[26];
  assign popcount29_7rcu_core_096 = popcount29_7rcu_core_057 ^ popcount29_7rcu_core_086;
  assign popcount29_7rcu_core_097 = popcount29_7rcu_core_057 & popcount29_7rcu_core_086;
  assign popcount29_7rcu_core_098 = popcount29_7rcu_core_096 ^ popcount29_7rcu_core_094;
  assign popcount29_7rcu_core_099 = popcount29_7rcu_core_096 & popcount29_7rcu_core_094;
  assign popcount29_7rcu_core_100 = popcount29_7rcu_core_097 | popcount29_7rcu_core_099;
  assign popcount29_7rcu_core_102 = ~input_a[7];
  assign popcount29_7rcu_core_104 = ~input_a[21];
  assign popcount29_7rcu_core_108 = ~input_a[14];
  assign popcount29_7rcu_core_112 = input_a[16] ^ input_a[11];
  assign popcount29_7rcu_core_113 = input_a[17] & input_a[18];
  assign popcount29_7rcu_core_114 = input_a[19] ^ input_a[20];
  assign popcount29_7rcu_core_115 = input_a[19] & input_a[20];
  assign popcount29_7rcu_core_116 = ~input_a[0];
  assign popcount29_7rcu_core_117 = input_a[14] & popcount29_7rcu_core_114;
  assign popcount29_7rcu_core_118 = popcount29_7rcu_core_113 ^ popcount29_7rcu_core_115;
  assign popcount29_7rcu_core_119 = input_a[17] & input_a[18];
  assign popcount29_7rcu_core_120 = popcount29_7rcu_core_118 | popcount29_7rcu_core_117;
  assign popcount29_7rcu_core_122 = popcount29_7rcu_core_119 | popcount29_7rcu_core_118;
  assign popcount29_7rcu_core_123 = ~(input_a[17] ^ input_a[10]);
  assign popcount29_7rcu_core_125 = input_a[14] ^ popcount29_7rcu_core_120;
  assign popcount29_7rcu_core_126 = input_a[14] & popcount29_7rcu_core_120;
  assign popcount29_7rcu_core_127 = popcount29_7rcu_core_125 ^ popcount29_7rcu_core_108;
  assign popcount29_7rcu_core_131 = ~(input_a[26] | input_a[11]);
  assign popcount29_7rcu_core_132 = popcount29_7rcu_core_122 | popcount29_7rcu_core_126;
  assign popcount29_7rcu_core_133 = ~(input_a[12] | input_a[2]);
  assign popcount29_7rcu_core_135 = input_a[21] ^ input_a[22];
  assign popcount29_7rcu_core_136 = input_a[21] & input_a[22];
  assign popcount29_7rcu_core_137 = input_a[23] ^ input_a[24];
  assign popcount29_7rcu_core_138 = input_a[23] & input_a[24];
  assign popcount29_7rcu_core_139 = popcount29_7rcu_core_135 ^ popcount29_7rcu_core_137;
  assign popcount29_7rcu_core_140 = popcount29_7rcu_core_135 & popcount29_7rcu_core_137;
  assign popcount29_7rcu_core_141 = popcount29_7rcu_core_136 ^ popcount29_7rcu_core_138;
  assign popcount29_7rcu_core_142 = popcount29_7rcu_core_136 & popcount29_7rcu_core_138;
  assign popcount29_7rcu_core_143 = popcount29_7rcu_core_141 | popcount29_7rcu_core_140;
  assign popcount29_7rcu_core_146 = ~(input_a[8] | input_a[15]);
  assign popcount29_7rcu_core_149 = input_a[15] | input_a[16];
  assign popcount29_7rcu_core_150 = input_a[22] & input_a[19];
  assign popcount29_7rcu_core_151 = ~(input_a[22] ^ input_a[19]);
  assign popcount29_7rcu_core_152 = ~(input_a[22] & input_a[25]);
  assign popcount29_7rcu_core_153 = ~(input_a[13] ^ input_a[9]);
  assign popcount29_7rcu_core_154 = ~input_a[25];
  assign popcount29_7rcu_core_156 = ~(input_a[12] | input_a[21]);
  assign popcount29_7rcu_core_157 = ~(input_a[12] ^ input_a[18]);
  assign popcount29_7rcu_core_158 = popcount29_7rcu_core_139 & input_a[7];
  assign popcount29_7rcu_core_159 = popcount29_7rcu_core_143 ^ popcount29_7rcu_core_154;
  assign popcount29_7rcu_core_160 = popcount29_7rcu_core_143 & popcount29_7rcu_core_154;
  assign popcount29_7rcu_core_161 = popcount29_7rcu_core_159 ^ popcount29_7rcu_core_158;
  assign popcount29_7rcu_core_162 = popcount29_7rcu_core_159 & popcount29_7rcu_core_158;
  assign popcount29_7rcu_core_163 = popcount29_7rcu_core_160 | popcount29_7rcu_core_162;
  assign popcount29_7rcu_core_164 = popcount29_7rcu_core_142 ^ input_a[25];
  assign popcount29_7rcu_core_166 = popcount29_7rcu_core_164 ^ popcount29_7rcu_core_163;
  assign popcount29_7rcu_core_167 = input_a[25] & popcount29_7rcu_core_163;
  assign popcount29_7rcu_core_168 = popcount29_7rcu_core_142 | popcount29_7rcu_core_167;
  assign popcount29_7rcu_core_169 = ~(input_a[24] & input_a[9]);
  assign popcount29_7rcu_core_170 = ~(input_a[4] | input_a[22]);
  assign popcount29_7rcu_core_171 = popcount29_7rcu_core_127 ^ popcount29_7rcu_core_161;
  assign popcount29_7rcu_core_172 = popcount29_7rcu_core_127 & popcount29_7rcu_core_161;
  assign popcount29_7rcu_core_174 = ~(input_a[20] ^ input_a[24]);
  assign popcount29_7rcu_core_176 = popcount29_7rcu_core_132 ^ popcount29_7rcu_core_166;
  assign popcount29_7rcu_core_177 = popcount29_7rcu_core_132 & popcount29_7rcu_core_166;
  assign popcount29_7rcu_core_178 = popcount29_7rcu_core_176 ^ popcount29_7rcu_core_172;
  assign popcount29_7rcu_core_179 = popcount29_7rcu_core_176 & popcount29_7rcu_core_172;
  assign popcount29_7rcu_core_180 = popcount29_7rcu_core_177 | popcount29_7rcu_core_179;
  assign popcount29_7rcu_core_183 = popcount29_7rcu_core_168 | popcount29_7rcu_core_180;
  assign popcount29_7rcu_core_185 = ~(input_a[3] & input_a[1]);
  assign popcount29_7rcu_core_186 = input_a[9] ^ input_a[25];
  assign popcount29_7rcu_core_187 = input_a[12] & input_a[28];
  assign popcount29_7rcu_core_188 = popcount29_7rcu_core_093 ^ popcount29_7rcu_core_171;
  assign popcount29_7rcu_core_189 = popcount29_7rcu_core_093 & popcount29_7rcu_core_171;
  assign popcount29_7rcu_core_190 = popcount29_7rcu_core_188 ^ popcount29_7rcu_core_187;
  assign popcount29_7rcu_core_191 = popcount29_7rcu_core_188 & popcount29_7rcu_core_187;
  assign popcount29_7rcu_core_192 = popcount29_7rcu_core_189 | popcount29_7rcu_core_191;
  assign popcount29_7rcu_core_193 = popcount29_7rcu_core_098 ^ popcount29_7rcu_core_178;
  assign popcount29_7rcu_core_194 = popcount29_7rcu_core_098 & popcount29_7rcu_core_178;
  assign popcount29_7rcu_core_195 = popcount29_7rcu_core_193 ^ popcount29_7rcu_core_192;
  assign popcount29_7rcu_core_196 = popcount29_7rcu_core_193 & popcount29_7rcu_core_192;
  assign popcount29_7rcu_core_197 = popcount29_7rcu_core_194 | popcount29_7rcu_core_196;
  assign popcount29_7rcu_core_198 = popcount29_7rcu_core_100 ^ popcount29_7rcu_core_183;
  assign popcount29_7rcu_core_199 = popcount29_7rcu_core_100 & popcount29_7rcu_core_183;
  assign popcount29_7rcu_core_200 = popcount29_7rcu_core_198 ^ popcount29_7rcu_core_197;
  assign popcount29_7rcu_core_201 = popcount29_7rcu_core_198 & popcount29_7rcu_core_197;
  assign popcount29_7rcu_core_202 = popcount29_7rcu_core_199 | popcount29_7rcu_core_201;
  assign popcount29_7rcu_core_203 = input_a[22] | input_a[23];
  assign popcount29_7rcu_core_205 = input_a[10] ^ input_a[19];

  assign popcount29_7rcu_out[0] = popcount29_7rcu_core_154;
  assign popcount29_7rcu_out[1] = popcount29_7rcu_core_190;
  assign popcount29_7rcu_out[2] = popcount29_7rcu_core_195;
  assign popcount29_7rcu_out[3] = popcount29_7rcu_core_200;
  assign popcount29_7rcu_out[4] = popcount29_7rcu_core_202;
endmodule