// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.69524
// WCE=19.0
// EP=0.884291%
// Printed PDK parameters:
//  Area=2151060.0
//  Delay=6783958.5
//  Power=116290.0

module popcount38_2oru(input [37:0] input_a, output [5:0] popcount38_2oru_out);
  wire popcount38_2oru_core_040;
  wire popcount38_2oru_core_041;
  wire popcount38_2oru_core_042;
  wire popcount38_2oru_core_043;
  wire popcount38_2oru_core_044;
  wire popcount38_2oru_core_045;
  wire popcount38_2oru_core_046;
  wire popcount38_2oru_core_048;
  wire popcount38_2oru_core_050;
  wire popcount38_2oru_core_051;
  wire popcount38_2oru_core_052;
  wire popcount38_2oru_core_053_not;
  wire popcount38_2oru_core_054;
  wire popcount38_2oru_core_055;
  wire popcount38_2oru_core_056;
  wire popcount38_2oru_core_057;
  wire popcount38_2oru_core_059;
  wire popcount38_2oru_core_060;
  wire popcount38_2oru_core_061;
  wire popcount38_2oru_core_066;
  wire popcount38_2oru_core_067;
  wire popcount38_2oru_core_068;
  wire popcount38_2oru_core_072;
  wire popcount38_2oru_core_073;
  wire popcount38_2oru_core_076;
  wire popcount38_2oru_core_077;
  wire popcount38_2oru_core_078;
  wire popcount38_2oru_core_079;
  wire popcount38_2oru_core_080;
  wire popcount38_2oru_core_082;
  wire popcount38_2oru_core_084;
  wire popcount38_2oru_core_085;
  wire popcount38_2oru_core_086;
  wire popcount38_2oru_core_087;
  wire popcount38_2oru_core_088;
  wire popcount38_2oru_core_090;
  wire popcount38_2oru_core_093;
  wire popcount38_2oru_core_094;
  wire popcount38_2oru_core_095;
  wire popcount38_2oru_core_096;
  wire popcount38_2oru_core_097;
  wire popcount38_2oru_core_098;
  wire popcount38_2oru_core_102;
  wire popcount38_2oru_core_103_not;
  wire popcount38_2oru_core_104;
  wire popcount38_2oru_core_105;
  wire popcount38_2oru_core_106;
  wire popcount38_2oru_core_110;
  wire popcount38_2oru_core_111;
  wire popcount38_2oru_core_113;
  wire popcount38_2oru_core_114;
  wire popcount38_2oru_core_115;
  wire popcount38_2oru_core_116;
  wire popcount38_2oru_core_121;
  wire popcount38_2oru_core_122;
  wire popcount38_2oru_core_124;
  wire popcount38_2oru_core_126;
  wire popcount38_2oru_core_128;
  wire popcount38_2oru_core_129;
  wire popcount38_2oru_core_131;
  wire popcount38_2oru_core_132;
  wire popcount38_2oru_core_137;
  wire popcount38_2oru_core_138;
  wire popcount38_2oru_core_139;
  wire popcount38_2oru_core_141;
  wire popcount38_2oru_core_142;
  wire popcount38_2oru_core_143;
  wire popcount38_2oru_core_151;
  wire popcount38_2oru_core_152;
  wire popcount38_2oru_core_153;
  wire popcount38_2oru_core_154;
  wire popcount38_2oru_core_155;
  wire popcount38_2oru_core_156;
  wire popcount38_2oru_core_157_not;
  wire popcount38_2oru_core_158;
  wire popcount38_2oru_core_160;
  wire popcount38_2oru_core_161;
  wire popcount38_2oru_core_166;
  wire popcount38_2oru_core_168;
  wire popcount38_2oru_core_169;
  wire popcount38_2oru_core_171;
  wire popcount38_2oru_core_174;
  wire popcount38_2oru_core_175;
  wire popcount38_2oru_core_176;
  wire popcount38_2oru_core_177;
  wire popcount38_2oru_core_179;
  wire popcount38_2oru_core_181;
  wire popcount38_2oru_core_182;
  wire popcount38_2oru_core_184;
  wire popcount38_2oru_core_185;
  wire popcount38_2oru_core_186;
  wire popcount38_2oru_core_187;
  wire popcount38_2oru_core_188;
  wire popcount38_2oru_core_189;
  wire popcount38_2oru_core_190;
  wire popcount38_2oru_core_192;
  wire popcount38_2oru_core_193;
  wire popcount38_2oru_core_194;
  wire popcount38_2oru_core_195;
  wire popcount38_2oru_core_197;
  wire popcount38_2oru_core_199;
  wire popcount38_2oru_core_201;
  wire popcount38_2oru_core_202;
  wire popcount38_2oru_core_204;
  wire popcount38_2oru_core_208;
  wire popcount38_2oru_core_209;
  wire popcount38_2oru_core_210_not;
  wire popcount38_2oru_core_213;
  wire popcount38_2oru_core_215;
  wire popcount38_2oru_core_219_not;
  wire popcount38_2oru_core_220;
  wire popcount38_2oru_core_222;
  wire popcount38_2oru_core_223;
  wire popcount38_2oru_core_224;
  wire popcount38_2oru_core_225;
  wire popcount38_2oru_core_227;
  wire popcount38_2oru_core_228;
  wire popcount38_2oru_core_229;
  wire popcount38_2oru_core_231;
  wire popcount38_2oru_core_233;
  wire popcount38_2oru_core_234;
  wire popcount38_2oru_core_235;
  wire popcount38_2oru_core_236;
  wire popcount38_2oru_core_239;
  wire popcount38_2oru_core_241;
  wire popcount38_2oru_core_243;
  wire popcount38_2oru_core_244;
  wire popcount38_2oru_core_245;
  wire popcount38_2oru_core_246;
  wire popcount38_2oru_core_247;
  wire popcount38_2oru_core_249;
  wire popcount38_2oru_core_251;
  wire popcount38_2oru_core_252;
  wire popcount38_2oru_core_254;
  wire popcount38_2oru_core_255;
  wire popcount38_2oru_core_257;
  wire popcount38_2oru_core_258;
  wire popcount38_2oru_core_260;
  wire popcount38_2oru_core_262;
  wire popcount38_2oru_core_263;
  wire popcount38_2oru_core_265;
  wire popcount38_2oru_core_266;
  wire popcount38_2oru_core_267;
  wire popcount38_2oru_core_268;
  wire popcount38_2oru_core_269;
  wire popcount38_2oru_core_270;
  wire popcount38_2oru_core_271;
  wire popcount38_2oru_core_272;
  wire popcount38_2oru_core_273;
  wire popcount38_2oru_core_274;
  wire popcount38_2oru_core_275;
  wire popcount38_2oru_core_277;
  wire popcount38_2oru_core_278;
  wire popcount38_2oru_core_280;
  wire popcount38_2oru_core_281;
  wire popcount38_2oru_core_282_not;
  wire popcount38_2oru_core_283;
  wire popcount38_2oru_core_284;
  wire popcount38_2oru_core_285;
  wire popcount38_2oru_core_286;
  wire popcount38_2oru_core_287;
  wire popcount38_2oru_core_288;
  wire popcount38_2oru_core_289;
  wire popcount38_2oru_core_291;
  wire popcount38_2oru_core_292;
  wire popcount38_2oru_core_295;
  wire popcount38_2oru_core_296;

  assign popcount38_2oru_core_040 = input_a[21] ^ input_a[1];
  assign popcount38_2oru_core_041 = ~(input_a[35] & input_a[37]);
  assign popcount38_2oru_core_042 = ~input_a[28];
  assign popcount38_2oru_core_043 = ~input_a[26];
  assign popcount38_2oru_core_044 = input_a[10] ^ input_a[14];
  assign popcount38_2oru_core_045 = input_a[6] & input_a[15];
  assign popcount38_2oru_core_046 = input_a[7] | input_a[21];
  assign popcount38_2oru_core_048 = ~(input_a[28] & input_a[20]);
  assign popcount38_2oru_core_050 = ~(input_a[26] ^ input_a[36]);
  assign popcount38_2oru_core_051 = input_a[3] | input_a[9];
  assign popcount38_2oru_core_052 = input_a[12] ^ input_a[29];
  assign popcount38_2oru_core_053_not = ~input_a[28];
  assign popcount38_2oru_core_054 = ~input_a[4];
  assign popcount38_2oru_core_055 = ~input_a[0];
  assign popcount38_2oru_core_056 = input_a[25] ^ input_a[5];
  assign popcount38_2oru_core_057 = ~(input_a[13] & input_a[24]);
  assign popcount38_2oru_core_059 = input_a[0] ^ input_a[8];
  assign popcount38_2oru_core_060 = ~(input_a[31] | input_a[8]);
  assign popcount38_2oru_core_061 = input_a[4] ^ input_a[3];
  assign popcount38_2oru_core_066 = ~(input_a[2] ^ input_a[34]);
  assign popcount38_2oru_core_067 = ~(input_a[33] ^ input_a[3]);
  assign popcount38_2oru_core_068 = ~input_a[15];
  assign popcount38_2oru_core_072 = input_a[10] | input_a[13];
  assign popcount38_2oru_core_073 = input_a[30] | input_a[28];
  assign popcount38_2oru_core_076 = input_a[31] ^ input_a[13];
  assign popcount38_2oru_core_077 = input_a[20] | input_a[10];
  assign popcount38_2oru_core_078 = ~input_a[32];
  assign popcount38_2oru_core_079 = ~(input_a[25] & input_a[27]);
  assign popcount38_2oru_core_080 = input_a[20] ^ input_a[24];
  assign popcount38_2oru_core_082 = input_a[8] & input_a[31];
  assign popcount38_2oru_core_084 = ~(input_a[20] & input_a[0]);
  assign popcount38_2oru_core_085 = ~(input_a[2] ^ input_a[15]);
  assign popcount38_2oru_core_086 = input_a[29] ^ input_a[22];
  assign popcount38_2oru_core_087 = input_a[22] & input_a[8];
  assign popcount38_2oru_core_088 = input_a[33] | input_a[25];
  assign popcount38_2oru_core_090 = ~(input_a[0] & input_a[9]);
  assign popcount38_2oru_core_093 = ~(input_a[34] & input_a[25]);
  assign popcount38_2oru_core_094 = ~(input_a[35] | input_a[19]);
  assign popcount38_2oru_core_095 = ~(input_a[31] | input_a[12]);
  assign popcount38_2oru_core_096 = ~(input_a[17] & input_a[24]);
  assign popcount38_2oru_core_097 = input_a[12] | input_a[18];
  assign popcount38_2oru_core_098 = input_a[37] & input_a[15];
  assign popcount38_2oru_core_102 = ~(input_a[8] & input_a[17]);
  assign popcount38_2oru_core_103_not = ~input_a[20];
  assign popcount38_2oru_core_104 = ~(input_a[27] ^ input_a[25]);
  assign popcount38_2oru_core_105 = input_a[5] | input_a[5];
  assign popcount38_2oru_core_106 = input_a[33] ^ input_a[33];
  assign popcount38_2oru_core_110 = input_a[6] | input_a[1];
  assign popcount38_2oru_core_111 = input_a[13] ^ input_a[12];
  assign popcount38_2oru_core_113 = input_a[16] & input_a[18];
  assign popcount38_2oru_core_114 = input_a[9] | input_a[4];
  assign popcount38_2oru_core_115 = input_a[24] | input_a[15];
  assign popcount38_2oru_core_116 = ~input_a[29];
  assign popcount38_2oru_core_121 = input_a[8] ^ input_a[35];
  assign popcount38_2oru_core_122 = ~(input_a[4] ^ input_a[0]);
  assign popcount38_2oru_core_124 = ~(input_a[27] | input_a[32]);
  assign popcount38_2oru_core_126 = ~(input_a[16] | input_a[22]);
  assign popcount38_2oru_core_128 = input_a[14] ^ input_a[10];
  assign popcount38_2oru_core_129 = input_a[12] & input_a[9];
  assign popcount38_2oru_core_131 = input_a[0] | input_a[18];
  assign popcount38_2oru_core_132 = input_a[22] & input_a[12];
  assign popcount38_2oru_core_137 = ~input_a[12];
  assign popcount38_2oru_core_138 = ~input_a[24];
  assign popcount38_2oru_core_139 = input_a[23] | input_a[26];
  assign popcount38_2oru_core_141 = input_a[0] | input_a[28];
  assign popcount38_2oru_core_142 = ~(input_a[10] ^ input_a[18]);
  assign popcount38_2oru_core_143 = input_a[18] & input_a[22];
  assign popcount38_2oru_core_151 = ~input_a[11];
  assign popcount38_2oru_core_152 = input_a[37] & input_a[20];
  assign popcount38_2oru_core_153 = input_a[23] & input_a[25];
  assign popcount38_2oru_core_154 = input_a[0] & input_a[30];
  assign popcount38_2oru_core_155 = ~input_a[7];
  assign popcount38_2oru_core_156 = ~(input_a[29] ^ input_a[27]);
  assign popcount38_2oru_core_157_not = ~input_a[5];
  assign popcount38_2oru_core_158 = ~(input_a[16] | input_a[18]);
  assign popcount38_2oru_core_160 = ~(input_a[9] & input_a[6]);
  assign popcount38_2oru_core_161 = ~(input_a[8] ^ input_a[12]);
  assign popcount38_2oru_core_166 = ~(input_a[8] & input_a[11]);
  assign popcount38_2oru_core_168 = ~input_a[19];
  assign popcount38_2oru_core_169 = input_a[37] | input_a[1];
  assign popcount38_2oru_core_171 = ~(input_a[1] | input_a[19]);
  assign popcount38_2oru_core_174 = ~input_a[2];
  assign popcount38_2oru_core_175 = input_a[28] | input_a[5];
  assign popcount38_2oru_core_176 = ~(input_a[0] ^ input_a[4]);
  assign popcount38_2oru_core_177 = input_a[7] ^ input_a[36];
  assign popcount38_2oru_core_179 = ~(input_a[33] | input_a[35]);
  assign popcount38_2oru_core_181 = input_a[8] | input_a[37];
  assign popcount38_2oru_core_182 = input_a[0] | input_a[29];
  assign popcount38_2oru_core_184 = input_a[2] & input_a[12];
  assign popcount38_2oru_core_185 = ~(input_a[27] | input_a[37]);
  assign popcount38_2oru_core_186 = ~(input_a[33] & input_a[13]);
  assign popcount38_2oru_core_187 = input_a[3] ^ input_a[5];
  assign popcount38_2oru_core_188 = ~(input_a[32] ^ input_a[5]);
  assign popcount38_2oru_core_189 = ~(input_a[2] ^ input_a[26]);
  assign popcount38_2oru_core_190 = input_a[5] | popcount38_2oru_core_181;
  assign popcount38_2oru_core_192 = popcount38_2oru_core_190 | input_a[1];
  assign popcount38_2oru_core_193 = ~(input_a[21] & input_a[8]);
  assign popcount38_2oru_core_194 = input_a[9] ^ input_a[19];
  assign popcount38_2oru_core_195 = ~(input_a[20] ^ input_a[37]);
  assign popcount38_2oru_core_197 = ~input_a[2];
  assign popcount38_2oru_core_199 = ~(input_a[14] ^ input_a[1]);
  assign popcount38_2oru_core_201 = input_a[26] & input_a[24];
  assign popcount38_2oru_core_202 = ~input_a[0];
  assign popcount38_2oru_core_204 = ~(input_a[7] | input_a[35]);
  assign popcount38_2oru_core_208 = ~(input_a[10] ^ input_a[16]);
  assign popcount38_2oru_core_209 = ~input_a[12];
  assign popcount38_2oru_core_210_not = ~input_a[18];
  assign popcount38_2oru_core_213 = input_a[8] ^ input_a[23];
  assign popcount38_2oru_core_215 = ~(input_a[19] ^ input_a[14]);
  assign popcount38_2oru_core_219_not = ~input_a[8];
  assign popcount38_2oru_core_220 = input_a[28] & input_a[7];
  assign popcount38_2oru_core_222 = input_a[7] ^ input_a[2];
  assign popcount38_2oru_core_223 = ~(input_a[26] & input_a[30]);
  assign popcount38_2oru_core_224 = input_a[18] ^ input_a[0];
  assign popcount38_2oru_core_225 = input_a[20] ^ input_a[22];
  assign popcount38_2oru_core_227 = input_a[25] | input_a[27];
  assign popcount38_2oru_core_228 = input_a[37] | input_a[17];
  assign popcount38_2oru_core_229 = input_a[15] ^ input_a[30];
  assign popcount38_2oru_core_231 = ~(input_a[17] ^ input_a[35]);
  assign popcount38_2oru_core_233 = ~(input_a[37] & input_a[4]);
  assign popcount38_2oru_core_234 = ~(input_a[15] | input_a[3]);
  assign popcount38_2oru_core_235 = ~(input_a[35] | input_a[23]);
  assign popcount38_2oru_core_236 = input_a[11] & input_a[15];
  assign popcount38_2oru_core_239 = ~(input_a[36] & input_a[5]);
  assign popcount38_2oru_core_241 = ~(input_a[33] & input_a[16]);
  assign popcount38_2oru_core_243 = ~(input_a[30] & input_a[13]);
  assign popcount38_2oru_core_244 = ~(input_a[22] | input_a[9]);
  assign popcount38_2oru_core_245 = ~(input_a[21] & input_a[6]);
  assign popcount38_2oru_core_246 = input_a[0] ^ input_a[16];
  assign popcount38_2oru_core_247 = ~(input_a[30] & input_a[25]);
  assign popcount38_2oru_core_249 = input_a[28] | input_a[16];
  assign popcount38_2oru_core_251 = ~(input_a[30] ^ input_a[18]);
  assign popcount38_2oru_core_252 = input_a[1] ^ input_a[6];
  assign popcount38_2oru_core_254 = input_a[9] ^ input_a[29];
  assign popcount38_2oru_core_255 = popcount38_2oru_core_192 | input_a[6];
  assign popcount38_2oru_core_257 = ~popcount38_2oru_core_255;
  assign popcount38_2oru_core_258 = input_a[25] | input_a[12];
  assign popcount38_2oru_core_260 = input_a[8] | input_a[19];
  assign popcount38_2oru_core_262 = ~input_a[3];
  assign popcount38_2oru_core_263 = input_a[29] & input_a[28];
  assign popcount38_2oru_core_265 = ~(input_a[9] ^ input_a[19]);
  assign popcount38_2oru_core_266 = ~(input_a[16] ^ input_a[15]);
  assign popcount38_2oru_core_267 = ~(input_a[35] & input_a[0]);
  assign popcount38_2oru_core_268 = input_a[2] ^ input_a[8];
  assign popcount38_2oru_core_269 = input_a[23] ^ input_a[13];
  assign popcount38_2oru_core_270 = ~input_a[21];
  assign popcount38_2oru_core_271 = input_a[32] & input_a[17];
  assign popcount38_2oru_core_272 = input_a[6] & input_a[10];
  assign popcount38_2oru_core_273 = input_a[21] & input_a[28];
  assign popcount38_2oru_core_274 = ~input_a[12];
  assign popcount38_2oru_core_275 = ~(input_a[1] & input_a[2]);
  assign popcount38_2oru_core_277 = input_a[20] | popcount38_2oru_core_257;
  assign popcount38_2oru_core_278 = input_a[4] | input_a[2];
  assign popcount38_2oru_core_280 = ~input_a[8];
  assign popcount38_2oru_core_281 = ~(input_a[15] | input_a[23]);
  assign popcount38_2oru_core_282_not = ~input_a[17];
  assign popcount38_2oru_core_283 = ~(input_a[2] | input_a[35]);
  assign popcount38_2oru_core_284 = input_a[37] ^ input_a[6];
  assign popcount38_2oru_core_285 = ~input_a[32];
  assign popcount38_2oru_core_286 = ~(input_a[21] & input_a[20]);
  assign popcount38_2oru_core_287 = input_a[24] | input_a[18];
  assign popcount38_2oru_core_288 = input_a[25] & input_a[30];
  assign popcount38_2oru_core_289 = input_a[26] | input_a[24];
  assign popcount38_2oru_core_291 = ~(input_a[17] & input_a[11]);
  assign popcount38_2oru_core_292 = input_a[22] & input_a[7];
  assign popcount38_2oru_core_295 = input_a[3] | input_a[1];
  assign popcount38_2oru_core_296 = input_a[29] | input_a[35];

  assign popcount38_2oru_out[0] = input_a[17];
  assign popcount38_2oru_out[1] = input_a[28];
  assign popcount38_2oru_out[2] = popcount38_2oru_core_277;
  assign popcount38_2oru_out[3] = popcount38_2oru_core_257;
  assign popcount38_2oru_out[4] = popcount38_2oru_core_255;
  assign popcount38_2oru_out[5] = 1'b0;
endmodule