// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.25
// WCE=4.0
// EP=0.765625%
// Printed PDK parameters:
//  Area=41206787.0
//  Delay=65198924.0
//  Power=2066600.0

module popcount20_zl4x(input [19:0] input_a, output [4:0] popcount20_zl4x_out);
  wire popcount20_zl4x_core_022;
  wire popcount20_zl4x_core_023;
  wire popcount20_zl4x_core_024;
  wire popcount20_zl4x_core_026;
  wire popcount20_zl4x_core_028;
  wire popcount20_zl4x_core_030;
  wire popcount20_zl4x_core_031;
  wire popcount20_zl4x_core_032;
  wire popcount20_zl4x_core_033;
  wire popcount20_zl4x_core_034;
  wire popcount20_zl4x_core_035;
  wire popcount20_zl4x_core_036;
  wire popcount20_zl4x_core_038;
  wire popcount20_zl4x_core_039;
  wire popcount20_zl4x_core_040;
  wire popcount20_zl4x_core_041;
  wire popcount20_zl4x_core_042;
  wire popcount20_zl4x_core_044;
  wire popcount20_zl4x_core_045;
  wire popcount20_zl4x_core_047_not;
  wire popcount20_zl4x_core_048;
  wire popcount20_zl4x_core_049;
  wire popcount20_zl4x_core_050;
  wire popcount20_zl4x_core_051;
  wire popcount20_zl4x_core_052;
  wire popcount20_zl4x_core_053;
  wire popcount20_zl4x_core_056;
  wire popcount20_zl4x_core_058;
  wire popcount20_zl4x_core_059;
  wire popcount20_zl4x_core_061;
  wire popcount20_zl4x_core_063;
  wire popcount20_zl4x_core_064;
  wire popcount20_zl4x_core_065;
  wire popcount20_zl4x_core_066;
  wire popcount20_zl4x_core_067;
  wire popcount20_zl4x_core_071;
  wire popcount20_zl4x_core_073;
  wire popcount20_zl4x_core_075;
  wire popcount20_zl4x_core_076;
  wire popcount20_zl4x_core_077;
  wire popcount20_zl4x_core_078;
  wire popcount20_zl4x_core_079;
  wire popcount20_zl4x_core_082;
  wire popcount20_zl4x_core_083;
  wire popcount20_zl4x_core_084;
  wire popcount20_zl4x_core_086;
  wire popcount20_zl4x_core_089;
  wire popcount20_zl4x_core_090;
  wire popcount20_zl4x_core_091;
  wire popcount20_zl4x_core_092;
  wire popcount20_zl4x_core_093;
  wire popcount20_zl4x_core_094;
  wire popcount20_zl4x_core_095;
  wire popcount20_zl4x_core_096;
  wire popcount20_zl4x_core_098;
  wire popcount20_zl4x_core_099;
  wire popcount20_zl4x_core_100;
  wire popcount20_zl4x_core_101;
  wire popcount20_zl4x_core_102;
  wire popcount20_zl4x_core_103;
  wire popcount20_zl4x_core_104;
  wire popcount20_zl4x_core_106;
  wire popcount20_zl4x_core_107;
  wire popcount20_zl4x_core_108;
  wire popcount20_zl4x_core_109;
  wire popcount20_zl4x_core_110;
  wire popcount20_zl4x_core_111;
  wire popcount20_zl4x_core_112;
  wire popcount20_zl4x_core_113;
  wire popcount20_zl4x_core_114;
  wire popcount20_zl4x_core_115;
  wire popcount20_zl4x_core_116;
  wire popcount20_zl4x_core_117;
  wire popcount20_zl4x_core_118;
  wire popcount20_zl4x_core_120;
  wire popcount20_zl4x_core_123;
  wire popcount20_zl4x_core_124;
  wire popcount20_zl4x_core_126;
  wire popcount20_zl4x_core_127;
  wire popcount20_zl4x_core_128;
  wire popcount20_zl4x_core_131;
  wire popcount20_zl4x_core_132;
  wire popcount20_zl4x_core_133;
  wire popcount20_zl4x_core_134;
  wire popcount20_zl4x_core_135;
  wire popcount20_zl4x_core_136;
  wire popcount20_zl4x_core_137;
  wire popcount20_zl4x_core_138;
  wire popcount20_zl4x_core_139;
  wire popcount20_zl4x_core_140;
  wire popcount20_zl4x_core_141;
  wire popcount20_zl4x_core_142;
  wire popcount20_zl4x_core_143;

  assign popcount20_zl4x_core_022 = input_a[0] ^ input_a[1];
  assign popcount20_zl4x_core_023 = input_a[0] & input_a[1];
  assign popcount20_zl4x_core_024 = ~input_a[3];
  assign popcount20_zl4x_core_026 = input_a[2] ^ popcount20_zl4x_core_024;
  assign popcount20_zl4x_core_028 = input_a[3] | input_a[2];
  assign popcount20_zl4x_core_030 = ~input_a[7];
  assign popcount20_zl4x_core_031 = popcount20_zl4x_core_022 & popcount20_zl4x_core_026;
  assign popcount20_zl4x_core_032 = popcount20_zl4x_core_023 ^ popcount20_zl4x_core_028;
  assign popcount20_zl4x_core_033 = popcount20_zl4x_core_023 & popcount20_zl4x_core_028;
  assign popcount20_zl4x_core_034 = popcount20_zl4x_core_032 ^ popcount20_zl4x_core_031;
  assign popcount20_zl4x_core_035 = input_a[3] & popcount20_zl4x_core_031;
  assign popcount20_zl4x_core_036 = popcount20_zl4x_core_033 | popcount20_zl4x_core_035;
  assign popcount20_zl4x_core_038 = ~(input_a[5] & input_a[11]);
  assign popcount20_zl4x_core_039 = ~(input_a[18] | input_a[6]);
  assign popcount20_zl4x_core_040 = input_a[10] & input_a[6];
  assign popcount20_zl4x_core_041 = input_a[8] | input_a[9];
  assign popcount20_zl4x_core_042 = input_a[8] & input_a[9];
  assign popcount20_zl4x_core_044 = input_a[7] & popcount20_zl4x_core_041;
  assign popcount20_zl4x_core_045 = popcount20_zl4x_core_042 | popcount20_zl4x_core_044;
  assign popcount20_zl4x_core_047_not = ~input_a[18];
  assign popcount20_zl4x_core_048 = input_a[7] & input_a[6];
  assign popcount20_zl4x_core_049 = popcount20_zl4x_core_040 ^ popcount20_zl4x_core_045;
  assign popcount20_zl4x_core_050 = popcount20_zl4x_core_040 & popcount20_zl4x_core_045;
  assign popcount20_zl4x_core_051 = popcount20_zl4x_core_049 ^ input_a[11];
  assign popcount20_zl4x_core_052 = popcount20_zl4x_core_049 & input_a[11];
  assign popcount20_zl4x_core_053 = popcount20_zl4x_core_050 | popcount20_zl4x_core_052;
  assign popcount20_zl4x_core_056 = ~(input_a[13] ^ input_a[10]);
  assign popcount20_zl4x_core_058 = popcount20_zl4x_core_034 ^ popcount20_zl4x_core_051;
  assign popcount20_zl4x_core_059 = popcount20_zl4x_core_034 & popcount20_zl4x_core_051;
  assign popcount20_zl4x_core_061 = ~(input_a[0] & input_a[12]);
  assign popcount20_zl4x_core_063 = popcount20_zl4x_core_036 ^ popcount20_zl4x_core_053;
  assign popcount20_zl4x_core_064 = popcount20_zl4x_core_036 & popcount20_zl4x_core_053;
  assign popcount20_zl4x_core_065 = popcount20_zl4x_core_063 ^ popcount20_zl4x_core_059;
  assign popcount20_zl4x_core_066 = popcount20_zl4x_core_063 & popcount20_zl4x_core_059;
  assign popcount20_zl4x_core_067 = popcount20_zl4x_core_064 | popcount20_zl4x_core_066;
  assign popcount20_zl4x_core_071 = input_a[2] ^ input_a[13];
  assign popcount20_zl4x_core_073 = ~input_a[4];
  assign popcount20_zl4x_core_075 = ~input_a[2];
  assign popcount20_zl4x_core_076 = input_a[18] | input_a[0];
  assign popcount20_zl4x_core_077 = ~input_a[17];
  assign popcount20_zl4x_core_078 = input_a[5] | input_a[8];
  assign popcount20_zl4x_core_079 = input_a[4] | input_a[12];
  assign popcount20_zl4x_core_082 = input_a[17] & input_a[14];
  assign popcount20_zl4x_core_083 = ~input_a[13];
  assign popcount20_zl4x_core_084 = input_a[13] & popcount20_zl4x_core_079;
  assign popcount20_zl4x_core_086 = ~input_a[16];
  assign popcount20_zl4x_core_089 = input_a[12] | input_a[6];
  assign popcount20_zl4x_core_090 = input_a[15] ^ input_a[16];
  assign popcount20_zl4x_core_091 = input_a[15] & input_a[16];
  assign popcount20_zl4x_core_092 = input_a[18] ^ input_a[19];
  assign popcount20_zl4x_core_093 = input_a[18] & input_a[19];
  assign popcount20_zl4x_core_094 = input_a[17] ^ popcount20_zl4x_core_092;
  assign popcount20_zl4x_core_095 = input_a[17] & popcount20_zl4x_core_092;
  assign popcount20_zl4x_core_096 = popcount20_zl4x_core_093 | popcount20_zl4x_core_095;
  assign popcount20_zl4x_core_098 = popcount20_zl4x_core_090 ^ popcount20_zl4x_core_094;
  assign popcount20_zl4x_core_099 = popcount20_zl4x_core_090 & popcount20_zl4x_core_094;
  assign popcount20_zl4x_core_100 = popcount20_zl4x_core_091 ^ popcount20_zl4x_core_096;
  assign popcount20_zl4x_core_101 = popcount20_zl4x_core_091 & popcount20_zl4x_core_096;
  assign popcount20_zl4x_core_102 = popcount20_zl4x_core_100 ^ popcount20_zl4x_core_099;
  assign popcount20_zl4x_core_103 = popcount20_zl4x_core_100 & popcount20_zl4x_core_099;
  assign popcount20_zl4x_core_104 = popcount20_zl4x_core_101 | popcount20_zl4x_core_103;
  assign popcount20_zl4x_core_106 = ~input_a[15];
  assign popcount20_zl4x_core_107 = input_a[7] & input_a[13];
  assign popcount20_zl4x_core_108 = input_a[5] & popcount20_zl4x_core_098;
  assign popcount20_zl4x_core_109 = popcount20_zl4x_core_083 ^ popcount20_zl4x_core_102;
  assign popcount20_zl4x_core_110 = popcount20_zl4x_core_083 & popcount20_zl4x_core_102;
  assign popcount20_zl4x_core_111 = popcount20_zl4x_core_109 ^ popcount20_zl4x_core_108;
  assign popcount20_zl4x_core_112 = popcount20_zl4x_core_109 & popcount20_zl4x_core_108;
  assign popcount20_zl4x_core_113 = popcount20_zl4x_core_110 | popcount20_zl4x_core_112;
  assign popcount20_zl4x_core_114 = popcount20_zl4x_core_084 ^ popcount20_zl4x_core_104;
  assign popcount20_zl4x_core_115 = popcount20_zl4x_core_084 & popcount20_zl4x_core_104;
  assign popcount20_zl4x_core_116 = popcount20_zl4x_core_114 ^ popcount20_zl4x_core_113;
  assign popcount20_zl4x_core_117 = popcount20_zl4x_core_114 & popcount20_zl4x_core_113;
  assign popcount20_zl4x_core_118 = popcount20_zl4x_core_115 | popcount20_zl4x_core_117;
  assign popcount20_zl4x_core_120 = input_a[6] | input_a[0];
  assign popcount20_zl4x_core_123 = ~(input_a[17] & input_a[12]);
  assign popcount20_zl4x_core_124 = ~(input_a[7] & input_a[15]);
  assign popcount20_zl4x_core_126 = popcount20_zl4x_core_058 ^ popcount20_zl4x_core_111;
  assign popcount20_zl4x_core_127 = popcount20_zl4x_core_058 & popcount20_zl4x_core_111;
  assign popcount20_zl4x_core_128 = input_a[4] | input_a[18];
  assign popcount20_zl4x_core_131 = popcount20_zl4x_core_065 ^ popcount20_zl4x_core_116;
  assign popcount20_zl4x_core_132 = popcount20_zl4x_core_065 & popcount20_zl4x_core_116;
  assign popcount20_zl4x_core_133 = popcount20_zl4x_core_131 ^ popcount20_zl4x_core_127;
  assign popcount20_zl4x_core_134 = popcount20_zl4x_core_131 & popcount20_zl4x_core_127;
  assign popcount20_zl4x_core_135 = popcount20_zl4x_core_132 | popcount20_zl4x_core_134;
  assign popcount20_zl4x_core_136 = popcount20_zl4x_core_067 ^ popcount20_zl4x_core_118;
  assign popcount20_zl4x_core_137 = popcount20_zl4x_core_067 & popcount20_zl4x_core_118;
  assign popcount20_zl4x_core_138 = popcount20_zl4x_core_136 ^ popcount20_zl4x_core_135;
  assign popcount20_zl4x_core_139 = popcount20_zl4x_core_136 & popcount20_zl4x_core_135;
  assign popcount20_zl4x_core_140 = popcount20_zl4x_core_137 | popcount20_zl4x_core_139;
  assign popcount20_zl4x_core_141 = ~(input_a[12] | input_a[3]);
  assign popcount20_zl4x_core_142 = ~input_a[18];
  assign popcount20_zl4x_core_143 = input_a[0] ^ input_a[18];

  assign popcount20_zl4x_out[0] = input_a[14];
  assign popcount20_zl4x_out[1] = popcount20_zl4x_core_126;
  assign popcount20_zl4x_out[2] = popcount20_zl4x_core_133;
  assign popcount20_zl4x_out[3] = popcount20_zl4x_core_138;
  assign popcount20_zl4x_out[4] = popcount20_zl4x_core_140;
endmodule