// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=2.37915
// WCE=17.0
// EP=0.868282%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount33_5zjr(input [32:0] input_a, output [5:0] popcount33_5zjr_out);
  wire popcount33_5zjr_core_035;
  wire popcount33_5zjr_core_037;
  wire popcount33_5zjr_core_038;
  wire popcount33_5zjr_core_040_not;
  wire popcount33_5zjr_core_041;
  wire popcount33_5zjr_core_042;
  wire popcount33_5zjr_core_043;
  wire popcount33_5zjr_core_044;
  wire popcount33_5zjr_core_045;
  wire popcount33_5zjr_core_051;
  wire popcount33_5zjr_core_052;
  wire popcount33_5zjr_core_053;
  wire popcount33_5zjr_core_056;
  wire popcount33_5zjr_core_057;
  wire popcount33_5zjr_core_060;
  wire popcount33_5zjr_core_061;
  wire popcount33_5zjr_core_062;
  wire popcount33_5zjr_core_064;
  wire popcount33_5zjr_core_065;
  wire popcount33_5zjr_core_066;
  wire popcount33_5zjr_core_067;
  wire popcount33_5zjr_core_068;
  wire popcount33_5zjr_core_069;
  wire popcount33_5zjr_core_071;
  wire popcount33_5zjr_core_072;
  wire popcount33_5zjr_core_073;
  wire popcount33_5zjr_core_074;
  wire popcount33_5zjr_core_075;
  wire popcount33_5zjr_core_076;
  wire popcount33_5zjr_core_079;
  wire popcount33_5zjr_core_080;
  wire popcount33_5zjr_core_081;
  wire popcount33_5zjr_core_084;
  wire popcount33_5zjr_core_085;
  wire popcount33_5zjr_core_086;
  wire popcount33_5zjr_core_087;
  wire popcount33_5zjr_core_088;
  wire popcount33_5zjr_core_090;
  wire popcount33_5zjr_core_091;
  wire popcount33_5zjr_core_092;
  wire popcount33_5zjr_core_093;
  wire popcount33_5zjr_core_094;
  wire popcount33_5zjr_core_095;
  wire popcount33_5zjr_core_096;
  wire popcount33_5zjr_core_097;
  wire popcount33_5zjr_core_098;
  wire popcount33_5zjr_core_099;
  wire popcount33_5zjr_core_100;
  wire popcount33_5zjr_core_101;
  wire popcount33_5zjr_core_103;
  wire popcount33_5zjr_core_104;
  wire popcount33_5zjr_core_106_not;
  wire popcount33_5zjr_core_107;
  wire popcount33_5zjr_core_108;
  wire popcount33_5zjr_core_109;
  wire popcount33_5zjr_core_110;
  wire popcount33_5zjr_core_111;
  wire popcount33_5zjr_core_114;
  wire popcount33_5zjr_core_116;
  wire popcount33_5zjr_core_117;
  wire popcount33_5zjr_core_118;
  wire popcount33_5zjr_core_119;
  wire popcount33_5zjr_core_123;
  wire popcount33_5zjr_core_124;
  wire popcount33_5zjr_core_126;
  wire popcount33_5zjr_core_130;
  wire popcount33_5zjr_core_132;
  wire popcount33_5zjr_core_133;
  wire popcount33_5zjr_core_135;
  wire popcount33_5zjr_core_136;
  wire popcount33_5zjr_core_137_not;
  wire popcount33_5zjr_core_140;
  wire popcount33_5zjr_core_141;
  wire popcount33_5zjr_core_143;
  wire popcount33_5zjr_core_145;
  wire popcount33_5zjr_core_148;
  wire popcount33_5zjr_core_149;
  wire popcount33_5zjr_core_152;
  wire popcount33_5zjr_core_154;
  wire popcount33_5zjr_core_155_not;
  wire popcount33_5zjr_core_156;
  wire popcount33_5zjr_core_157;
  wire popcount33_5zjr_core_158;
  wire popcount33_5zjr_core_159;
  wire popcount33_5zjr_core_161;
  wire popcount33_5zjr_core_162;
  wire popcount33_5zjr_core_165;
  wire popcount33_5zjr_core_167;
  wire popcount33_5zjr_core_168;
  wire popcount33_5zjr_core_169;
  wire popcount33_5zjr_core_170;
  wire popcount33_5zjr_core_173;
  wire popcount33_5zjr_core_174;
  wire popcount33_5zjr_core_176;
  wire popcount33_5zjr_core_177;
  wire popcount33_5zjr_core_178;
  wire popcount33_5zjr_core_179;
  wire popcount33_5zjr_core_180;
  wire popcount33_5zjr_core_182;
  wire popcount33_5zjr_core_183;
  wire popcount33_5zjr_core_185;
  wire popcount33_5zjr_core_186;
  wire popcount33_5zjr_core_188;
  wire popcount33_5zjr_core_190;
  wire popcount33_5zjr_core_191;
  wire popcount33_5zjr_core_198;
  wire popcount33_5zjr_core_200_not;
  wire popcount33_5zjr_core_201;
  wire popcount33_5zjr_core_202;
  wire popcount33_5zjr_core_204;
  wire popcount33_5zjr_core_206;
  wire popcount33_5zjr_core_207;
  wire popcount33_5zjr_core_208;
  wire popcount33_5zjr_core_210;
  wire popcount33_5zjr_core_211;
  wire popcount33_5zjr_core_212;
  wire popcount33_5zjr_core_213;
  wire popcount33_5zjr_core_216;
  wire popcount33_5zjr_core_217;
  wire popcount33_5zjr_core_218;
  wire popcount33_5zjr_core_219;
  wire popcount33_5zjr_core_220;
  wire popcount33_5zjr_core_221;
  wire popcount33_5zjr_core_222;
  wire popcount33_5zjr_core_225;
  wire popcount33_5zjr_core_227;
  wire popcount33_5zjr_core_231;
  wire popcount33_5zjr_core_232;
  wire popcount33_5zjr_core_233;
  wire popcount33_5zjr_core_235;
  wire popcount33_5zjr_core_236;
  wire popcount33_5zjr_core_237;

  assign popcount33_5zjr_core_035 = ~(input_a[7] ^ input_a[25]);
  assign popcount33_5zjr_core_037 = ~(input_a[21] ^ input_a[23]);
  assign popcount33_5zjr_core_038 = input_a[0] ^ input_a[3];
  assign popcount33_5zjr_core_040_not = ~input_a[32];
  assign popcount33_5zjr_core_041 = input_a[21] | input_a[16];
  assign popcount33_5zjr_core_042 = ~(input_a[1] | input_a[25]);
  assign popcount33_5zjr_core_043 = input_a[2] & input_a[4];
  assign popcount33_5zjr_core_044 = ~input_a[4];
  assign popcount33_5zjr_core_045 = input_a[23] ^ input_a[15];
  assign popcount33_5zjr_core_051 = ~input_a[0];
  assign popcount33_5zjr_core_052 = ~input_a[17];
  assign popcount33_5zjr_core_053 = input_a[16] & input_a[23];
  assign popcount33_5zjr_core_056 = ~input_a[4];
  assign popcount33_5zjr_core_057 = input_a[6] ^ input_a[9];
  assign popcount33_5zjr_core_060 = ~input_a[6];
  assign popcount33_5zjr_core_061 = input_a[20] ^ input_a[20];
  assign popcount33_5zjr_core_062 = input_a[12] ^ input_a[24];
  assign popcount33_5zjr_core_064 = ~(input_a[7] | input_a[7]);
  assign popcount33_5zjr_core_065 = input_a[2] & input_a[1];
  assign popcount33_5zjr_core_066 = input_a[0] & input_a[26];
  assign popcount33_5zjr_core_067 = ~(input_a[29] | input_a[0]);
  assign popcount33_5zjr_core_068 = input_a[32] | input_a[10];
  assign popcount33_5zjr_core_069 = input_a[6] ^ input_a[1];
  assign popcount33_5zjr_core_071 = ~(input_a[11] ^ input_a[0]);
  assign popcount33_5zjr_core_072 = input_a[7] & input_a[19];
  assign popcount33_5zjr_core_073 = ~input_a[27];
  assign popcount33_5zjr_core_074 = ~(input_a[9] & input_a[10]);
  assign popcount33_5zjr_core_075 = input_a[32] | input_a[18];
  assign popcount33_5zjr_core_076 = input_a[31] | input_a[12];
  assign popcount33_5zjr_core_079 = ~input_a[22];
  assign popcount33_5zjr_core_080 = input_a[2] | input_a[13];
  assign popcount33_5zjr_core_081 = input_a[1] | input_a[11];
  assign popcount33_5zjr_core_084 = ~(input_a[20] ^ input_a[3]);
  assign popcount33_5zjr_core_085 = ~(input_a[32] ^ input_a[7]);
  assign popcount33_5zjr_core_086 = input_a[27] | input_a[14];
  assign popcount33_5zjr_core_087 = input_a[24] ^ input_a[26];
  assign popcount33_5zjr_core_088 = ~input_a[10];
  assign popcount33_5zjr_core_090 = input_a[24] | input_a[29];
  assign popcount33_5zjr_core_091 = ~(input_a[23] | input_a[11]);
  assign popcount33_5zjr_core_092 = ~(input_a[27] & input_a[11]);
  assign popcount33_5zjr_core_093 = ~input_a[9];
  assign popcount33_5zjr_core_094 = ~input_a[13];
  assign popcount33_5zjr_core_095 = input_a[17] | input_a[21];
  assign popcount33_5zjr_core_096 = ~(input_a[18] ^ input_a[1]);
  assign popcount33_5zjr_core_097 = ~(input_a[32] | input_a[26]);
  assign popcount33_5zjr_core_098 = ~input_a[6];
  assign popcount33_5zjr_core_099 = ~(input_a[11] & input_a[2]);
  assign popcount33_5zjr_core_100 = ~(input_a[27] | input_a[7]);
  assign popcount33_5zjr_core_101 = ~(input_a[26] & input_a[20]);
  assign popcount33_5zjr_core_103 = ~input_a[26];
  assign popcount33_5zjr_core_104 = input_a[18] | input_a[15];
  assign popcount33_5zjr_core_106_not = ~input_a[10];
  assign popcount33_5zjr_core_107 = input_a[27] & input_a[0];
  assign popcount33_5zjr_core_108 = ~input_a[23];
  assign popcount33_5zjr_core_109 = ~(input_a[14] | input_a[0]);
  assign popcount33_5zjr_core_110 = ~input_a[19];
  assign popcount33_5zjr_core_111 = input_a[31] & input_a[30];
  assign popcount33_5zjr_core_114 = ~(input_a[8] ^ input_a[3]);
  assign popcount33_5zjr_core_116 = ~(input_a[4] & input_a[11]);
  assign popcount33_5zjr_core_117 = ~input_a[19];
  assign popcount33_5zjr_core_118 = ~input_a[0];
  assign popcount33_5zjr_core_119 = input_a[29] | input_a[20];
  assign popcount33_5zjr_core_123 = ~(input_a[29] & input_a[19]);
  assign popcount33_5zjr_core_124 = ~(input_a[9] | input_a[18]);
  assign popcount33_5zjr_core_126 = input_a[32] & input_a[22];
  assign popcount33_5zjr_core_130 = ~(input_a[8] | input_a[30]);
  assign popcount33_5zjr_core_132 = ~(input_a[17] & input_a[13]);
  assign popcount33_5zjr_core_133 = ~(input_a[2] & input_a[21]);
  assign popcount33_5zjr_core_135 = ~(input_a[23] ^ input_a[4]);
  assign popcount33_5zjr_core_136 = input_a[13] | input_a[16];
  assign popcount33_5zjr_core_137_not = ~input_a[13];
  assign popcount33_5zjr_core_140 = ~(input_a[8] ^ input_a[29]);
  assign popcount33_5zjr_core_141 = input_a[7] & input_a[6];
  assign popcount33_5zjr_core_143 = input_a[7] & input_a[0];
  assign popcount33_5zjr_core_145 = input_a[23] & input_a[19];
  assign popcount33_5zjr_core_148 = ~input_a[20];
  assign popcount33_5zjr_core_149 = input_a[7] ^ input_a[1];
  assign popcount33_5zjr_core_152 = input_a[4] ^ input_a[10];
  assign popcount33_5zjr_core_154 = ~(input_a[26] ^ input_a[11]);
  assign popcount33_5zjr_core_155_not = ~input_a[32];
  assign popcount33_5zjr_core_156 = input_a[15] & input_a[21];
  assign popcount33_5zjr_core_157 = input_a[15] & input_a[9];
  assign popcount33_5zjr_core_158 = input_a[30] & input_a[1];
  assign popcount33_5zjr_core_159 = input_a[16] & input_a[16];
  assign popcount33_5zjr_core_161 = ~(input_a[7] ^ input_a[13]);
  assign popcount33_5zjr_core_162 = ~(input_a[0] & input_a[29]);
  assign popcount33_5zjr_core_165 = input_a[26] | input_a[15];
  assign popcount33_5zjr_core_167 = ~input_a[3];
  assign popcount33_5zjr_core_168 = input_a[29] | input_a[31];
  assign popcount33_5zjr_core_169 = ~(input_a[18] ^ input_a[4]);
  assign popcount33_5zjr_core_170 = ~input_a[11];
  assign popcount33_5zjr_core_173 = ~(input_a[9] | input_a[19]);
  assign popcount33_5zjr_core_174 = ~(input_a[20] & input_a[13]);
  assign popcount33_5zjr_core_176 = input_a[11] | input_a[15];
  assign popcount33_5zjr_core_177 = ~(input_a[26] & input_a[4]);
  assign popcount33_5zjr_core_178 = ~(input_a[28] | input_a[1]);
  assign popcount33_5zjr_core_179 = ~input_a[8];
  assign popcount33_5zjr_core_180 = input_a[1] ^ input_a[10];
  assign popcount33_5zjr_core_182 = ~(input_a[20] ^ input_a[3]);
  assign popcount33_5zjr_core_183 = input_a[2] | input_a[26];
  assign popcount33_5zjr_core_185 = ~input_a[13];
  assign popcount33_5zjr_core_186 = input_a[0] | input_a[15];
  assign popcount33_5zjr_core_188 = input_a[32] | input_a[21];
  assign popcount33_5zjr_core_190 = ~input_a[32];
  assign popcount33_5zjr_core_191 = ~(input_a[31] & input_a[30]);
  assign popcount33_5zjr_core_198 = input_a[30] | input_a[8];
  assign popcount33_5zjr_core_200_not = ~input_a[18];
  assign popcount33_5zjr_core_201 = input_a[21] | input_a[12];
  assign popcount33_5zjr_core_202 = input_a[7] & input_a[12];
  assign popcount33_5zjr_core_204 = input_a[17] ^ input_a[4];
  assign popcount33_5zjr_core_206 = ~input_a[21];
  assign popcount33_5zjr_core_207 = ~(input_a[32] & input_a[18]);
  assign popcount33_5zjr_core_208 = ~(input_a[1] & input_a[20]);
  assign popcount33_5zjr_core_210 = ~(input_a[27] | input_a[30]);
  assign popcount33_5zjr_core_211 = input_a[27] | input_a[28];
  assign popcount33_5zjr_core_212 = input_a[9] & input_a[13];
  assign popcount33_5zjr_core_213 = input_a[0] & input_a[2];
  assign popcount33_5zjr_core_216 = input_a[30] ^ input_a[31];
  assign popcount33_5zjr_core_217 = input_a[32] | input_a[29];
  assign popcount33_5zjr_core_218 = ~(input_a[13] & input_a[8]);
  assign popcount33_5zjr_core_219 = input_a[22] ^ input_a[8];
  assign popcount33_5zjr_core_220 = ~(input_a[15] & input_a[5]);
  assign popcount33_5zjr_core_221 = input_a[4] ^ input_a[7];
  assign popcount33_5zjr_core_222 = input_a[29] | input_a[30];
  assign popcount33_5zjr_core_225 = input_a[22] ^ input_a[9];
  assign popcount33_5zjr_core_227 = ~input_a[18];
  assign popcount33_5zjr_core_231 = input_a[24] ^ input_a[12];
  assign popcount33_5zjr_core_232 = ~(input_a[8] & input_a[15]);
  assign popcount33_5zjr_core_233 = input_a[24] | input_a[30];
  assign popcount33_5zjr_core_235 = ~(input_a[21] | input_a[31]);
  assign popcount33_5zjr_core_236 = input_a[1] | input_a[7];
  assign popcount33_5zjr_core_237 = ~(input_a[19] | input_a[12]);

  assign popcount33_5zjr_out[0] = input_a[29];
  assign popcount33_5zjr_out[1] = input_a[9];
  assign popcount33_5zjr_out[2] = 1'b0;
  assign popcount33_5zjr_out[3] = 1'b0;
  assign popcount33_5zjr_out[4] = 1'b1;
  assign popcount33_5zjr_out[5] = 1'b0;
endmodule