// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=6.72199
// WCE=24.0
// EP=0.958637%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount28_elja(input [27:0] input_a, output [4:0] popcount28_elja_out);
  wire popcount28_elja_core_031;
  wire popcount28_elja_core_032;
  wire popcount28_elja_core_033;
  wire popcount28_elja_core_034;
  wire popcount28_elja_core_036;
  wire popcount28_elja_core_037;
  wire popcount28_elja_core_040_not;
  wire popcount28_elja_core_042;
  wire popcount28_elja_core_043;
  wire popcount28_elja_core_050;
  wire popcount28_elja_core_051;
  wire popcount28_elja_core_052;
  wire popcount28_elja_core_054;
  wire popcount28_elja_core_055;
  wire popcount28_elja_core_056;
  wire popcount28_elja_core_061;
  wire popcount28_elja_core_063;
  wire popcount28_elja_core_065;
  wire popcount28_elja_core_066;
  wire popcount28_elja_core_067;
  wire popcount28_elja_core_069;
  wire popcount28_elja_core_072;
  wire popcount28_elja_core_073;
  wire popcount28_elja_core_074;
  wire popcount28_elja_core_075;
  wire popcount28_elja_core_076;
  wire popcount28_elja_core_078;
  wire popcount28_elja_core_079;
  wire popcount28_elja_core_080;
  wire popcount28_elja_core_084;
  wire popcount28_elja_core_086;
  wire popcount28_elja_core_089;
  wire popcount28_elja_core_090;
  wire popcount28_elja_core_094;
  wire popcount28_elja_core_097;
  wire popcount28_elja_core_098;
  wire popcount28_elja_core_100;
  wire popcount28_elja_core_102;
  wire popcount28_elja_core_103;
  wire popcount28_elja_core_104;
  wire popcount28_elja_core_105;
  wire popcount28_elja_core_107;
  wire popcount28_elja_core_110;
  wire popcount28_elja_core_112;
  wire popcount28_elja_core_113;
  wire popcount28_elja_core_114;
  wire popcount28_elja_core_115;
  wire popcount28_elja_core_116;
  wire popcount28_elja_core_117;
  wire popcount28_elja_core_118;
  wire popcount28_elja_core_119;
  wire popcount28_elja_core_120;
  wire popcount28_elja_core_121;
  wire popcount28_elja_core_123;
  wire popcount28_elja_core_124;
  wire popcount28_elja_core_125;
  wire popcount28_elja_core_128;
  wire popcount28_elja_core_129;
  wire popcount28_elja_core_130;
  wire popcount28_elja_core_131;
  wire popcount28_elja_core_132;
  wire popcount28_elja_core_134;
  wire popcount28_elja_core_135;
  wire popcount28_elja_core_136_not;
  wire popcount28_elja_core_138_not;
  wire popcount28_elja_core_139;
  wire popcount28_elja_core_141;
  wire popcount28_elja_core_142;
  wire popcount28_elja_core_144;
  wire popcount28_elja_core_145;
  wire popcount28_elja_core_146;
  wire popcount28_elja_core_147;
  wire popcount28_elja_core_148;
  wire popcount28_elja_core_149;
  wire popcount28_elja_core_150;
  wire popcount28_elja_core_151;
  wire popcount28_elja_core_153;
  wire popcount28_elja_core_154;
  wire popcount28_elja_core_158;
  wire popcount28_elja_core_160;
  wire popcount28_elja_core_163;
  wire popcount28_elja_core_165;
  wire popcount28_elja_core_167;
  wire popcount28_elja_core_168;
  wire popcount28_elja_core_170;
  wire popcount28_elja_core_171;
  wire popcount28_elja_core_174;
  wire popcount28_elja_core_175;
  wire popcount28_elja_core_176;
  wire popcount28_elja_core_177;
  wire popcount28_elja_core_178;
  wire popcount28_elja_core_179;
  wire popcount28_elja_core_180;
  wire popcount28_elja_core_183;
  wire popcount28_elja_core_184;
  wire popcount28_elja_core_188;
  wire popcount28_elja_core_190;
  wire popcount28_elja_core_191;
  wire popcount28_elja_core_192;
  wire popcount28_elja_core_194;
  wire popcount28_elja_core_197_not;
  wire popcount28_elja_core_199;
  wire popcount28_elja_core_200;

  assign popcount28_elja_core_031 = ~(input_a[12] ^ input_a[21]);
  assign popcount28_elja_core_032 = ~(input_a[16] & input_a[22]);
  assign popcount28_elja_core_033 = ~input_a[8];
  assign popcount28_elja_core_034 = input_a[25] ^ input_a[19];
  assign popcount28_elja_core_036 = input_a[8] | input_a[17];
  assign popcount28_elja_core_037 = ~input_a[5];
  assign popcount28_elja_core_040_not = ~input_a[2];
  assign popcount28_elja_core_042 = ~(input_a[27] | input_a[2]);
  assign popcount28_elja_core_043 = ~input_a[20];
  assign popcount28_elja_core_050 = input_a[22] ^ input_a[5];
  assign popcount28_elja_core_051 = ~input_a[9];
  assign popcount28_elja_core_052 = ~(input_a[7] & input_a[9]);
  assign popcount28_elja_core_054 = ~input_a[23];
  assign popcount28_elja_core_055 = input_a[17] | input_a[1];
  assign popcount28_elja_core_056 = ~input_a[1];
  assign popcount28_elja_core_061 = ~(input_a[9] ^ input_a[6]);
  assign popcount28_elja_core_063 = ~(input_a[8] & input_a[5]);
  assign popcount28_elja_core_065 = ~(input_a[0] & input_a[14]);
  assign popcount28_elja_core_066 = ~(input_a[15] | input_a[26]);
  assign popcount28_elja_core_067 = ~input_a[0];
  assign popcount28_elja_core_069 = input_a[14] & input_a[9];
  assign popcount28_elja_core_072 = ~(input_a[2] ^ input_a[0]);
  assign popcount28_elja_core_073 = input_a[16] | input_a[19];
  assign popcount28_elja_core_074 = ~(input_a[15] & input_a[3]);
  assign popcount28_elja_core_075 = input_a[4] & input_a[15];
  assign popcount28_elja_core_076 = input_a[26] & input_a[14];
  assign popcount28_elja_core_078 = ~input_a[0];
  assign popcount28_elja_core_079 = ~(input_a[3] | input_a[8]);
  assign popcount28_elja_core_080 = ~input_a[0];
  assign popcount28_elja_core_084 = ~input_a[19];
  assign popcount28_elja_core_086 = ~(input_a[24] & input_a[27]);
  assign popcount28_elja_core_089 = ~(input_a[25] | input_a[9]);
  assign popcount28_elja_core_090 = ~input_a[1];
  assign popcount28_elja_core_094 = ~(input_a[21] ^ input_a[20]);
  assign popcount28_elja_core_097 = ~(input_a[26] & input_a[7]);
  assign popcount28_elja_core_098 = ~(input_a[18] ^ input_a[10]);
  assign popcount28_elja_core_100 = input_a[1] | input_a[7];
  assign popcount28_elja_core_102 = input_a[16] ^ input_a[6];
  assign popcount28_elja_core_103 = ~(input_a[14] | input_a[6]);
  assign popcount28_elja_core_104 = ~(input_a[12] ^ input_a[17]);
  assign popcount28_elja_core_105 = ~(input_a[5] | input_a[16]);
  assign popcount28_elja_core_107 = ~(input_a[4] ^ input_a[23]);
  assign popcount28_elja_core_110 = ~(input_a[26] | input_a[20]);
  assign popcount28_elja_core_112 = ~(input_a[20] | input_a[2]);
  assign popcount28_elja_core_113 = ~(input_a[3] | input_a[9]);
  assign popcount28_elja_core_114 = input_a[12] & input_a[22];
  assign popcount28_elja_core_115 = input_a[24] ^ input_a[19];
  assign popcount28_elja_core_116 = ~input_a[1];
  assign popcount28_elja_core_117 = ~(input_a[18] & input_a[15]);
  assign popcount28_elja_core_118 = input_a[23] ^ input_a[5];
  assign popcount28_elja_core_119 = input_a[4] | input_a[1];
  assign popcount28_elja_core_120 = ~(input_a[14] | input_a[14]);
  assign popcount28_elja_core_121 = input_a[8] | input_a[27];
  assign popcount28_elja_core_123 = ~(input_a[6] ^ input_a[20]);
  assign popcount28_elja_core_124 = ~(input_a[18] | input_a[2]);
  assign popcount28_elja_core_125 = ~(input_a[13] | input_a[1]);
  assign popcount28_elja_core_128 = ~(input_a[8] & input_a[10]);
  assign popcount28_elja_core_129 = input_a[19] | input_a[12];
  assign popcount28_elja_core_130 = ~(input_a[2] | input_a[20]);
  assign popcount28_elja_core_131 = input_a[5] & input_a[14];
  assign popcount28_elja_core_132 = ~input_a[26];
  assign popcount28_elja_core_134 = ~input_a[3];
  assign popcount28_elja_core_135 = input_a[3] | input_a[10];
  assign popcount28_elja_core_136_not = ~input_a[21];
  assign popcount28_elja_core_138_not = ~input_a[24];
  assign popcount28_elja_core_139 = input_a[22] ^ input_a[18];
  assign popcount28_elja_core_141 = ~(input_a[5] & input_a[2]);
  assign popcount28_elja_core_142 = ~input_a[9];
  assign popcount28_elja_core_144 = ~input_a[20];
  assign popcount28_elja_core_145 = input_a[0] | input_a[23];
  assign popcount28_elja_core_146 = ~input_a[17];
  assign popcount28_elja_core_147 = ~input_a[14];
  assign popcount28_elja_core_148 = ~input_a[13];
  assign popcount28_elja_core_149 = ~(input_a[2] & input_a[1]);
  assign popcount28_elja_core_150 = ~input_a[17];
  assign popcount28_elja_core_151 = ~(input_a[19] ^ input_a[8]);
  assign popcount28_elja_core_153 = input_a[13] ^ input_a[8];
  assign popcount28_elja_core_154 = ~input_a[9];
  assign popcount28_elja_core_158 = ~(input_a[22] | input_a[27]);
  assign popcount28_elja_core_160 = input_a[21] & input_a[20];
  assign popcount28_elja_core_163 = ~(input_a[23] ^ input_a[17]);
  assign popcount28_elja_core_165 = input_a[14] | input_a[27];
  assign popcount28_elja_core_167 = ~(input_a[9] ^ input_a[24]);
  assign popcount28_elja_core_168 = ~(input_a[17] & input_a[23]);
  assign popcount28_elja_core_170 = ~(input_a[5] & input_a[0]);
  assign popcount28_elja_core_171 = ~(input_a[20] | input_a[5]);
  assign popcount28_elja_core_174 = ~(input_a[20] ^ input_a[22]);
  assign popcount28_elja_core_175 = ~(input_a[16] & input_a[16]);
  assign popcount28_elja_core_176 = input_a[10] ^ input_a[2];
  assign popcount28_elja_core_177 = ~input_a[18];
  assign popcount28_elja_core_178 = ~(input_a[22] | input_a[14]);
  assign popcount28_elja_core_179 = ~(input_a[13] & input_a[9]);
  assign popcount28_elja_core_180 = ~(input_a[19] ^ input_a[26]);
  assign popcount28_elja_core_183 = ~(input_a[24] & input_a[15]);
  assign popcount28_elja_core_184 = ~input_a[25];
  assign popcount28_elja_core_188 = input_a[16] & input_a[25];
  assign popcount28_elja_core_190 = input_a[25] & input_a[6];
  assign popcount28_elja_core_191 = input_a[21] ^ input_a[15];
  assign popcount28_elja_core_192 = ~(input_a[20] & input_a[22]);
  assign popcount28_elja_core_194 = input_a[19] | input_a[11];
  assign popcount28_elja_core_197_not = ~input_a[24];
  assign popcount28_elja_core_199 = ~(input_a[20] | input_a[1]);
  assign popcount28_elja_core_200 = input_a[22] ^ input_a[15];

  assign popcount28_elja_out[0] = input_a[15];
  assign popcount28_elja_out[1] = input_a[11];
  assign popcount28_elja_out[2] = input_a[3];
  assign popcount28_elja_out[3] = input_a[20];
  assign popcount28_elja_out[4] = 1'b0;
endmodule