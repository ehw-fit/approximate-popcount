// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=1.52052
// WCE=6.0
// EP=0.801678%
// Printed PDK parameters:
//  Area=46227717.0
//  Delay=68233896.0
//  Power=2502500.0

module popcount29_2bwi(input [28:0] input_a, output [4:0] popcount29_2bwi_out);
  wire popcount29_2bwi_core_032;
  wire popcount29_2bwi_core_034;
  wire popcount29_2bwi_core_037;
  wire popcount29_2bwi_core_038;
  wire popcount29_2bwi_core_039;
  wire popcount29_2bwi_core_040;
  wire popcount29_2bwi_core_041;
  wire popcount29_2bwi_core_042;
  wire popcount29_2bwi_core_043;
  wire popcount29_2bwi_core_044;
  wire popcount29_2bwi_core_045;
  wire popcount29_2bwi_core_046;
  wire popcount29_2bwi_core_047;
  wire popcount29_2bwi_core_048;
  wire popcount29_2bwi_core_050;
  wire popcount29_2bwi_core_051;
  wire popcount29_2bwi_core_053;
  wire popcount29_2bwi_core_056;
  wire popcount29_2bwi_core_057;
  wire popcount29_2bwi_core_059;
  wire popcount29_2bwi_core_060;
  wire popcount29_2bwi_core_062;
  wire popcount29_2bwi_core_063;
  wire popcount29_2bwi_core_065;
  wire popcount29_2bwi_core_066;
  wire popcount29_2bwi_core_067;
  wire popcount29_2bwi_core_069;
  wire popcount29_2bwi_core_070;
  wire popcount29_2bwi_core_071;
  wire popcount29_2bwi_core_073;
  wire popcount29_2bwi_core_074;
  wire popcount29_2bwi_core_076;
  wire popcount29_2bwi_core_077;
  wire popcount29_2bwi_core_079;
  wire popcount29_2bwi_core_084;
  wire popcount29_2bwi_core_085;
  wire popcount29_2bwi_core_086;
  wire popcount29_2bwi_core_088;
  wire popcount29_2bwi_core_089;
  wire popcount29_2bwi_core_091;
  wire popcount29_2bwi_core_093;
  wire popcount29_2bwi_core_094_not;
  wire popcount29_2bwi_core_098;
  wire popcount29_2bwi_core_102;
  wire popcount29_2bwi_core_104;
  wire popcount29_2bwi_core_105;
  wire popcount29_2bwi_core_108;
  wire popcount29_2bwi_core_109;
  wire popcount29_2bwi_core_113;
  wire popcount29_2bwi_core_114;
  wire popcount29_2bwi_core_115;
  wire popcount29_2bwi_core_116;
  wire popcount29_2bwi_core_117;
  wire popcount29_2bwi_core_118;
  wire popcount29_2bwi_core_119;
  wire popcount29_2bwi_core_124;
  wire popcount29_2bwi_core_125;
  wire popcount29_2bwi_core_126;
  wire popcount29_2bwi_core_127;
  wire popcount29_2bwi_core_128;
  wire popcount29_2bwi_core_129;
  wire popcount29_2bwi_core_131;
  wire popcount29_2bwi_core_132;
  wire popcount29_2bwi_core_135;
  wire popcount29_2bwi_core_136;
  wire popcount29_2bwi_core_137;
  wire popcount29_2bwi_core_138;
  wire popcount29_2bwi_core_139;
  wire popcount29_2bwi_core_140;
  wire popcount29_2bwi_core_141;
  wire popcount29_2bwi_core_142;
  wire popcount29_2bwi_core_143;
  wire popcount29_2bwi_core_144;
  wire popcount29_2bwi_core_146;
  wire popcount29_2bwi_core_147;
  wire popcount29_2bwi_core_148;
  wire popcount29_2bwi_core_149;
  wire popcount29_2bwi_core_150;
  wire popcount29_2bwi_core_151;
  wire popcount29_2bwi_core_152;
  wire popcount29_2bwi_core_153;
  wire popcount29_2bwi_core_154;
  wire popcount29_2bwi_core_155;
  wire popcount29_2bwi_core_157;
  wire popcount29_2bwi_core_158;
  wire popcount29_2bwi_core_159;
  wire popcount29_2bwi_core_160;
  wire popcount29_2bwi_core_161;
  wire popcount29_2bwi_core_162;
  wire popcount29_2bwi_core_163;
  wire popcount29_2bwi_core_164;
  wire popcount29_2bwi_core_165;
  wire popcount29_2bwi_core_166;
  wire popcount29_2bwi_core_167;
  wire popcount29_2bwi_core_169;
  wire popcount29_2bwi_core_170;
  wire popcount29_2bwi_core_171;
  wire popcount29_2bwi_core_172;
  wire popcount29_2bwi_core_173;
  wire popcount29_2bwi_core_174;
  wire popcount29_2bwi_core_175;
  wire popcount29_2bwi_core_176;
  wire popcount29_2bwi_core_177;
  wire popcount29_2bwi_core_178;
  wire popcount29_2bwi_core_179;
  wire popcount29_2bwi_core_180;
  wire popcount29_2bwi_core_183;
  wire popcount29_2bwi_core_184_not;
  wire popcount29_2bwi_core_186;
  wire popcount29_2bwi_core_187;
  wire popcount29_2bwi_core_188;
  wire popcount29_2bwi_core_189;
  wire popcount29_2bwi_core_190;
  wire popcount29_2bwi_core_191;
  wire popcount29_2bwi_core_192;
  wire popcount29_2bwi_core_193;
  wire popcount29_2bwi_core_194;
  wire popcount29_2bwi_core_195;
  wire popcount29_2bwi_core_196;
  wire popcount29_2bwi_core_197;
  wire popcount29_2bwi_core_198;
  wire popcount29_2bwi_core_199;
  wire popcount29_2bwi_core_200;
  wire popcount29_2bwi_core_201;
  wire popcount29_2bwi_core_202;
  wire popcount29_2bwi_core_203;
  wire popcount29_2bwi_core_204;
  wire popcount29_2bwi_core_205;
  wire popcount29_2bwi_core_206;
  wire popcount29_2bwi_core_207;

  assign popcount29_2bwi_core_032 = input_a[3] & input_a[1];
  assign popcount29_2bwi_core_034 = input_a[26] ^ input_a[4];
  assign popcount29_2bwi_core_037 = input_a[11] ^ input_a[3];
  assign popcount29_2bwi_core_038 = input_a[0] & input_a[13];
  assign popcount29_2bwi_core_039 = ~input_a[25];
  assign popcount29_2bwi_core_040 = input_a[9] & input_a[10];
  assign popcount29_2bwi_core_041 = input_a[22] | input_a[28];
  assign popcount29_2bwi_core_042 = input_a[19] & input_a[12];
  assign popcount29_2bwi_core_043 = popcount29_2bwi_core_038 | popcount29_2bwi_core_040;
  assign popcount29_2bwi_core_044 = popcount29_2bwi_core_038 & popcount29_2bwi_core_040;
  assign popcount29_2bwi_core_045 = popcount29_2bwi_core_043 | popcount29_2bwi_core_042;
  assign popcount29_2bwi_core_046 = popcount29_2bwi_core_043 & popcount29_2bwi_core_042;
  assign popcount29_2bwi_core_047 = popcount29_2bwi_core_044 | popcount29_2bwi_core_046;
  assign popcount29_2bwi_core_048 = ~(input_a[15] | input_a[28]);
  assign popcount29_2bwi_core_050 = ~input_a[12];
  assign popcount29_2bwi_core_051 = popcount29_2bwi_core_032 & popcount29_2bwi_core_045;
  assign popcount29_2bwi_core_053 = ~(input_a[14] & input_a[19]);
  assign popcount29_2bwi_core_056 = ~(input_a[28] ^ input_a[8]);
  assign popcount29_2bwi_core_057 = popcount29_2bwi_core_047 | popcount29_2bwi_core_051;
  assign popcount29_2bwi_core_059 = ~(input_a[2] & input_a[26]);
  assign popcount29_2bwi_core_060 = ~input_a[20];
  assign popcount29_2bwi_core_062 = ~(input_a[10] ^ input_a[26]);
  assign popcount29_2bwi_core_063 = input_a[15] ^ input_a[22];
  assign popcount29_2bwi_core_065 = ~(input_a[28] | input_a[9]);
  assign popcount29_2bwi_core_066 = ~(input_a[19] ^ input_a[14]);
  assign popcount29_2bwi_core_067 = ~(input_a[24] & input_a[18]);
  assign popcount29_2bwi_core_069 = ~(input_a[19] & input_a[10]);
  assign popcount29_2bwi_core_070 = ~input_a[12];
  assign popcount29_2bwi_core_071 = ~(input_a[18] ^ input_a[25]);
  assign popcount29_2bwi_core_073 = ~(input_a[24] & input_a[6]);
  assign popcount29_2bwi_core_074 = ~(input_a[27] | input_a[28]);
  assign popcount29_2bwi_core_076 = input_a[15] & input_a[20];
  assign popcount29_2bwi_core_077 = ~(input_a[27] & input_a[17]);
  assign popcount29_2bwi_core_079 = input_a[10] ^ input_a[17];
  assign popcount29_2bwi_core_084 = ~(input_a[16] & input_a[4]);
  assign popcount29_2bwi_core_085 = ~(input_a[18] ^ input_a[12]);
  assign popcount29_2bwi_core_086 = input_a[15] | input_a[23];
  assign popcount29_2bwi_core_088 = input_a[21] ^ input_a[25];
  assign popcount29_2bwi_core_089 = input_a[18] & input_a[10];
  assign popcount29_2bwi_core_091 = input_a[21] ^ input_a[21];
  assign popcount29_2bwi_core_093 = input_a[4] | input_a[7];
  assign popcount29_2bwi_core_094_not = ~input_a[2];
  assign popcount29_2bwi_core_098 = ~popcount29_2bwi_core_057;
  assign popcount29_2bwi_core_102 = ~(input_a[10] & input_a[7]);
  assign popcount29_2bwi_core_104 = ~(input_a[25] & input_a[15]);
  assign popcount29_2bwi_core_105 = ~(input_a[16] & input_a[25]);
  assign popcount29_2bwi_core_108 = ~(input_a[3] ^ input_a[22]);
  assign popcount29_2bwi_core_109 = input_a[14] & input_a[6];
  assign popcount29_2bwi_core_113 = input_a[16] & input_a[18];
  assign popcount29_2bwi_core_114 = input_a[1] ^ input_a[1];
  assign popcount29_2bwi_core_115 = input_a[15] & input_a[20];
  assign popcount29_2bwi_core_116 = ~(input_a[16] | input_a[0]);
  assign popcount29_2bwi_core_117 = ~(input_a[23] ^ input_a[27]);
  assign popcount29_2bwi_core_118 = popcount29_2bwi_core_113 ^ popcount29_2bwi_core_115;
  assign popcount29_2bwi_core_119 = popcount29_2bwi_core_113 & popcount29_2bwi_core_115;
  assign popcount29_2bwi_core_124 = input_a[8] & input_a[17];
  assign popcount29_2bwi_core_125 = popcount29_2bwi_core_109 ^ popcount29_2bwi_core_118;
  assign popcount29_2bwi_core_126 = popcount29_2bwi_core_109 & popcount29_2bwi_core_118;
  assign popcount29_2bwi_core_127 = popcount29_2bwi_core_125 ^ popcount29_2bwi_core_124;
  assign popcount29_2bwi_core_128 = popcount29_2bwi_core_125 & popcount29_2bwi_core_124;
  assign popcount29_2bwi_core_129 = popcount29_2bwi_core_126 | popcount29_2bwi_core_128;
  assign popcount29_2bwi_core_131 = ~(input_a[17] ^ input_a[16]);
  assign popcount29_2bwi_core_132 = popcount29_2bwi_core_119 | popcount29_2bwi_core_129;
  assign popcount29_2bwi_core_135 = input_a[21] ^ input_a[22];
  assign popcount29_2bwi_core_136 = input_a[21] & input_a[22];
  assign popcount29_2bwi_core_137 = input_a[23] ^ input_a[24];
  assign popcount29_2bwi_core_138 = input_a[23] & input_a[24];
  assign popcount29_2bwi_core_139 = popcount29_2bwi_core_135 ^ popcount29_2bwi_core_137;
  assign popcount29_2bwi_core_140 = popcount29_2bwi_core_135 & popcount29_2bwi_core_137;
  assign popcount29_2bwi_core_141 = popcount29_2bwi_core_136 ^ popcount29_2bwi_core_138;
  assign popcount29_2bwi_core_142 = popcount29_2bwi_core_136 & popcount29_2bwi_core_138;
  assign popcount29_2bwi_core_143 = popcount29_2bwi_core_141 | popcount29_2bwi_core_140;
  assign popcount29_2bwi_core_144 = ~(input_a[23] ^ input_a[21]);
  assign popcount29_2bwi_core_146 = input_a[25] ^ input_a[26];
  assign popcount29_2bwi_core_147 = input_a[25] & input_a[26];
  assign popcount29_2bwi_core_148 = input_a[27] ^ input_a[28];
  assign popcount29_2bwi_core_149 = input_a[27] & input_a[28];
  assign popcount29_2bwi_core_150 = popcount29_2bwi_core_146 ^ popcount29_2bwi_core_148;
  assign popcount29_2bwi_core_151 = popcount29_2bwi_core_146 & popcount29_2bwi_core_148;
  assign popcount29_2bwi_core_152 = popcount29_2bwi_core_147 ^ popcount29_2bwi_core_149;
  assign popcount29_2bwi_core_153 = popcount29_2bwi_core_147 & popcount29_2bwi_core_149;
  assign popcount29_2bwi_core_154 = popcount29_2bwi_core_152 | popcount29_2bwi_core_151;
  assign popcount29_2bwi_core_155 = ~(input_a[17] & input_a[0]);
  assign popcount29_2bwi_core_157 = popcount29_2bwi_core_139 ^ popcount29_2bwi_core_150;
  assign popcount29_2bwi_core_158 = popcount29_2bwi_core_139 & popcount29_2bwi_core_150;
  assign popcount29_2bwi_core_159 = popcount29_2bwi_core_143 ^ popcount29_2bwi_core_154;
  assign popcount29_2bwi_core_160 = popcount29_2bwi_core_143 & popcount29_2bwi_core_154;
  assign popcount29_2bwi_core_161 = popcount29_2bwi_core_159 ^ popcount29_2bwi_core_158;
  assign popcount29_2bwi_core_162 = popcount29_2bwi_core_159 & popcount29_2bwi_core_158;
  assign popcount29_2bwi_core_163 = popcount29_2bwi_core_160 | popcount29_2bwi_core_162;
  assign popcount29_2bwi_core_164 = popcount29_2bwi_core_142 ^ popcount29_2bwi_core_153;
  assign popcount29_2bwi_core_165 = popcount29_2bwi_core_142 & popcount29_2bwi_core_153;
  assign popcount29_2bwi_core_166 = popcount29_2bwi_core_164 | popcount29_2bwi_core_163;
  assign popcount29_2bwi_core_167 = ~(input_a[2] ^ input_a[19]);
  assign popcount29_2bwi_core_169 = input_a[1] | input_a[2];
  assign popcount29_2bwi_core_170 = input_a[2] & popcount29_2bwi_core_157;
  assign popcount29_2bwi_core_171 = popcount29_2bwi_core_127 ^ popcount29_2bwi_core_161;
  assign popcount29_2bwi_core_172 = popcount29_2bwi_core_127 & popcount29_2bwi_core_161;
  assign popcount29_2bwi_core_173 = popcount29_2bwi_core_171 ^ popcount29_2bwi_core_170;
  assign popcount29_2bwi_core_174 = popcount29_2bwi_core_171 & popcount29_2bwi_core_170;
  assign popcount29_2bwi_core_175 = popcount29_2bwi_core_172 | popcount29_2bwi_core_174;
  assign popcount29_2bwi_core_176 = popcount29_2bwi_core_132 ^ popcount29_2bwi_core_166;
  assign popcount29_2bwi_core_177 = popcount29_2bwi_core_132 & popcount29_2bwi_core_166;
  assign popcount29_2bwi_core_178 = popcount29_2bwi_core_176 ^ popcount29_2bwi_core_175;
  assign popcount29_2bwi_core_179 = popcount29_2bwi_core_176 & popcount29_2bwi_core_175;
  assign popcount29_2bwi_core_180 = popcount29_2bwi_core_177 | popcount29_2bwi_core_179;
  assign popcount29_2bwi_core_183 = popcount29_2bwi_core_165 | popcount29_2bwi_core_180;
  assign popcount29_2bwi_core_184_not = ~input_a[22];
  assign popcount29_2bwi_core_186 = ~(input_a[17] | input_a[24]);
  assign popcount29_2bwi_core_187 = ~(input_a[13] | input_a[11]);
  assign popcount29_2bwi_core_188 = popcount29_2bwi_core_093 ^ popcount29_2bwi_core_173;
  assign popcount29_2bwi_core_189 = popcount29_2bwi_core_093 & popcount29_2bwi_core_173;
  assign popcount29_2bwi_core_190 = popcount29_2bwi_core_188 ^ input_a[11];
  assign popcount29_2bwi_core_191 = popcount29_2bwi_core_188 & input_a[11];
  assign popcount29_2bwi_core_192 = popcount29_2bwi_core_189 | popcount29_2bwi_core_191;
  assign popcount29_2bwi_core_193 = popcount29_2bwi_core_098 ^ popcount29_2bwi_core_178;
  assign popcount29_2bwi_core_194 = popcount29_2bwi_core_098 & popcount29_2bwi_core_178;
  assign popcount29_2bwi_core_195 = popcount29_2bwi_core_193 ^ popcount29_2bwi_core_192;
  assign popcount29_2bwi_core_196 = popcount29_2bwi_core_193 & popcount29_2bwi_core_192;
  assign popcount29_2bwi_core_197 = popcount29_2bwi_core_194 | popcount29_2bwi_core_196;
  assign popcount29_2bwi_core_198 = popcount29_2bwi_core_057 ^ popcount29_2bwi_core_183;
  assign popcount29_2bwi_core_199 = popcount29_2bwi_core_057 & popcount29_2bwi_core_183;
  assign popcount29_2bwi_core_200 = popcount29_2bwi_core_198 ^ popcount29_2bwi_core_197;
  assign popcount29_2bwi_core_201 = popcount29_2bwi_core_198 & popcount29_2bwi_core_197;
  assign popcount29_2bwi_core_202 = popcount29_2bwi_core_199 | popcount29_2bwi_core_201;
  assign popcount29_2bwi_core_203 = input_a[25] ^ input_a[19];
  assign popcount29_2bwi_core_204 = ~input_a[7];
  assign popcount29_2bwi_core_205 = ~(input_a[9] ^ input_a[16]);
  assign popcount29_2bwi_core_206 = input_a[4] ^ input_a[5];
  assign popcount29_2bwi_core_207 = ~(input_a[13] ^ input_a[12]);

  assign popcount29_2bwi_out[0] = input_a[5];
  assign popcount29_2bwi_out[1] = popcount29_2bwi_core_190;
  assign popcount29_2bwi_out[2] = popcount29_2bwi_core_195;
  assign popcount29_2bwi_out[3] = popcount29_2bwi_core_200;
  assign popcount29_2bwi_out[4] = popcount29_2bwi_core_202;
endmodule