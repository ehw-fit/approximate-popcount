
module cmp_pos(input [46:0] input_a, output [5:0] cgp_out);
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_059;
  wire cgp_core_060;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_065;
  wire cgp_core_066;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_071;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_081;
  wire cgp_core_082;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_086;
  wire cgp_core_088;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_094;
  wire cgp_core_095;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_099;
  wire cgp_core_100;
  wire cgp_core_101;
  wire cgp_core_103;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_111;
  wire cgp_core_113;
  wire cgp_core_114;
  wire cgp_core_115;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_119;
  wire cgp_core_120;
  wire cgp_core_121;
  wire cgp_core_122;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_127;
  wire cgp_core_129;
  wire cgp_core_130;
  wire cgp_core_131;
  wire cgp_core_132;
  wire cgp_core_133;
  wire cgp_core_134;
  wire cgp_core_135;
  wire cgp_core_136;
  wire cgp_core_137;
  wire cgp_core_138;
  wire cgp_core_139;
  wire cgp_core_140;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_146;
  wire cgp_core_147;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_158;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_161;
  wire cgp_core_162;
  wire cgp_core_163;
  wire cgp_core_164;
  wire cgp_core_165;
  wire cgp_core_166;
  wire cgp_core_170;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_174;
  wire cgp_core_175;
  wire cgp_core_176;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_180;
  wire cgp_core_181;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_187;
  wire cgp_core_188;
  wire cgp_core_192;
  wire cgp_core_193;
  wire cgp_core_194;
  wire cgp_core_195;
  wire cgp_core_196;
  wire cgp_core_197;
  wire cgp_core_198;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_203;
  wire cgp_core_204;
  wire cgp_core_206;
  wire cgp_core_207;
  wire cgp_core_208;
  wire cgp_core_209;
  wire cgp_core_210;
  wire cgp_core_211;
  wire cgp_core_212;
  wire cgp_core_216;
  wire cgp_core_217;
  wire cgp_core_218;
  wire cgp_core_219;
  wire cgp_core_220;
  wire cgp_core_221;
  wire cgp_core_222;
  wire cgp_core_223;
  wire cgp_core_224;
  wire cgp_core_225;
  wire cgp_core_226;
  wire cgp_core_227;
  wire cgp_core_228;
  wire cgp_core_229;
  wire cgp_core_230;
  wire cgp_core_231;
  wire cgp_core_232;
  wire cgp_core_233;
  wire cgp_core_234;
  wire cgp_core_235;
  wire cgp_core_236;
  wire cgp_core_240;
  wire cgp_core_242;
  wire cgp_core_243;
  wire cgp_core_244;
  wire cgp_core_245;
  wire cgp_core_246;
  wire cgp_core_247;
  wire cgp_core_248;
  wire cgp_core_249;
  wire cgp_core_250;
  wire cgp_core_251;
  wire cgp_core_252;
  wire cgp_core_253;
  wire cgp_core_255;
  wire cgp_core_257;
  wire cgp_core_258;
  wire cgp_core_259;
  wire cgp_core_260;
  wire cgp_core_261;
  wire cgp_core_262;
  wire cgp_core_263;
  wire cgp_core_265;
  wire cgp_core_266;
  wire cgp_core_267;
  wire cgp_core_268;
  wire cgp_core_269;
  wire cgp_core_272;
  wire cgp_core_273;
  wire cgp_core_274;
  wire cgp_core_276;
  wire cgp_core_279;
  wire cgp_core_281;
  wire cgp_core_282;
  wire cgp_core_283;
  wire cgp_core_284;
  wire cgp_core_285;
  wire cgp_core_286;
  wire cgp_core_287;
  wire cgp_core_288;
  wire cgp_core_289;
  wire cgp_core_290;
  wire cgp_core_291;
  wire cgp_core_292;
  wire cgp_core_293;
  wire cgp_core_294;
  wire cgp_core_295;
  wire cgp_core_296;
  wire cgp_core_297;
  wire cgp_core_298;
  wire cgp_core_299;
  wire cgp_core_300;
  wire cgp_core_301;
  wire cgp_core_303;
  wire cgp_core_305;
  wire cgp_core_306;
  wire cgp_core_307;
  wire cgp_core_309;
  wire cgp_core_310;
  wire cgp_core_311;
  wire cgp_core_312;
  wire cgp_core_313;
  wire cgp_core_314;
  wire cgp_core_315;
  wire cgp_core_316;
  wire cgp_core_317;
  wire cgp_core_318;
  wire cgp_core_320;
  wire cgp_core_324;
  wire cgp_core_325;
  wire cgp_core_326;
  wire cgp_core_327;
  wire cgp_core_328;
  wire cgp_core_329;
  wire cgp_core_330;
  wire cgp_core_331;
  wire cgp_core_332;
  wire cgp_core_333;
  wire cgp_core_334;
  wire cgp_core_335;
  wire cgp_core_336;
  wire cgp_core_337;
  wire cgp_core_338;
  wire cgp_core_339;
  wire cgp_core_340;
  wire cgp_core_345;
  wire cgp_core_346;
  wire cgp_core_347;
  wire cgp_core_348;
  wire cgp_core_349;
  wire cgp_core_350;
  wire cgp_core_351;
  wire cgp_core_352;
  wire cgp_core_353;
  wire cgp_core_354;
  wire cgp_core_355;
  wire cgp_core_356;
  wire cgp_core_357;
  wire cgp_core_358;
  wire cgp_core_359;
  wire cgp_core_360;
  wire cgp_core_361;
  wire cgp_core_362;
  wire cgp_core_363;
  wire cgp_core_364;
  wire cgp_core_365;
  wire cgp_core_366;
  wire cgp_core_367;
  wire cgp_core_369;
  wire cgp_core_370;

  assign cgp_core_049 = input_a[0] ^ input_a[1];
  assign cgp_core_050 = input_a[0] & input_a[1];
  assign cgp_core_051 = input_a[3] ^ input_a[4];
  assign cgp_core_052 = input_a[3] & input_a[4];
  assign cgp_core_053 = input_a[2] ^ cgp_core_051;
  assign cgp_core_054 = input_a[2] & cgp_core_051;
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_057 = cgp_core_049 ^ cgp_core_053;
  assign cgp_core_058 = cgp_core_049 & cgp_core_053;
  assign cgp_core_059 = cgp_core_050 ^ cgp_core_055;
  assign cgp_core_060 = cgp_core_050 & cgp_core_055;
  assign cgp_core_061 = cgp_core_059 ^ cgp_core_058;
  assign cgp_core_062 = cgp_core_059 & cgp_core_058;
  assign cgp_core_063 = cgp_core_060 | cgp_core_062;
  assign cgp_core_065 = input_a[20] & input_a[32];
  assign cgp_core_066 = input_a[6] ^ input_a[7];
  assign cgp_core_067 = input_a[6] & input_a[7];
  assign cgp_core_068 = input_a[5] ^ cgp_core_066;
  assign cgp_core_069 = input_a[5] & cgp_core_066;
  assign cgp_core_070 = cgp_core_067 | cgp_core_069;
  assign cgp_core_071 = input_a[44] | input_a[23];
  assign cgp_core_072 = input_a[9] ^ input_a[10];
  assign cgp_core_073 = input_a[9] & input_a[10];
  assign cgp_core_074 = input_a[8] ^ cgp_core_072;
  assign cgp_core_075 = input_a[8] & cgp_core_072;
  assign cgp_core_076 = cgp_core_073 | cgp_core_075;
  assign cgp_core_077 = input_a[46] ^ input_a[4];
  assign cgp_core_078 = cgp_core_068 ^ cgp_core_074;
  assign cgp_core_079 = cgp_core_068 & cgp_core_074;
  assign cgp_core_080 = cgp_core_070 ^ cgp_core_076;
  assign cgp_core_081 = cgp_core_070 & cgp_core_076;
  assign cgp_core_082 = cgp_core_080 ^ cgp_core_079;
  assign cgp_core_083 = cgp_core_080 & cgp_core_079;
  assign cgp_core_084 = cgp_core_081 | cgp_core_083;
  assign cgp_core_086 = ~input_a[36];
  assign cgp_core_088 = input_a[43] & input_a[4];
  assign cgp_core_090 = cgp_core_057 ^ cgp_core_078;
  assign cgp_core_091 = cgp_core_057 & cgp_core_078;
  assign cgp_core_092 = cgp_core_061 ^ cgp_core_082;
  assign cgp_core_093 = cgp_core_061 & cgp_core_082;
  assign cgp_core_094 = cgp_core_092 ^ cgp_core_091;
  assign cgp_core_095 = cgp_core_092 & cgp_core_091;
  assign cgp_core_096 = cgp_core_093 | cgp_core_095;
  assign cgp_core_097 = cgp_core_063 ^ cgp_core_084;
  assign cgp_core_098 = cgp_core_063 & cgp_core_084;
  assign cgp_core_099 = cgp_core_097 ^ cgp_core_096;
  assign cgp_core_100 = cgp_core_097 & cgp_core_096;
  assign cgp_core_101 = cgp_core_098 | cgp_core_100;
  assign cgp_core_103 = ~(input_a[17] ^ input_a[4]);
  assign cgp_core_107 = input_a[12] ^ input_a[13];
  assign cgp_core_108 = input_a[12] & input_a[13];
  assign cgp_core_109 = input_a[11] ^ cgp_core_107;
  assign cgp_core_110 = input_a[11] & cgp_core_107;
  assign cgp_core_111 = cgp_core_108 | cgp_core_110;
  assign cgp_core_113 = input_a[15] ^ input_a[16];
  assign cgp_core_114 = input_a[15] & input_a[16];
  assign cgp_core_115 = input_a[14] ^ cgp_core_113;
  assign cgp_core_116 = input_a[14] & cgp_core_113;
  assign cgp_core_117 = cgp_core_114 | cgp_core_116;
  assign cgp_core_119 = cgp_core_109 ^ cgp_core_115;
  assign cgp_core_120 = cgp_core_109 & cgp_core_115;
  assign cgp_core_121 = cgp_core_111 ^ cgp_core_117;
  assign cgp_core_122 = cgp_core_111 & cgp_core_117;
  assign cgp_core_123 = cgp_core_121 ^ cgp_core_120;
  assign cgp_core_124 = cgp_core_121 & cgp_core_120;
  assign cgp_core_125 = cgp_core_122 | cgp_core_124;
  assign cgp_core_127 = input_a[5] ^ input_a[32];
  assign cgp_core_129 = input_a[11] ^ input_a[9];
  assign cgp_core_130 = ~input_a[35];
  assign cgp_core_131 = input_a[18] ^ input_a[19];
  assign cgp_core_132 = input_a[18] & input_a[19];
  assign cgp_core_133 = input_a[17] ^ cgp_core_131;
  assign cgp_core_134 = input_a[17] & cgp_core_131;
  assign cgp_core_135 = cgp_core_132 | cgp_core_134;
  assign cgp_core_136 = ~(input_a[1] ^ input_a[9]);
  assign cgp_core_137 = input_a[21] ^ input_a[22];
  assign cgp_core_138 = input_a[21] & input_a[22];
  assign cgp_core_139 = input_a[20] ^ cgp_core_137;
  assign cgp_core_140 = input_a[20] & cgp_core_137;
  assign cgp_core_141 = cgp_core_138 | cgp_core_140;
  assign cgp_core_142 = ~(input_a[25] & input_a[42]);
  assign cgp_core_143 = cgp_core_133 ^ cgp_core_139;
  assign cgp_core_144 = cgp_core_133 & cgp_core_139;
  assign cgp_core_145 = cgp_core_135 ^ cgp_core_141;
  assign cgp_core_146 = cgp_core_135 & cgp_core_141;
  assign cgp_core_147 = cgp_core_145 ^ cgp_core_144;
  assign cgp_core_148 = cgp_core_145 & cgp_core_144;
  assign cgp_core_149 = cgp_core_146 | cgp_core_148;
  assign cgp_core_153 = input_a[25] ^ input_a[42];
  assign cgp_core_154 = input_a[28] | input_a[8];
  assign cgp_core_155 = cgp_core_119 ^ cgp_core_143;
  assign cgp_core_156 = cgp_core_119 & cgp_core_143;
  assign cgp_core_157 = cgp_core_123 ^ cgp_core_147;
  assign cgp_core_158 = cgp_core_123 & cgp_core_147;
  assign cgp_core_159 = cgp_core_157 ^ cgp_core_156;
  assign cgp_core_160 = cgp_core_157 & cgp_core_156;
  assign cgp_core_161 = cgp_core_158 | cgp_core_160;
  assign cgp_core_162 = cgp_core_125 ^ cgp_core_149;
  assign cgp_core_163 = cgp_core_125 & cgp_core_149;
  assign cgp_core_164 = cgp_core_162 ^ cgp_core_161;
  assign cgp_core_165 = cgp_core_162 & cgp_core_161;
  assign cgp_core_166 = cgp_core_163 | cgp_core_165;
  assign cgp_core_170 = ~(input_a[38] & input_a[15]);
  assign cgp_core_172 = cgp_core_090 ^ cgp_core_155;
  assign cgp_core_173 = cgp_core_090 & cgp_core_155;
  assign cgp_core_174 = cgp_core_094 ^ cgp_core_159;
  assign cgp_core_175 = cgp_core_094 & cgp_core_159;
  assign cgp_core_176 = cgp_core_174 ^ cgp_core_173;
  assign cgp_core_177 = cgp_core_174 & cgp_core_173;
  assign cgp_core_178 = cgp_core_175 | cgp_core_177;
  assign cgp_core_179 = cgp_core_099 ^ cgp_core_164;
  assign cgp_core_180 = cgp_core_099 & cgp_core_164;
  assign cgp_core_181 = cgp_core_179 ^ cgp_core_178;
  assign cgp_core_182 = cgp_core_179 & cgp_core_178;
  assign cgp_core_183 = cgp_core_180 | cgp_core_182;
  assign cgp_core_184 = cgp_core_101 ^ cgp_core_166;
  assign cgp_core_185 = cgp_core_101 & cgp_core_166;
  assign cgp_core_186 = cgp_core_184 ^ cgp_core_183;
  assign cgp_core_187 = cgp_core_184 & cgp_core_183;
  assign cgp_core_188 = cgp_core_185 | cgp_core_187;
  assign cgp_core_192 = ~input_a[19];
  assign cgp_core_193 = ~input_a[36];
  assign cgp_core_194 = input_a[24] ^ input_a[25];
  assign cgp_core_195 = input_a[24] & input_a[25];
  assign cgp_core_196 = input_a[23] ^ cgp_core_194;
  assign cgp_core_197 = input_a[23] & cgp_core_194;
  assign cgp_core_198 = cgp_core_195 | cgp_core_197;
  assign cgp_core_199 = ~(input_a[45] & input_a[28]);
  assign cgp_core_200 = input_a[27] ^ input_a[28];
  assign cgp_core_201 = input_a[27] & input_a[28];
  assign cgp_core_202 = input_a[26] ^ cgp_core_200;
  assign cgp_core_203 = input_a[26] & cgp_core_200;
  assign cgp_core_204 = cgp_core_201 | cgp_core_203;
  assign cgp_core_206 = cgp_core_196 ^ cgp_core_202;
  assign cgp_core_207 = cgp_core_196 & cgp_core_202;
  assign cgp_core_208 = cgp_core_198 ^ cgp_core_204;
  assign cgp_core_209 = cgp_core_198 & cgp_core_204;
  assign cgp_core_210 = cgp_core_208 ^ cgp_core_207;
  assign cgp_core_211 = cgp_core_208 & cgp_core_207;
  assign cgp_core_212 = cgp_core_209 | cgp_core_211;
  assign cgp_core_216 = input_a[18] & input_a[20];
  assign cgp_core_217 = input_a[18] & input_a[36];
  assign cgp_core_218 = input_a[30] ^ input_a[31];
  assign cgp_core_219 = input_a[30] & input_a[31];
  assign cgp_core_220 = input_a[29] ^ cgp_core_218;
  assign cgp_core_221 = input_a[29] & cgp_core_218;
  assign cgp_core_222 = cgp_core_219 | cgp_core_221;
  assign cgp_core_223 = input_a[10] ^ input_a[32];
  assign cgp_core_224 = input_a[33] ^ input_a[34];
  assign cgp_core_225 = input_a[33] & input_a[34];
  assign cgp_core_226 = input_a[32] ^ cgp_core_224;
  assign cgp_core_227 = input_a[32] & cgp_core_224;
  assign cgp_core_228 = cgp_core_225 | cgp_core_227;
  assign cgp_core_229 = input_a[35] | input_a[23];
  assign cgp_core_230 = cgp_core_220 ^ cgp_core_226;
  assign cgp_core_231 = cgp_core_220 & cgp_core_226;
  assign cgp_core_232 = cgp_core_222 ^ cgp_core_228;
  assign cgp_core_233 = cgp_core_222 & cgp_core_228;
  assign cgp_core_234 = cgp_core_232 ^ cgp_core_231;
  assign cgp_core_235 = cgp_core_232 & cgp_core_231;
  assign cgp_core_236 = cgp_core_233 | cgp_core_235;
  assign cgp_core_240 = ~(input_a[34] ^ input_a[40]);
  assign cgp_core_242 = cgp_core_206 ^ cgp_core_230;
  assign cgp_core_243 = cgp_core_206 & cgp_core_230;
  assign cgp_core_244 = cgp_core_210 ^ cgp_core_234;
  assign cgp_core_245 = cgp_core_210 & cgp_core_234;
  assign cgp_core_246 = cgp_core_244 ^ cgp_core_243;
  assign cgp_core_247 = cgp_core_244 & cgp_core_243;
  assign cgp_core_248 = cgp_core_245 | cgp_core_247;
  assign cgp_core_249 = cgp_core_212 ^ cgp_core_236;
  assign cgp_core_250 = cgp_core_212 & cgp_core_236;
  assign cgp_core_251 = cgp_core_249 ^ cgp_core_248;
  assign cgp_core_252 = cgp_core_249 & cgp_core_248;
  assign cgp_core_253 = cgp_core_250 | cgp_core_252;
  assign cgp_core_255 = input_a[15] | input_a[16];
  assign cgp_core_257 = input_a[9] ^ input_a[9];
  assign cgp_core_258 = ~input_a[12];
  assign cgp_core_259 = input_a[36] | input_a[37];
  assign cgp_core_260 = input_a[36] & input_a[37];
  assign cgp_core_261 = input_a[2] | input_a[2];
  assign cgp_core_262 = input_a[35] & cgp_core_259;
  assign cgp_core_263 = cgp_core_260 | cgp_core_262;
  assign cgp_core_265 = input_a[39] | input_a[40];
  assign cgp_core_266 = input_a[39] & input_a[40];
  assign cgp_core_267 = ~(input_a[30] ^ input_a[27]);
  assign cgp_core_268 = input_a[38] & cgp_core_265;
  assign cgp_core_269 = cgp_core_266 | cgp_core_268;
  assign cgp_core_272 = ~input_a[26];
  assign cgp_core_273 = cgp_core_263 ^ cgp_core_269;
  assign cgp_core_274 = cgp_core_263 & cgp_core_269;
  assign cgp_core_276 = ~input_a[24];
  assign cgp_core_279 = input_a[33] | input_a[31];
  assign cgp_core_281 = ~(input_a[20] ^ input_a[18]);
  assign cgp_core_282 = input_a[32] ^ input_a[9];
  assign cgp_core_283 = input_a[42] ^ input_a[43];
  assign cgp_core_284 = input_a[42] & input_a[43];
  assign cgp_core_285 = input_a[41] ^ cgp_core_283;
  assign cgp_core_286 = input_a[41] & cgp_core_283;
  assign cgp_core_287 = cgp_core_284 | cgp_core_286;
  assign cgp_core_288 = ~input_a[7];
  assign cgp_core_289 = input_a[45] ^ input_a[46];
  assign cgp_core_290 = input_a[45] & input_a[46];
  assign cgp_core_291 = input_a[44] ^ cgp_core_289;
  assign cgp_core_292 = input_a[44] & cgp_core_289;
  assign cgp_core_293 = cgp_core_290 | cgp_core_292;
  assign cgp_core_294 = ~(input_a[39] | input_a[15]);
  assign cgp_core_295 = cgp_core_285 ^ cgp_core_291;
  assign cgp_core_296 = cgp_core_285 & cgp_core_291;
  assign cgp_core_297 = cgp_core_287 ^ cgp_core_293;
  assign cgp_core_298 = cgp_core_287 & cgp_core_293;
  assign cgp_core_299 = cgp_core_297 ^ cgp_core_296;
  assign cgp_core_300 = cgp_core_297 & cgp_core_296;
  assign cgp_core_301 = cgp_core_298 | cgp_core_300;
  assign cgp_core_303 = ~input_a[31];
  assign cgp_core_305 = ~input_a[44];
  assign cgp_core_306 = input_a[44] & input_a[45];
  assign cgp_core_307 = ~cgp_core_295;
  assign cgp_core_309 = cgp_core_273 ^ cgp_core_299;
  assign cgp_core_310 = cgp_core_273 & cgp_core_299;
  assign cgp_core_311 = cgp_core_309 ^ cgp_core_295;
  assign cgp_core_312 = cgp_core_309 & cgp_core_295;
  assign cgp_core_313 = cgp_core_310 | cgp_core_312;
  assign cgp_core_314 = cgp_core_274 ^ cgp_core_301;
  assign cgp_core_315 = cgp_core_274 & cgp_core_301;
  assign cgp_core_316 = cgp_core_314 ^ cgp_core_313;
  assign cgp_core_317 = cgp_core_314 & cgp_core_313;
  assign cgp_core_318 = cgp_core_315 | cgp_core_317;
  assign cgp_core_320 = ~(input_a[34] | input_a[37]);
  assign cgp_core_324 = cgp_core_242 ^ cgp_core_307;
  assign cgp_core_325 = cgp_core_242 & cgp_core_307;
  assign cgp_core_326 = cgp_core_246 ^ cgp_core_311;
  assign cgp_core_327 = cgp_core_246 & cgp_core_311;
  assign cgp_core_328 = cgp_core_326 ^ cgp_core_325;
  assign cgp_core_329 = cgp_core_326 & cgp_core_325;
  assign cgp_core_330 = cgp_core_327 | cgp_core_329;
  assign cgp_core_331 = cgp_core_251 ^ cgp_core_316;
  assign cgp_core_332 = cgp_core_251 & cgp_core_316;
  assign cgp_core_333 = cgp_core_331 ^ cgp_core_330;
  assign cgp_core_334 = cgp_core_331 & cgp_core_330;
  assign cgp_core_335 = cgp_core_332 | cgp_core_334;
  assign cgp_core_336 = cgp_core_253 ^ cgp_core_318;
  assign cgp_core_337 = cgp_core_253 & cgp_core_318;
  assign cgp_core_338 = cgp_core_336 ^ cgp_core_335;
  assign cgp_core_339 = cgp_core_336 & cgp_core_335;
  assign cgp_core_340 = cgp_core_337 | cgp_core_339;
  assign cgp_core_345 = input_a[5] & input_a[26];
  assign cgp_core_346 = cgp_core_172 ^ cgp_core_324;
  assign cgp_core_347 = cgp_core_172 & cgp_core_324;
  assign cgp_core_348 = cgp_core_176 ^ cgp_core_328;
  assign cgp_core_349 = cgp_core_176 & cgp_core_328;
  assign cgp_core_350 = cgp_core_348 ^ cgp_core_347;
  assign cgp_core_351 = cgp_core_348 & cgp_core_347;
  assign cgp_core_352 = cgp_core_349 | cgp_core_351;
  assign cgp_core_353 = cgp_core_181 ^ cgp_core_333;
  assign cgp_core_354 = cgp_core_181 & cgp_core_333;
  assign cgp_core_355 = cgp_core_353 ^ cgp_core_352;
  assign cgp_core_356 = cgp_core_353 & cgp_core_352;
  assign cgp_core_357 = cgp_core_354 | cgp_core_356;
  assign cgp_core_358 = cgp_core_186 ^ cgp_core_338;
  assign cgp_core_359 = cgp_core_186 & cgp_core_338;
  assign cgp_core_360 = cgp_core_358 ^ cgp_core_357;
  assign cgp_core_361 = cgp_core_358 & cgp_core_357;
  assign cgp_core_362 = cgp_core_359 | cgp_core_361;
  assign cgp_core_363 = cgp_core_188 ^ cgp_core_340;
  assign cgp_core_364 = cgp_core_188 & cgp_core_340;
  assign cgp_core_365 = cgp_core_363 ^ cgp_core_362;
  assign cgp_core_366 = cgp_core_363 & cgp_core_362;
  assign cgp_core_367 = cgp_core_364 | cgp_core_366;
  assign cgp_core_369 = input_a[41] & input_a[1];
  assign cgp_core_370 = input_a[2] | input_a[10];

  assign cgp_out[0] = cgp_core_346;
  assign cgp_out[1] = cgp_core_350;
  assign cgp_out[2] = cgp_core_355;
  assign cgp_out[3] = cgp_core_360;
  assign cgp_out[4] = cgp_core_365;
  assign cgp_out[5] = cgp_core_367;
endmodule

module cmp_neg(input [29:0] input_a, output [4:0] cgp_out);
  wire cgp_core_033;
  wire cgp_core_034;
  wire cgp_core_036;
  wire cgp_core_037;
  wire cgp_core_038;
  wire cgp_core_039;
  wire cgp_core_040;
  wire cgp_core_041;
  wire cgp_core_044;
  wire cgp_core_045;
  wire cgp_core_047;
  wire cgp_core_049;
  wire cgp_core_050;
  wire cgp_core_051;
  wire cgp_core_052;
  wire cgp_core_053;
  wire cgp_core_054;
  wire cgp_core_055;
  wire cgp_core_056;
  wire cgp_core_057;
  wire cgp_core_058;
  wire cgp_core_061;
  wire cgp_core_062;
  wire cgp_core_063;
  wire cgp_core_064;
  wire cgp_core_065;
  wire cgp_core_067;
  wire cgp_core_068;
  wire cgp_core_069;
  wire cgp_core_070;
  wire cgp_core_072;
  wire cgp_core_073;
  wire cgp_core_074;
  wire cgp_core_075;
  wire cgp_core_076;
  wire cgp_core_077;
  wire cgp_core_078;
  wire cgp_core_079;
  wire cgp_core_080;
  wire cgp_core_083;
  wire cgp_core_084;
  wire cgp_core_085;
  wire cgp_core_086;
  wire cgp_core_087;
  wire cgp_core_088;
  wire cgp_core_089;
  wire cgp_core_090;
  wire cgp_core_091;
  wire cgp_core_092;
  wire cgp_core_093;
  wire cgp_core_096;
  wire cgp_core_097;
  wire cgp_core_098;
  wire cgp_core_100;
  wire cgp_core_102;
  wire cgp_core_103;
  wire cgp_core_104;
  wire cgp_core_105;
  wire cgp_core_106;
  wire cgp_core_107;
  wire cgp_core_108;
  wire cgp_core_109;
  wire cgp_core_110;
  wire cgp_core_112;
  wire cgp_core_113;
  wire cgp_core_114;
  wire cgp_core_115;
  wire cgp_core_116;
  wire cgp_core_117;
  wire cgp_core_118;
  wire cgp_core_119;
  wire cgp_core_122;
  wire cgp_core_123;
  wire cgp_core_124;
  wire cgp_core_125;
  wire cgp_core_126;
  wire cgp_core_128;
  wire cgp_core_130;
  wire cgp_core_131;
  wire cgp_core_137;
  wire cgp_core_141;
  wire cgp_core_142;
  wire cgp_core_143;
  wire cgp_core_144;
  wire cgp_core_145;
  wire cgp_core_146;
  wire cgp_core_147;
  wire cgp_core_148;
  wire cgp_core_149;
  wire cgp_core_152;
  wire cgp_core_153;
  wire cgp_core_154;
  wire cgp_core_155;
  wire cgp_core_156;
  wire cgp_core_157;
  wire cgp_core_158;
  wire cgp_core_159;
  wire cgp_core_160;
  wire cgp_core_163;
  wire cgp_core_164;
  wire cgp_core_165;
  wire cgp_core_166;
  wire cgp_core_167;
  wire cgp_core_168;
  wire cgp_core_169;
  wire cgp_core_170;
  wire cgp_core_171;
  wire cgp_core_172;
  wire cgp_core_173;
  wire cgp_core_175;
  wire cgp_core_177;
  wire cgp_core_178;
  wire cgp_core_179;
  wire cgp_core_180;
  wire cgp_core_181;
  wire cgp_core_182;
  wire cgp_core_183;
  wire cgp_core_184;
  wire cgp_core_185;
  wire cgp_core_186;
  wire cgp_core_188;
  wire cgp_core_189;
  wire cgp_core_190;
  wire cgp_core_191;
  wire cgp_core_192;
  wire cgp_core_193;
  wire cgp_core_196;
  wire cgp_core_197;
  wire cgp_core_199;
  wire cgp_core_200;
  wire cgp_core_201;
  wire cgp_core_202;
  wire cgp_core_203;
  wire cgp_core_204;
  wire cgp_core_205;
  wire cgp_core_206;
  wire cgp_core_207;
  wire cgp_core_208;
  wire cgp_core_211;
  wire cgp_core_212;
  wire cgp_core_213;

  assign cgp_core_033 = input_a[1] & input_a[18];
  assign cgp_core_034 = ~input_a[0];
  assign cgp_core_036 = cgp_core_033 ^ input_a[0];
  assign cgp_core_037 = cgp_core_033 & input_a[0];
  assign cgp_core_038 = input_a[15] & input_a[23];
  assign cgp_core_039 = input_a[3] & input_a[4];
  assign cgp_core_040 = input_a[7] & input_a[20];
  assign cgp_core_041 = input_a[2] & input_a[19];
  assign cgp_core_044 = cgp_core_039 ^ cgp_core_041;
  assign cgp_core_045 = cgp_core_039 & cgp_core_041;
  assign cgp_core_047 = input_a[18] | input_a[16];
  assign cgp_core_049 = ~(input_a[11] & input_a[17]);
  assign cgp_core_050 = cgp_core_034 & input_a[20];
  assign cgp_core_051 = cgp_core_036 ^ cgp_core_044;
  assign cgp_core_052 = cgp_core_036 & cgp_core_044;
  assign cgp_core_053 = cgp_core_051 ^ cgp_core_050;
  assign cgp_core_054 = cgp_core_051 & cgp_core_050;
  assign cgp_core_055 = cgp_core_052 | cgp_core_054;
  assign cgp_core_056 = cgp_core_037 ^ cgp_core_045;
  assign cgp_core_057 = cgp_core_037 & cgp_core_045;
  assign cgp_core_058 = cgp_core_056 | cgp_core_055;
  assign cgp_core_061 = input_a[7] ^ input_a[8];
  assign cgp_core_062 = input_a[7] & input_a[8];
  assign cgp_core_063 = ~(input_a[9] & input_a[10]);
  assign cgp_core_064 = input_a[9] & input_a[10];
  assign cgp_core_065 = cgp_core_061 ^ cgp_core_063;
  assign cgp_core_067 = input_a[8] ^ cgp_core_064;
  assign cgp_core_068 = cgp_core_062 & cgp_core_064;
  assign cgp_core_069 = cgp_core_067 | cgp_core_061;
  assign cgp_core_070 = input_a[7] & input_a[20];
  assign cgp_core_072 = input_a[11] ^ input_a[12];
  assign cgp_core_073 = input_a[11] & input_a[12];
  assign cgp_core_074 = input_a[13] ^ input_a[14];
  assign cgp_core_075 = input_a[13] & input_a[14];
  assign cgp_core_076 = cgp_core_072 ^ cgp_core_074;
  assign cgp_core_077 = cgp_core_072 & cgp_core_074;
  assign cgp_core_078 = cgp_core_073 ^ cgp_core_075;
  assign cgp_core_079 = cgp_core_073 & cgp_core_075;
  assign cgp_core_080 = cgp_core_078 | cgp_core_077;
  assign cgp_core_083 = ~input_a[19];
  assign cgp_core_084 = cgp_core_065 & cgp_core_076;
  assign cgp_core_085 = cgp_core_069 ^ cgp_core_080;
  assign cgp_core_086 = cgp_core_069 & cgp_core_080;
  assign cgp_core_087 = cgp_core_085 ^ cgp_core_084;
  assign cgp_core_088 = cgp_core_085 & cgp_core_084;
  assign cgp_core_089 = cgp_core_086 | cgp_core_088;
  assign cgp_core_090 = cgp_core_068 ^ cgp_core_079;
  assign cgp_core_091 = cgp_core_068 & cgp_core_079;
  assign cgp_core_092 = cgp_core_090 | cgp_core_089;
  assign cgp_core_093 = ~(input_a[28] & input_a[18]);
  assign cgp_core_096 = input_a[11] ^ input_a[17];
  assign cgp_core_097 = ~input_a[2];
  assign cgp_core_098 = cgp_core_053 & cgp_core_087;
  assign cgp_core_100 = ~(input_a[0] ^ input_a[18]);
  assign cgp_core_102 = cgp_core_058 ^ cgp_core_092;
  assign cgp_core_103 = cgp_core_058 & cgp_core_092;
  assign cgp_core_104 = cgp_core_102 ^ cgp_core_098;
  assign cgp_core_105 = cgp_core_102 & cgp_core_098;
  assign cgp_core_106 = cgp_core_103 | cgp_core_105;
  assign cgp_core_107 = cgp_core_057 ^ cgp_core_091;
  assign cgp_core_108 = cgp_core_057 & cgp_core_091;
  assign cgp_core_109 = cgp_core_107 | cgp_core_106;
  assign cgp_core_110 = ~(input_a[8] | input_a[18]);
  assign cgp_core_112 = ~(input_a[20] | input_a[4]);
  assign cgp_core_113 = input_a[17] & input_a[21];
  assign cgp_core_114 = ~(input_a[22] & input_a[0]);
  assign cgp_core_115 = input_a[6] & input_a[5];
  assign cgp_core_116 = cgp_core_113 | cgp_core_115;
  assign cgp_core_117 = ~(input_a[29] | input_a[24]);
  assign cgp_core_118 = ~input_a[27];
  assign cgp_core_119 = input_a[23] ^ input_a[21];
  assign cgp_core_122 = input_a[9] | input_a[4];
  assign cgp_core_123 = ~(input_a[14] & input_a[27]);
  assign cgp_core_124 = ~input_a[0];
  assign cgp_core_125 = input_a[9] ^ input_a[11];
  assign cgp_core_126 = ~(input_a[13] | input_a[20]);
  assign cgp_core_128 = input_a[26] | input_a[17];
  assign cgp_core_130 = input_a[17] ^ input_a[29];
  assign cgp_core_131 = ~cgp_core_116;
  assign cgp_core_137 = input_a[17] & input_a[21];
  assign cgp_core_141 = ~input_a[23];
  assign cgp_core_142 = input_a[26] | input_a[22];
  assign cgp_core_143 = input_a[24] ^ input_a[25];
  assign cgp_core_144 = input_a[24] & input_a[25];
  assign cgp_core_145 = cgp_core_141 ^ cgp_core_143;
  assign cgp_core_146 = cgp_core_141 & cgp_core_143;
  assign cgp_core_147 = input_a[23] ^ cgp_core_144;
  assign cgp_core_148 = input_a[23] & cgp_core_144;
  assign cgp_core_149 = cgp_core_147 | cgp_core_146;
  assign cgp_core_152 = input_a[26] ^ input_a[27];
  assign cgp_core_153 = input_a[26] & input_a[27];
  assign cgp_core_154 = input_a[28] ^ input_a[29];
  assign cgp_core_155 = input_a[28] & input_a[29];
  assign cgp_core_156 = cgp_core_152 ^ cgp_core_154;
  assign cgp_core_157 = cgp_core_152 & cgp_core_154;
  assign cgp_core_158 = cgp_core_153 ^ cgp_core_155;
  assign cgp_core_159 = cgp_core_153 & cgp_core_155;
  assign cgp_core_160 = cgp_core_158 | cgp_core_157;
  assign cgp_core_163 = cgp_core_145 ^ cgp_core_156;
  assign cgp_core_164 = cgp_core_145 & cgp_core_156;
  assign cgp_core_165 = cgp_core_149 ^ cgp_core_160;
  assign cgp_core_166 = cgp_core_149 & cgp_core_160;
  assign cgp_core_167 = cgp_core_165 ^ cgp_core_164;
  assign cgp_core_168 = cgp_core_165 & cgp_core_164;
  assign cgp_core_169 = cgp_core_166 | cgp_core_168;
  assign cgp_core_170 = cgp_core_148 ^ cgp_core_159;
  assign cgp_core_171 = input_a[23] & cgp_core_159;
  assign cgp_core_172 = cgp_core_170 | cgp_core_169;
  assign cgp_core_173 = ~input_a[19];
  assign cgp_core_175 = input_a[23] ^ input_a[3];
  assign cgp_core_177 = cgp_core_131 ^ cgp_core_167;
  assign cgp_core_178 = cgp_core_131 & cgp_core_167;
  assign cgp_core_179 = cgp_core_177 ^ cgp_core_163;
  assign cgp_core_180 = cgp_core_177 & cgp_core_163;
  assign cgp_core_181 = cgp_core_178 | cgp_core_180;
  assign cgp_core_182 = cgp_core_116 ^ cgp_core_172;
  assign cgp_core_183 = cgp_core_116 & cgp_core_172;
  assign cgp_core_184 = cgp_core_182 ^ cgp_core_181;
  assign cgp_core_185 = cgp_core_182 & cgp_core_181;
  assign cgp_core_186 = cgp_core_183 | cgp_core_185;
  assign cgp_core_188 = ~input_a[18];
  assign cgp_core_189 = cgp_core_171 | cgp_core_186;
  assign cgp_core_190 = input_a[23] & input_a[17];
  assign cgp_core_191 = ~(input_a[8] | input_a[28]);
  assign cgp_core_192 = ~input_a[1];
  assign cgp_core_193 = input_a[16] & input_a[22];
  assign cgp_core_196 = cgp_core_179 ^ cgp_core_193;
  assign cgp_core_197 = cgp_core_179 & cgp_core_193;
  assign cgp_core_199 = cgp_core_104 ^ cgp_core_184;
  assign cgp_core_200 = cgp_core_104 & cgp_core_184;
  assign cgp_core_201 = cgp_core_199 ^ cgp_core_197;
  assign cgp_core_202 = cgp_core_199 & cgp_core_197;
  assign cgp_core_203 = cgp_core_200 | cgp_core_202;
  assign cgp_core_204 = cgp_core_109 ^ cgp_core_189;
  assign cgp_core_205 = cgp_core_109 & cgp_core_189;
  assign cgp_core_206 = cgp_core_204 ^ cgp_core_203;
  assign cgp_core_207 = cgp_core_204 & cgp_core_203;
  assign cgp_core_208 = cgp_core_205 | cgp_core_207;
  assign cgp_core_211 = cgp_core_108 | cgp_core_208;
  assign cgp_core_212 = ~(input_a[18] & input_a[20]);
  assign cgp_core_213 = ~input_a[16];

  assign cgp_out[0] = input_a[15];
  assign cgp_out[1] = cgp_core_196;
  assign cgp_out[2] = cgp_core_201;
  assign cgp_out[3] = cgp_core_206;
  assign cgp_out[4] = cgp_core_211;
endmodule
module pcc(input [46:0] pos, input [29:0] neg, output outval);
    wire [5:0] cnt_pos;
    wire [4:0] cnt_neg;

    cmp_pos ipos(pos, cnt_pos);
    cmp_neg ineg(neg, cnt_neg);

    assign outval = (cnt_pos >= cnt_neg);
endmodule
