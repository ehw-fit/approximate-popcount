// 
// This code is a part of TNNApprox library distributed under The MIT License.
// When used, please cite the following article: V. Mrazek, A. Kokkinis, P. Papanikolaou, Z. Vasicek, K. Siozis, G. Tzimpragos, M. Tahoori, G. Zervakis "Evolutionary Approximation of Ternary Neurons \for On-sensor Printed Neural Networks" International Conference on Computer Aided Design (ICCAD), 2024
// 
// MAE=4.34694
// WCE=18.0
// EP=0.92618%
// Printed PDK parameters:
//  Area=0.0
//  Delay=0.0
//  Power=0.0

module popcount23_2it3(input [22:0] input_a, output [4:0] popcount23_2it3_out);
  wire popcount23_2it3_core_025;
  wire popcount23_2it3_core_026;
  wire popcount23_2it3_core_027;
  wire popcount23_2it3_core_029;
  wire popcount23_2it3_core_033;
  wire popcount23_2it3_core_034;
  wire popcount23_2it3_core_035;
  wire popcount23_2it3_core_038;
  wire popcount23_2it3_core_040;
  wire popcount23_2it3_core_043;
  wire popcount23_2it3_core_045;
  wire popcount23_2it3_core_046;
  wire popcount23_2it3_core_047;
  wire popcount23_2it3_core_048;
  wire popcount23_2it3_core_052;
  wire popcount23_2it3_core_056;
  wire popcount23_2it3_core_058;
  wire popcount23_2it3_core_059;
  wire popcount23_2it3_core_062;
  wire popcount23_2it3_core_064;
  wire popcount23_2it3_core_066;
  wire popcount23_2it3_core_067;
  wire popcount23_2it3_core_069;
  wire popcount23_2it3_core_070;
  wire popcount23_2it3_core_072_not;
  wire popcount23_2it3_core_073;
  wire popcount23_2it3_core_074;
  wire popcount23_2it3_core_078;
  wire popcount23_2it3_core_080;
  wire popcount23_2it3_core_081;
  wire popcount23_2it3_core_082;
  wire popcount23_2it3_core_083;
  wire popcount23_2it3_core_084;
  wire popcount23_2it3_core_085;
  wire popcount23_2it3_core_087;
  wire popcount23_2it3_core_088;
  wire popcount23_2it3_core_090;
  wire popcount23_2it3_core_092;
  wire popcount23_2it3_core_094;
  wire popcount23_2it3_core_095;
  wire popcount23_2it3_core_096;
  wire popcount23_2it3_core_097;
  wire popcount23_2it3_core_098;
  wire popcount23_2it3_core_099;
  wire popcount23_2it3_core_103;
  wire popcount23_2it3_core_104_not;
  wire popcount23_2it3_core_105;
  wire popcount23_2it3_core_107;
  wire popcount23_2it3_core_108;
  wire popcount23_2it3_core_110;
  wire popcount23_2it3_core_112;
  wire popcount23_2it3_core_115;
  wire popcount23_2it3_core_121;
  wire popcount23_2it3_core_122;
  wire popcount23_2it3_core_123;
  wire popcount23_2it3_core_124;
  wire popcount23_2it3_core_125;
  wire popcount23_2it3_core_126;
  wire popcount23_2it3_core_128;
  wire popcount23_2it3_core_129;
  wire popcount23_2it3_core_130;
  wire popcount23_2it3_core_132;
  wire popcount23_2it3_core_134;
  wire popcount23_2it3_core_135;
  wire popcount23_2it3_core_138;
  wire popcount23_2it3_core_140;
  wire popcount23_2it3_core_141;
  wire popcount23_2it3_core_142_not;
  wire popcount23_2it3_core_143;
  wire popcount23_2it3_core_145;
  wire popcount23_2it3_core_146;
  wire popcount23_2it3_core_147;
  wire popcount23_2it3_core_148;
  wire popcount23_2it3_core_149;
  wire popcount23_2it3_core_150;
  wire popcount23_2it3_core_153;
  wire popcount23_2it3_core_154;
  wire popcount23_2it3_core_155;
  wire popcount23_2it3_core_160;
  wire popcount23_2it3_core_161;
  wire popcount23_2it3_core_162;
  wire popcount23_2it3_core_163;
  wire popcount23_2it3_core_165;
  wire popcount23_2it3_core_167;
  wire popcount23_2it3_core_168;

  assign popcount23_2it3_core_025 = ~input_a[8];
  assign popcount23_2it3_core_026 = ~input_a[6];
  assign popcount23_2it3_core_027 = ~input_a[1];
  assign popcount23_2it3_core_029 = ~(input_a[16] | input_a[1]);
  assign popcount23_2it3_core_033 = ~(input_a[5] & input_a[9]);
  assign popcount23_2it3_core_034 = input_a[18] | input_a[10];
  assign popcount23_2it3_core_035 = input_a[18] | input_a[7];
  assign popcount23_2it3_core_038 = ~(input_a[0] & input_a[21]);
  assign popcount23_2it3_core_040 = input_a[17] & input_a[21];
  assign popcount23_2it3_core_043 = ~(input_a[16] & input_a[22]);
  assign popcount23_2it3_core_045 = ~(input_a[5] | input_a[17]);
  assign popcount23_2it3_core_046 = input_a[13] ^ input_a[17];
  assign popcount23_2it3_core_047 = input_a[0] | input_a[6];
  assign popcount23_2it3_core_048 = ~(input_a[19] & input_a[3]);
  assign popcount23_2it3_core_052 = input_a[22] ^ input_a[2];
  assign popcount23_2it3_core_056 = ~(input_a[17] & input_a[18]);
  assign popcount23_2it3_core_058 = ~(input_a[10] ^ input_a[14]);
  assign popcount23_2it3_core_059 = input_a[6] | input_a[9];
  assign popcount23_2it3_core_062 = ~(input_a[15] ^ input_a[13]);
  assign popcount23_2it3_core_064 = input_a[21] ^ input_a[12];
  assign popcount23_2it3_core_066 = ~(input_a[5] | input_a[5]);
  assign popcount23_2it3_core_067 = ~(input_a[19] ^ input_a[13]);
  assign popcount23_2it3_core_069 = input_a[9] & input_a[21];
  assign popcount23_2it3_core_070 = input_a[19] | input_a[16];
  assign popcount23_2it3_core_072_not = ~input_a[21];
  assign popcount23_2it3_core_073 = input_a[12] & input_a[5];
  assign popcount23_2it3_core_074 = input_a[7] & input_a[19];
  assign popcount23_2it3_core_078 = input_a[1] & input_a[19];
  assign popcount23_2it3_core_080 = ~(input_a[5] & input_a[5]);
  assign popcount23_2it3_core_081 = input_a[12] & input_a[21];
  assign popcount23_2it3_core_082 = input_a[15] & input_a[22];
  assign popcount23_2it3_core_083 = ~(input_a[3] ^ input_a[17]);
  assign popcount23_2it3_core_084 = ~(input_a[13] & input_a[19]);
  assign popcount23_2it3_core_085 = ~(input_a[12] ^ input_a[20]);
  assign popcount23_2it3_core_087 = ~input_a[4];
  assign popcount23_2it3_core_088 = ~input_a[7];
  assign popcount23_2it3_core_090 = ~(input_a[17] | input_a[12]);
  assign popcount23_2it3_core_092 = ~(input_a[22] & input_a[14]);
  assign popcount23_2it3_core_094 = ~input_a[1];
  assign popcount23_2it3_core_095 = ~(input_a[20] | input_a[6]);
  assign popcount23_2it3_core_096 = ~(input_a[18] | input_a[5]);
  assign popcount23_2it3_core_097 = input_a[10] & input_a[7];
  assign popcount23_2it3_core_098 = input_a[5] ^ input_a[12];
  assign popcount23_2it3_core_099 = ~input_a[22];
  assign popcount23_2it3_core_103 = ~(input_a[6] ^ input_a[7]);
  assign popcount23_2it3_core_104_not = ~input_a[7];
  assign popcount23_2it3_core_105 = input_a[20] ^ input_a[21];
  assign popcount23_2it3_core_107 = ~(input_a[19] & input_a[19]);
  assign popcount23_2it3_core_108 = ~(input_a[0] ^ input_a[3]);
  assign popcount23_2it3_core_110 = input_a[21] & input_a[15];
  assign popcount23_2it3_core_112 = input_a[10] & input_a[3];
  assign popcount23_2it3_core_115 = input_a[16] & input_a[22];
  assign popcount23_2it3_core_121 = ~input_a[20];
  assign popcount23_2it3_core_122 = input_a[20] | input_a[17];
  assign popcount23_2it3_core_123 = input_a[19] | input_a[11];
  assign popcount23_2it3_core_124 = ~(input_a[4] | input_a[21]);
  assign popcount23_2it3_core_125 = ~(input_a[13] & input_a[3]);
  assign popcount23_2it3_core_126 = ~(input_a[14] & input_a[6]);
  assign popcount23_2it3_core_128 = ~input_a[9];
  assign popcount23_2it3_core_129 = ~input_a[11];
  assign popcount23_2it3_core_130 = input_a[10] | input_a[5];
  assign popcount23_2it3_core_132 = input_a[18] | input_a[17];
  assign popcount23_2it3_core_134 = ~(input_a[3] & input_a[4]);
  assign popcount23_2it3_core_135 = ~input_a[20];
  assign popcount23_2it3_core_138 = input_a[18] ^ input_a[21];
  assign popcount23_2it3_core_140 = ~(input_a[3] & input_a[3]);
  assign popcount23_2it3_core_141 = input_a[9] & input_a[11];
  assign popcount23_2it3_core_142_not = ~input_a[14];
  assign popcount23_2it3_core_143 = input_a[12] ^ input_a[4];
  assign popcount23_2it3_core_145 = input_a[0] & input_a[21];
  assign popcount23_2it3_core_146 = ~(input_a[21] | input_a[12]);
  assign popcount23_2it3_core_147 = ~(input_a[4] ^ input_a[1]);
  assign popcount23_2it3_core_148 = ~(input_a[1] & input_a[0]);
  assign popcount23_2it3_core_149 = input_a[21] ^ input_a[1];
  assign popcount23_2it3_core_150 = ~(input_a[9] & input_a[13]);
  assign popcount23_2it3_core_153 = input_a[10] & input_a[3];
  assign popcount23_2it3_core_154 = input_a[1] | input_a[7];
  assign popcount23_2it3_core_155 = ~(input_a[19] ^ input_a[10]);
  assign popcount23_2it3_core_160 = ~(input_a[13] & input_a[8]);
  assign popcount23_2it3_core_161 = ~(input_a[1] | input_a[0]);
  assign popcount23_2it3_core_162 = input_a[7] | input_a[6];
  assign popcount23_2it3_core_163 = input_a[8] | input_a[7];
  assign popcount23_2it3_core_165 = ~(input_a[19] ^ input_a[21]);
  assign popcount23_2it3_core_167 = input_a[6] & input_a[1];
  assign popcount23_2it3_core_168 = input_a[1] & input_a[11];

  assign popcount23_2it3_out[0] = input_a[20];
  assign popcount23_2it3_out[1] = 1'b1;
  assign popcount23_2it3_out[2] = input_a[19];
  assign popcount23_2it3_out[3] = input_a[13];
  assign popcount23_2it3_out[4] = 1'b0;
endmodule